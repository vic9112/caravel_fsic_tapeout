.GLOBAL VDD VSS
.GLOBAL VBP VBN

*.CONNECT VBP VDD
*.CONNECT VBN VSS


.subckt SAEDRVT14_ADDF_V1_0P5 VDD VSS VBP VBN S CO A B CI
Mxmn12 CO con VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn11 S net86 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn9 net102 con VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn8 VSS A net94 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn7 net94 B net102 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn6 net94 con net86 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn5 net86 CI net102 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn4 net82 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn3 con A net82 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn2 net70 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn1 net70 A VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn0 con CI net70 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp11 CO con VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp10 S net86 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp9 net135 con net86 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp8 net86 CI net139 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp7 net139 B net135 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp6 VDD A net135 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp5 net139 con VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp4 con A net123 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp3 net123 B VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp2 net111 B VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp1 con CI net111 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 net111 A VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ADDF_V1_0P5




.subckt SAEDRVT14_ADDF_V1_1 VDD VSS VBP VBN S CO A B CI
Mxmn12 CO con VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn11 S net86 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn9 net102 con VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn8 VSS A net94 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn7 net94 B net102 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn6 net94 con net86 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn5 net86 CI net102 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn4 net82 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 con A net82 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn2 net70 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn1 net70 A VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 con CI net70 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp11 CO con VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp10 S net86 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp9 net135 con net86 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp8 net86 CI net139 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp7 net139 B net135 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp6 VDD A net135 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp5 net139 con VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp4 con A net123 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp3 net123 B VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp2 net111 B VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 con CI net111 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp0 net111 A VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ADDF_V1_1




.subckt SAEDRVT14_ADDF_V1_2 VDD VSS VBP VBN S CO A B CI
Mxmn12 CO con VSS VBN n08 l=0.014u nf=2 m=2 nfin=4
Mxmn11 S net86 VSS VBN n08 l=0.014u nf=2 m=2 nfin=4
Mxmn9 net102 con VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn8 VSS A net94 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn7 net94 B net102 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn6 net94 con net86 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn5 net86 CI net102 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn4 net82 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 con A net82 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn2 net70 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn1 net70 A VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 con CI net70 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp11 CO con VDD VBP p08 l=0.014u nf=2 m=2 nfin=4
Mxmp10 S net86 VDD VBP p08 l=0.014u nf=2 m=2 nfin=4
Mxmp9 net135 con net86 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp8 net86 CI net139 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp7 net139 B net135 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp6 VDD A net135 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp5 net139 con VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp4 con A net123 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp3 net123 B VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp2 net111 B VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 con CI net111 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp0 net111 A VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ADDF_V1_2




.subckt SAEDRVT14_ADDF_V2_0P5 VDD VSS VBP VBN S CO A B CI
Mxmn28 net60 pn net74 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn27 net56 p net74 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn26 CO net74 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn25 S net67 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn24 pn p VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn23 net58 p net67 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn22 net56 pn net67 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn21 net56 CI VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmn20 net58 net56 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn18 net18 B p VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn17 net60 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn16 net59 net60 p VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn15 net59 net18 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn14 net18 A VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmpdummy VDD A VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp26 net60 p net74 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp25 CO net74 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp24 net56 pn net74 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp23 S net67 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp22 pn p VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp21 net56 p net67 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp20 net049 pn net67 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp19 net56 CI VDD VBP p08 l=0.014u nf=2 m=1 nfin=2
Mxmp18 net049 net56 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp16 net18 net60 p VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp15 net60 B VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp14 net050 B p VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp13 net050 net18 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp12 net18 A VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ADDF_V2_0P5




.subckt SAEDRVT14_ADDF_V2_1 VDD VSS VBP VBN S CO A B CI
Mxmp26 net60 p net74 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp25 CO net74 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp24 net56 pn net74 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp23 S net67 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp22 pn p VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp21 net56 p net67 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp20 net050 pn net67 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp19 net56 CI VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp18 net050 net56 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp16 net18 net60 p VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp15 net60 B VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp14 net051 B p VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp13 net051 net18 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp12 net18 A VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp13 VDD A VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmn28 net60 pn net74 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn27 net56 p net74 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn26 CO net74 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn25 S net67 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn24 pn p VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn23 net58 p net67 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn22 net56 pn net67 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn21 net56 CI VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn20 net58 net56 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn18 net18 B p VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn17 net60 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn16 net59 net60 p VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn15 net59 net18 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn14 net18 A VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ADDF_V2_1




.subckt SAEDRVT14_ADDF_V2_2 VDD VSS VBP VBN S CO A B CI
Mxmn28 net60 pn net74 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn27 net56 p net74 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn26 CO net74 VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmn25 S net67 VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmn24 pn p VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn23 net58 p net67 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn22 net56 pn net67 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn21 net56 CI VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn20 net58 net56 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn18 net18 B p VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn17 net60 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn16 net59 net60 p VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn15 net59 net18 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn14 net18 A VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmpdummy VDD A VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp26 net60 p net74 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp25 CO net74 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp24 net56 pn net74 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp23 S net67 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp22 pn p VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp21 net56 p net67 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp20 net049 pn net67 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp19 net56 CI VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp18 net049 net56 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp16 net18 net60 p VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp15 net60 B VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp14 net050 B p VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp13 net050 net18 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp12 net18 A VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ADDF_V2_2




.subckt SAEDRVT14_ADDH_0P5 VDD VSS VBP VBN S CO A B
Mxmi1#2fn2 CO i1#2fint_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi1#2fn1 i1#2fmidn_a_b B VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi1#2fn0 i1#2fint_zn A i1#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fn5 i0#2fab A VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fn4 S i0#2fint_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fi0#2fn3 i0#2fi0#2fbb i0#2fab i0#2fint_zn VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fi0#2fn2 i0#2fi0#2fbb B VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fi0#2fn1 i0#2fi0#2fbbb A i0#2fint_zn VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi1#2fp2 CO i1#2fint_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi1#2fp1 i1#2fint_zn A VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi1#2fp0 i1#2fint_zn B VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fp5 i0#2fab A VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fp4 S i0#2fint_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fi0#2fp3 i0#2fi0#2fbb A i0#2fint_zn VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fi0#2fp2 i0#2fi0#2fbb B VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fi0#2fp1 i0#2fi0#2fnet21 i0#2fab i0#2fint_zn VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ADDH_0P5




.subckt SAEDRVT14_ADDH_1 VDD VSS VBP VBN S CO A B
Mxmi1#2fn2 CO i1#2fint_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi1#2fn1 i1#2fmidn_a_b B VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi1#2fn0 i1#2fint_zn A i1#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fn5 i0#2fab A VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fn4 S i0#2fint_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fi0#2fn3 i0#2fi0#2fbb i0#2fab i0#2fint_zn VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fi0#2fn2 i0#2fi0#2fbb B VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fi0#2fn1 i0#2fi0#2fbbb A i0#2fint_zn VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi1#2fp2 CO i1#2fint_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi1#2fp1 i1#2fint_zn A VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi1#2fp0 i1#2fint_zn B VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fp5 i0#2fab A VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fp4 S i0#2fint_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fi0#2fp3 i0#2fi0#2fbb A i0#2fint_zn VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fi0#2fp2 i0#2fi0#2fbb B VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fi0#2fp1 i0#2fi0#2fnet21 i0#2fab i0#2fint_zn VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ADDH_1




.subckt SAEDRVT14_ADDH_2 VDD VSS VBP VBN S CO A B
Mxmmn0 VSS B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi1#2fn2 CO i1#2fint_zn VSS VBN n08 l=0.014u nf=2 m=2 nfin=4
Mxmi1#2fn1 i1#2fmidn_a_b B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi1#2fn0 i1#2fint_zn A i1#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn5 i0#2fab A VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fn4 S i0#2fint_zn VSS VBN n08 l=0.014u nf=2 m=2 nfin=4
Mxmi0#2fi0#2fn3 i0#2fi0#2fbb i0#2fab i0#2fint_zn VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fi0#2fn2 i0#2fi0#2fbb B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fi0#2fn1 i0#2fi0#2fbbb A i0#2fint_zn VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi1#2fp2 CO i1#2fint_zn VDD VBP p08 l=0.014u nf=2 m=2 nfin=4
Mxmi1#2fp1 i1#2fint_zn A VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi1#2fp0 i1#2fint_zn B VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp5 i0#2fab A VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fp4 S i0#2fint_zn VDD VBP p08 l=0.014u nf=2 m=2 nfin=4
Mxmi0#2fi0#2fp3 i0#2fi0#2fbb A i0#2fint_zn VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fi0#2fp2 i0#2fi0#2fbb B VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fi0#2fp1 i0#2fi0#2fnet21 i0#2fab i0#2fint_zn VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ADDH_2




.subckt SAEDRVT14_ADDH_4 VDD VSS VBP VBN S CO A B
Mxmi1#2fn11 i1#2fmidn_a_b1 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi1#2fn01 i1#2fint_zn A i1#2fmidn_a_b1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi1#2fn2 CO i1#2fint_zn VSS VBN n08 l=0.014u nf=4 m=4 nfin=4
Mxmi1#2fn1 i1#2fmidn_a_b B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi1#2fn0 i1#2fint_zn A i1#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn5 i0#2fab A VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn4 S i0#2fint_zn VSS VBN n08 l=0.014u nf=4 m=4 nfin=4
Mxmi0#2fi0#2fn3 i0#2fi0#2fbb i0#2fab i0#2fint_zn VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fi0#2fn2 i0#2fi0#2fbb B VSS VBN n08 l=0.014u nf=2 m=2 nfin=4
Mxmi0#2fi0#2fn1 i0#2fi0#2fbbb A i0#2fint_zn VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb VSS VBN n08 l=0.014u nf=2 m=2 nfin=4
Mxmi1#2fp2 CO i1#2fint_zn VDD VBP p08 l=0.014u nf=4 m=4 nfin=4
Mxmi1#2fp1 i1#2fint_zn A VDD VBP p08 l=0.014u nf=2 m=2 nfin=4
Mxmi1#2fp0 i1#2fint_zn B VDD VBP p08 l=0.014u nf=2 m=2 nfin=4
Mxmi0#2fp5 i0#2fab A VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp4 S i0#2fint_zn VDD VBP p08 l=0.014u nf=4 m=4 nfin=4
Mxmi0#2fi0#2fp3 i0#2fi0#2fbb A i0#2fint_zn VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fi0#2fp2 i0#2fi0#2fbb B VDD VBP p08 l=0.014u nf=2 m=2 nfin=4
Mxmi0#2fi0#2fp1 i0#2fi0#2fnet21 i0#2fab i0#2fint_zn VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb VDD VBP p08 l=0.014u nf=2 m=2 nfin=4
.ends SAEDRVT14_ADDH_4




.subckt SAEDRVT14_AN2_0P5 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn2 X i0#2fint_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmi0#2fn1 i0#2fmidn_a_b A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fn0 i0#2fint_zn A1 i0#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fp2 X i0#2fint_zn VDD VBP p08 l=0.014u nf=3 m=1 nfin=2
Mxmi0#2fp1 i0#2fint_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fp0 i0#2fint_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AN2_0P5




.subckt SAEDRVT14_AN2_0P75 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn2 X i0#2fint_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmi0#2fn1 i0#2fmidn_a_b A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fn0 i0#2fint_zn A1 i0#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fp2 X i0#2fint_zn VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmi0#2fp1 i0#2fint_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fp0 i0#2fint_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AN2_0P75




.subckt SAEDRVT14_AN2_1 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn2 X i0#2fint_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fn1 i0#2fmidn_a_b A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fn0 i0#2fint_zn A1 i0#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fp2 X i0#2fint_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp1 i0#2fint_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fp0 i0#2fint_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AN2_1




.subckt SAEDRVT14_AN2_2 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn2 X i0#2fint_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmi0#2fn1 i0#2fmidn_a_b A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 i0#2fint_zn A1 i0#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp2 X i0#2fint_zn VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmi0#2fp1 i0#2fint_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp0 i0#2fint_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AN2_2




.subckt SAEDRVT14_AN2_4 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn11 i0#2fmidn_a_b1 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn01 i0#2fint_zn A1 i0#2fmidn_a_b1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn2 X i0#2fint_zn VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmi0#2fn1 i0#2fmidn_a_b A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 i0#2fint_zn A1 i0#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp2 X i0#2fint_zn VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmi0#2fp1 i0#2fint_zn A1 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmi0#2fp0 i0#2fint_zn A2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_AN2_4




.subckt SAEDRVT14_AN2_8 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn2 X i0#2fint_zn VSS VBN n08 l=0.014u nf=8 m=1 nfin=3
Mxmi0#2fn1 i0#2fmidn_a_b A2 VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmi0#2fn0 i0#2fint_zn A1 i0#2fmidn_a_b VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmi0#2fp2 X i0#2fint_zn VDD VBP p08 l=0.014u nf=8 m=1 nfin=4
Mxmi0#2fp1 i0#2fint_zn A1 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmi0#2fp0 i0#2fint_zn A2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_AN2_8




.subckt SAEDRVT14_AN2B_MM_12 A B VBN VBP VDD VSS X
Mxmi0#2fn13 i0#2fmidn_a_b3 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn12 i0#2fmidn_a_b2 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn11 i0#2fmidn_a_b1 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn03 int_zn i0#2fckb i0#2fmidn_a_b3 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn02 int_zn i0#2fckb i0#2fmidn_a_b2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn01 int_zn i0#2fckb i0#2fmidn_a_b1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=12 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_a_b B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 int_zn i0#2fckb i0#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fmn2 i0#2fckb A VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=12 m=1 nfin=4
Mxmi0#2fp1 int_zn B VDD VBP p08 l=0.014u nf=4. m=1 nfin=3
Mxmi0#2fp0 int_zn i0#2fckb VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxmi0#2fmp2 i0#2fckb A VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AN2B_MM_12




.subckt SAEDRVT14_AN2B_MM_16 A B VBN VBP VDD VSS X
Mxmi0#2fn14 i0#2fmidn_a_b4 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn13 i0#2fmidn_a_b3 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn12 i0#2fmidn_a_b2 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn11 i0#2fmidn_a_b1 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn04 int_zn i0#2fckb i0#2fmidn_a_b4 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn03 int_zn i0#2fckb i0#2fmidn_a_b3 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn02 int_zn i0#2fckb i0#2fmidn_a_b2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn01 int_zn i0#2fckb i0#2fmidn_a_b1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=16 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_a_b B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 int_zn i0#2fckb i0#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fmn2 i0#2fckb A VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=16 m=1 nfin=4
Mxmi0#2fp1 int_zn B VDD VBP p08 l=0.014u nf=5 m=1 nfin=3
Mxmi0#2fp0 int_zn i0#2fckb VDD VBP p08 l=0.014u nf=5 m=1 nfin=3
Mxmi0#2fmp2 i0#2fckb A VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AN2B_MM_16




.subckt SAEDRVT14_AN2B_MM_1 A B VBN VBP VDD VSS X
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_a_b B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 int_zn i0#2fckb i0#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fmn2 i0#2fckb A VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp1 int_zn B VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp0 int_zn i0#2fckb VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fmp2 i0#2fckb A VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AN2B_MM_1




.subckt SAEDRVT14_AN2B_MM_20 A B VBN VBP VDD VSS X
Mxmi0#2fn15 i0#2fmidn_a_b5 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn14 i0#2fmidn_a_b4 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn13 i0#2fmidn_a_b3 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn12 i0#2fmidn_a_b2 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn11 i0#2fmidn_a_b1 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn05 int_zn i0#2fckb i0#2fmidn_a_b5 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn04 int_zn i0#2fckb i0#2fmidn_a_b4 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn03 int_zn i0#2fckb i0#2fmidn_a_b3 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn02 int_zn i0#2fckb i0#2fmidn_a_b2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn01 int_zn i0#2fckb i0#2fmidn_a_b1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=20 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_a_b B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 int_zn i0#2fckb i0#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fmn2 i0#2fckb A VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=20 m=1 nfin=4
Mxmi0#2fp1 int_zn B VDD VBP p08 l=0.014u nf=6 m=1 nfin=3
Mxmi0#2fp0 int_zn i0#2fckb VDD VBP p08 l=0.014u nf=6 m=1 nfin=3
Mxmi0#2fmp2 i0#2fckb A VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AN2B_MM_20




.subckt SAEDRVT14_AN2B_MM_2 A B VBN VBP VDD VSS X
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmi0#2fn1 i0#2fmidn_a_b B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 int_zn i0#2fckb i0#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fmn2 i0#2fckb A VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=6 m=1 nfin=4
Mxmi0#2fp1 int_zn B VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp0 int_zn i0#2fckb VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fmp2 i0#2fckb A VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AN2B_MM_2




.subckt SAEDRVT14_AN2B_MM_4 a b vbn vbp vdd vss x
xmi0#2fn2 x int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmi0#2fn1 i0#2fmidn_a_b b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 int_zn i0#2fckb i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn2 i0#2fckb a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 x int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fp1 int_zn b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0 int_zn i0#2fckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp2 i0#2fckb a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AN2B_MM_4




.subckt SAEDRVT14_AN2B_MM_6 A B VBN VBP VDD VSS X
Mxmi0#2fn11 i0#2fmidn_a_b1 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn01 int_zn i0#2fckb i0#2fmidn_a_b1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=6 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_a_b B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 int_zn i0#2fckb i0#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fmn2 i0#2fckb A VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=6 m=1 nfin=4
Mxmi0#2fp1 int_zn B VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmi0#2fp0 int_zn i0#2fckb VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmi0#2fmp2 i0#2fckb A VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AN2B_MM_6




.subckt SAEDRVT14_AN2B_MM_8 A B VBN VBP VDD VSS X
Mxmi0#2fn12 i0#2fmidn_a_b2 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn11 i0#2fmidn_a_b1 B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn02 int_zn i0#2fckb i0#2fmidn_a_b2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn01 int_zn i0#2fckb i0#2fmidn_a_b1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=8 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_a_b B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 int_zn i0#2fckb i0#2fmidn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fmn2 i0#2fckb A VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=8 m=1 nfin=4
Mxmi0#2fp1 int_zn B VDD VBP p08 l=0.014u nf=3 m=1 nfin=3
Mxmi0#2fp0 int_zn i0#2fckb VDD VBP p08 l=0.014u nf=3 m=1 nfin=3
Mxmi0#2fmp2 i0#2fckb A VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AN2B_MM_8




.subckt SAEDRVT14_AN2B_PMM_2 VDD VSS VDDR X A B
Mxn2 X int_zn VSS VSS n08 l=0.014u nf=2 m=2 nfin=3
Mxn1 net019 isob VSS VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxn0 int_zn B net019 VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 isob A VSS VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxp2 X int_zn VDDR VDDR p08 l=0.014u nf=2 m=2 nfin=3
Mxp1 int_zn B VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=3
Mxp0 int_zn isob VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=2
Mxmp3 isob A VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AN2B_PMM_2




.subckt SAEDRVT14_AN2B_PMM_8 VDD VSS VDDR X A B
Mxn2 X int_zn VSS VSS n08 l=0.014u nf=6 m=1 nfin=4
Mxn1 net019 isob VSS VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxn0 int_zn B net019 VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 isob A VSS VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxp2 X int_zn VDDR VDDR p08 l=0.014u nf=6 m=1 nfin=4
Mxp1 int_zn B VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=3
Mxp0 int_zn isob VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=2
Mxmp3 isob A VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AN2B_PMM_8




.subckt SAEDRVT14_AN2B_PSECO_1 VDD VSS VDDR X A B
Mxn2 X int_zn VSS VSS n08 l=0.014u nf=1 m=1 nfin=3
Mxn1 net019 isob VSS VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxn0 int_zn B net019 VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 isob A VSS VSS n08 l=0.014u nf=1 m=1 nfin=2
Mxmn2 VSS int_zn VSS VSS n08 l=0.014u nf=1 m=1 nfin=2
Mxp2 X int_zn VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=4
Mxp1 int_zn B VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=2
Mxp0 int_zn isob VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=4
Mxmp3 isob A VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=4
Mxmp2 VDDR int_zn VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AN2B_PSECO_1




.subckt SAEDRVT14_AN2B_PSECO_2 VDD VSS VDDR X A B
Mxn2 X int_zn VSS VSS n08 l=0.014u nf=2 m=1 nfin=3
Mxn1 net019 isob VSS VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxn0 int_zn B net019 VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 isob A VSS VSS n08 l=0.014u nf=1 m=1 nfin=2
Mxp2 X int_zn VDDR VDDR p08 l=0.014u nf=2 m=1 nfin=4
Mxp1 int_zn B VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=2
Mxp0 int_zn isob VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=4
Mxmp3 isob A VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AN2B_PSECO_2




.subckt SAEDRVT14_AN2B_PSECO_4 VDD VSS VDDR X A B
Mxn11 net0191 isob VSS VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxn01 int_zn B net0191 VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxn2 X int_zn VSS VSS n08 l=0.014u nf=4 m=1 nfin=3
Mxn1 net019 isob VSS VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxn0 int_zn B net019 VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 isob A VSS VSS n08 l=0.014u nf=1 m=1 nfin=2
Mxp2 X int_zn VDDR VDDR p08 l=0.014u nf=4 m=1 nfin=4
Mxp1 int_zn B VDDR VDDR p08 l=0.014u nf=2 m=1 nfin=2
Mxp0 int_zn isob VDDR VDDR p08 l=0.014u nf=2 m=1 nfin=4
Mxmp3 isob A VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AN2B_PSECO_4




.subckt SAEDRVT14_AN2B_PSECO_8 VDD VSS VDDR X A B
Mxn12 net0192 isob VSS VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxn11 net0191 isob VSS VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxn02 int_zn B net0192 VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxn01 int_zn B net0191 VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxn2 X int_zn VSS VSS n08 l=0.014u nf=8 m=1 nfin=3
Mxn1 net019 isob VSS VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxn0 int_zn B net019 VSS n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 isob A VSS VSS n08 l=0.014u nf=1 m=1 nfin=2
Mxp2 X int_zn VDDR VDDR p08 l=0.014u nf=8 m=1 nfin=4
Mxp1 int_zn B VDDR VDDR p08 l=0.014u nf=3 m=1 nfin=2
Mxp0 int_zn isob VDDR VDDR p08 l=0.014u nf=3 m=1 nfin=4
Mxmp3 isob A VDDR VDDR p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AN2B_PSECO_8




.subckt SAEDRVT14_AN2_ECO_2 VDD VSS VBP VBN X A1 A2
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmn1 midn_a_b A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=3 m=1 nfin=4
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AN2_ECO_2




.subckt SAEDRVT14_AN2_ISO_1 VDD VSS VBP VBN X CK EN
Mxn2 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxn1 midn_a_b EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxn0 int_zn CK midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxp2 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxp1 int_zn CK VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxp0 int_zn EN VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AN2_ISO_1




.subckt SAEDRVT14_AN2_ISO4_1 VDD VSS VBP VBN EN CK0 CK1 CK2 CK3 X0 X1 X2 X3
MM15 X0 int_zn_0 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
MM14 midn_a_b_0 EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
MM13 int_zn_0 CK0 midn_a_b_0 VBN n08 l=0.014u nf=1 m=1 nfin=3
MM9 X1 int_zn_1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
MM8 midn_a_b_1 EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
MM7 int_zn_1 CK1 midn_a_b_1 VBN n08 l=0.014u nf=1 m=1 nfin=3
MM2 X2 int_zn_2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
MM1 midn_a_b_2 EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
MM0 int_zn_2 CK2 midn_a_b_2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn2 X3 int_zn_3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn1 midn_a_b_3 EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn0 int_zn_3 CK3 midn_a_b_3 VBN n08 l=0.014u nf=1 m=1 nfin=3
MM18 X0 int_zn_0 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
MM17 int_zn_0 CK0 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
MM16 int_zn_0 EN VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
MM12 X1 int_zn_1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
MM11 int_zn_1 CK1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
MM10 int_zn_1 EN VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
MM5 X2 int_zn_2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
MM4 int_zn_2 CK2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
MM3 int_zn_2 EN VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxp2 X3 int_zn_3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp1 int_zn_3 CK3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxp0 int_zn_3 EN VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AN2_ISO4_1




.subckt SAEDRVT14_AN2_ISO4_4 VDD VSS VBP VBN EN CK0 CK1 CK2 CK3 X0 X1 X2 X3
MM20 midn_a_b1_0 EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
MM19 int_zn_0 CK0 midn_a_b1_0 VBN n08 l=0.014u nf=1 m=1 nfin=4
MM18 X0 int_zn_0 VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
MM17 midn_a_b_0 EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
MM16 int_zn_0 CK0 midn_a_b_0 VBN n08 l=0.014u nf=1 m=1 nfin=4
MM24 int_zn_1 CK1 midn_a_b_1 VBN n08 l=0.014u nf=1 m=1 nfin=4
MM25 midn_a_b_1 EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
MM26 X1 int_zn_1 VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
MM27 int_zn_1 CK1 midn_a_b1_1 VBN n08 l=0.014u nf=1 m=1 nfin=4
MM28 midn_a_b1_1 EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
MM38 midn_a_b_2 EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
MM39 int_zn_2 CK2 midn_a_b_2 VBN n08 l=0.014u nf=1 m=1 nfin=4
MM40 X3 int_zn_3 VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
MM41 int_zn_3 CK3 midn_a_b1_3 VBN n08 l=0.014u nf=1 m=1 nfin=4
MM42 midn_a_b1_3 EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
MM35 midn_a_b1_2 EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
MM36 int_zn_2 CK2 midn_a_b1_2 VBN n08 l=0.014u nf=1 m=1 nfin=4
MM37 X2 int_zn_2 VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
MM46 int_zn_3 CK3 midn_a_b_3 VBN n08 l=0.014u nf=1 m=1 nfin=4
MM47 midn_a_b_3 EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
MM23 X0 int_zn_0 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
MM22 int_zn_0 CK0 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
MM21 int_zn_0 EN VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
MM29 int_zn_1 EN VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
MM30 int_zn_1 CK1 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
MM31 X1 int_zn_1 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
MM32 X2 int_zn_2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
MM33 int_zn_2 CK2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
MM34 int_zn_2 EN VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
MM43 int_zn_3 EN VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
MM44 int_zn_3 CK3 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
MM45 X3 int_zn_3 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_AN2_ISO4_4




.subckt SAEDRVT14_AN2_ISO_4 VDD VSS VBP VBN X CK EN
Mxn11 midn_a_b1 EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn01 int_zn CK midn_a_b1 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn2 X int_zn VSS VBN n08 l=0.014u nf=1 m=4 nfin=4
Mxn1 midn_a_b EN VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn0 int_zn CK midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxp2 X int_zn VDD VBP p08 l=0.014u nf=1 m=4 nfin=4
Mxp1 int_zn CK VDD VBP p08 l=0.014u nf=1 m=2 nfin=3
Mxp0 int_zn EN VDD VBP p08 l=0.014u nf=1 m=2 nfin=3
.ends SAEDRVT14_AN2_ISO_4




.subckt SAEDRVT14_AN2_MM_0P5 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fn1 i0#2fmidn_en_ck A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fn0 int_zn A1 i0#2fmidn_en_ck VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AN2_MM_0P5




.subckt SAEDRVT14_AN2_MM_12 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn13 i0#2fmidn_en_ck3 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn12 i0#2fmidn_en_ck2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn11 i0#2fmidn_en_ck1 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn03 int_zn A1 i0#2fmidn_en_ck3 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn02 int_zn A1 i0#2fmidn_en_ck2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn01 int_zn A1 i0#2fmidn_en_ck1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=12 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_en_ck A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 int_zn A1 i0#2fmidn_en_ck VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=12 m=1 nfin=4
Mxmi0#2fp1 int_zn A1 VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxmi0#2fp0 int_zn A2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
.ends SAEDRVT14_AN2_MM_12




.subckt SAEDRVT14_AN2_MM_16 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn13 i0#2fmidn_en_ck3 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn12 i0#2fmidn_en_ck2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn11 i0#2fmidn_en_ck1 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn03 int_zn A1 i0#2fmidn_en_ck3 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn02 int_zn A1 i0#2fmidn_en_ck2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn01 int_zn A1 i0#2fmidn_en_ck1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=16 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_en_ck A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 int_zn A1 i0#2fmidn_en_ck VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=16 m=1 nfin=4
Mxmi0#2fp1 int_zn A1 VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxmi0#2fp0 int_zn A2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
.ends SAEDRVT14_AN2_MM_16




.subckt SAEDRVT14_AN2_MM_1 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_en_ck A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fn0 int_zn A1 i0#2fmidn_en_ck VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AN2_MM_1




.subckt SAEDRVT14_AN2_MM_20 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn14 i0#2fmidn_en_ck4 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn13 i0#2fmidn_en_ck3 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn12 i0#2fmidn_en_ck2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn11 i0#2fmidn_en_ck1 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn04 int_zn A1 i0#2fmidn_en_ck4 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn03 int_zn A1 i0#2fmidn_en_ck3 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn02 int_zn A1 i0#2fmidn_en_ck2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn01 int_zn A1 i0#2fmidn_en_ck1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=20 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_en_ck A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 int_zn A1 i0#2fmidn_en_ck VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=20 m=1 nfin=4
Mxmi0#2fp1 int_zn A1 VDD VBP p08 l=0.014u nf=5 m=1 nfin=3
Mxmi0#2fp0 int_zn A2 VDD VBP p08 l=0.014u nf=5 m=1 nfin=3
.ends SAEDRVT14_AN2_MM_20




.subckt SAEDRVT14_AN2_MM_2 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_en_ck A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fn0 int_zn A1 i0#2fmidn_en_ck VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmi0#2fp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AN2_MM_2




.subckt SAEDRVT14_AN2_MM_3 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=3 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_en_ck A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 int_zn A1 i0#2fmidn_en_ck VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=3 m=1 nfin=4
Mxmi0#2fp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AN2_MM_3




.subckt SAEDRVT14_AN2_MM_4 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn11 i0#2fmidn_en_ck1 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fn01 int_zn A1 i0#2fmidn_en_ck1 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_en_ck A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fn0 int_zn A1 i0#2fmidn_en_ck VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmi0#2fp1 int_zn A1 VDD VBP p08 l=0.014u nf=2 m=1 nfin=2
Mxmi0#2fp0 int_zn A2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_AN2_MM_4




.subckt SAEDRVT14_AN2_MM_6 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn11 i0#2fmidn_en_ck1 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn01 int_zn A1 i0#2fmidn_en_ck1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=6 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_en_ck A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 int_zn A1 i0#2fmidn_en_ck VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=6 m=1 nfin=4
Mxmi0#2fp1 int_zn A1 VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmi0#2fp0 int_zn A2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_AN2_MM_6




.subckt SAEDRVT14_AN2_MM_8 VDD VSS VBP VBN X A1 A2
Mxmi0#2fn12 i0#2fmidn_en_ck2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn11 i0#2fmidn_en_ck1 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn02 int_zn A1 i0#2fmidn_en_ck2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn01 int_zn A1 i0#2fmidn_en_ck1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn2 X int_zn VSS VBN n08 l=0.014u nf=8 m=1 nfin=4
Mxmi0#2fn1 i0#2fmidn_en_ck A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn0 int_zn A1 i0#2fmidn_en_ck VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp2 X int_zn VDD VBP p08 l=0.014u nf=8 m=1 nfin=4
Mxmi0#2fp1 int_zn A1 VDD VBP p08 l=0.014u nf=3 m=1 nfin=3
Mxmi0#2fp0 int_zn A2 VDD VBP p08 l=0.014u nf=3 m=1 nfin=3
.ends SAEDRVT14_AN2_MM_8




.subckt SAEDRVT14_AN3_0P5 VDD VSS VBP VBN X A1 A2 A3
Mxmn3 midn_b_c A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn1 midn_a_b A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmp3 int_zn A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AN3_0P5




.subckt SAEDRVT14_AN3_0P75 VDD VSS VBP VBN X A1 A2 A3
Mxmn3 midn_b_c A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn1 midn_a_b A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp3 int_zn A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AN3_0P75




.subckt SAEDRVT14_AN3_1 VDD VSS VBP VBN X A1 A2 A3
Mxmn3 midn_b_c A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn1 midn_a_b A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp3 int_zn A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AN3_1




.subckt SAEDRVT14_AN3_2 VDD VSS VBP VBN X A1 A2 A3
Mxmn3 midn_b_c A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn1 midn_a_b A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp3 int_zn A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AN3_2




.subckt SAEDRVT14_AN3_4 VDD VSS VBP VBN X A1 A2 A3
Mxmn31 midn_b_c1 A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn11 midn_a_b A2 midn_b_c1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 midn_b_c A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmn1 midn_a_b A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmp3 int_zn A3 VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=2 m=1 nfin=2
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_AN3_4




.subckt SAEDRVT14_AN3_8 VDD VSS VBP VBN X A1 A2 A3
Mxmn33 midn_b_c3 A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn32 midn_b_c2 A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn31 midn_b_c1 A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn13 midn_a_b A2 midn_b_c3 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn12 midn_a_b A2 midn_b_c2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn11 midn_a_b A2 midn_b_c1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 midn_b_c A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=8 m=1 nfin=3
Mxmn1 midn_a_b A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=4 m=1 nfin=2
Mxmp3 int_zn A3 VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=8 m=1 nfin=4
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=4 m=1 nfin=2
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
.ends SAEDRVT14_AN3_8




.subckt SAEDRVT14_AN3_ECO_1 VDD VSS VBP VBN X A1 A2 A3
Mxmn3 midn_b_c A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn1 midn_a_b A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp3 int_zn A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AN3_ECO_1




.subckt SAEDRVT14_AN4_0P5 VDD VSS VBP VBN X A1 A2 A3 A4
Mxmn4 midn_c_d A4 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn3 midn_b_c A3 midn_c_d VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn1 midn_a_b A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmp4 int_zn A4 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp3 int_zn A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AN4_0P5




.subckt SAEDRVT14_AN4_0P75 VDD VSS VBP VBN X A1 A2 A3 A4
Mxmn4 midn_c_d A4 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 midn_b_c A3 midn_c_d VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn1 midn_a_b A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp4 int_zn A4 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp3 int_zn A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AN4_0P75




.subckt SAEDRVT14_AN4_1 VDD VSS VBP VBN X A1 A2 A3 A4
Mxmn4 midn_c_d A4 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn3 midn_b_c A3 midn_c_d VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn1 midn_a_b A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmp4 int_zn A4 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp3 int_zn A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AN4_1




.subckt SAEDRVT14_AN4_2 VDD VSS VBP VBN X A1 A2 A3 A4
Mxmn4 midn_c_d A4 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 midn_b_c A3 midn_c_d VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn1 midn_a_b A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp4 int_zn A4 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp3 int_zn A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AN4_2




.subckt SAEDRVT14_AN4_4 VDD VSS VBP VBN X A1 A2 A3 A4
Mxmn41 midn_c_d1 A4 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn31 midn_b_c A3 midn_c_d1 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn11 midn_a_b1 A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn01 int_zn A1 midn_a_b1 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn4 midn_c_d A4 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn3 midn_b_c A3 midn_c_d VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmn1 midn_a_b A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmp4 int_zn A4 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp3 int_zn A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AN4_4




.subckt SAEDRVT14_AN4_8 VDD VSS VBP VBN X A1 A2 A3 A4
Mxmn43 midn_c_d3 A4 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn42 midn_c_d2 A4 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn41 midn_c_d1 A4 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn33 midn_b_c A3 midn_c_d3 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn32 midn_b_c A3 midn_c_d2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn31 midn_b_c A3 midn_c_d1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn13 midn_a_b3 A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn12 midn_a_b2 A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn11 midn_a_b1 A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn03 int_zn A1 midn_a_b3 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn02 int_zn A1 midn_a_b2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn01 int_zn A1 midn_a_b1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn4 midn_c_d A4 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 midn_b_c A3 midn_c_d VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=8 m=1 nfin=4
Mxmn1 midn_a_b A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp4 int_zn A4 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp3 int_zn A3 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=8 m=1 nfin=4
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_AN4_8




.subckt SAEDRVT14_AN4_ECO_2 VDD VSS VBP VBN X A1 A2 A3 A4
Mxmn4 midn_c_d A4 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 midn_b_c A3 midn_c_d VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn2 X int_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmn1 midn_a_b A2 midn_b_c VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 int_zn A1 midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp4 int_zn A4 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp3 int_zn A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp2 X int_zn VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp1 int_zn A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 int_zn A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AN4_ECO_2




.subckt SAEDRVT14_AO211_1 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmn7 midn_a1_a2 A2 VSS VBN n08 l=0.014u nf=3 m=1 nfin=3
Mxmn6 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn5 int_zn A1 midn_a1_a2 VBN n08 l=0.014u nf=3 m=1 nfin=3
Mxmn4 int_zn B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn3 int_zn B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmp5 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp4 VDD A2 midp_a1a2_b VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp2 midp_b_c B2 int_zn VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp1 VDD A1 midp_a1a2_b VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 midp_a1a2_b B1 midp_b_c VBP p08 l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_AO211_1




.subckt SAEDRVT14_AO211_2 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmn7 midn_a1_a2 A2 VSS VBN n08 l=0.014u nf=3 m=1 nfin=3
Mxmn6 X int_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmn5 int_zn A1 midn_a1_a2 VBN n08 l=0.014u nf=3 m=1 nfin=3
Mxmn4 int_zn B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn3 int_zn B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmp5 X int_zn VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp4 VDD A2 midp_a1a2_b VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp2 midp_b_c B2 int_zn VBP p08 l=0.014u nf=3 m=1 nfin=3
Mxmp1 VDD A1 midp_a1a2_b VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 midp_a1a2_b B1 midp_b_c VBP p08 l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_AO211_2




.subckt SAEDRVT14_AO211_4 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmn71 midn_a1_a21 A2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn51 int_zn A1 midn_a1_a21 VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn7 midn_a1_a2 A2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn6 X int_zn VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmn5 int_zn A1 midn_a1_a2 VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn4 int_zn B1 VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmn3 int_zn B2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmp21 midp_b_c1 B2 int_zn VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp01 midp_a1a2_b B1 midp_b_c1 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp5 X int_zn VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp4 VDD A2 midp_a1a2_b VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp2 midp_b_c B2 int_zn VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 VDD A1 midp_a1a2_b VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp0 midp_a1a2_b B1 midp_b_c VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AO211_4




.subckt SAEDRVT14_AO21_1 VDD VSS VBP VBN X A1 A2 B
Mxmn5 midn_a1_a2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn4 int_zn A1 midn_a1_a2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn3 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 int_zn B VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmp4 VDD A2 midp_a1a2_b VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp3 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 VDD A1 midp_a1a2_b VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 midp_a1a2_b B int_zn VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AO21_1




.subckt SAEDRVT14_AO211_U_0P5 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmn7 midn_a1_a2 A2 VSS VBN n08 l=0.014u nf=4 m=1 nfin=2
Mxmn6 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn5 int_zn A1 midn_a1_a2 VBN n08 l=0.014u nf=3 m=1 nfin=2
Mxmn4 int_zn B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn3 int_zn B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp5 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp4 VDD A2 midp_a1a2_b VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp2 midp_b_c B2 int_zn VBP p08 l=0.014u nf=2 m=1 nfin=2
Mxmp1 VDD A1 midp_a1a2_b VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 midp_a1a2_b B1 midp_b_c VBP p08 l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_AO211_U_0P5




.subckt SAEDRVT14_AO21_2 vdd vss vbp vbn x a1 a2 b
xmn5 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn4 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn3 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn0 int_zn b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp4 vdd a2 midp_a1a2_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 vdd a1 midp_a1a2_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_a1a2_b b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AO21_2




.subckt SAEDRVT14_AO21_4 VDD VSS VBP VBN X A1 A2 B
Mxmn51 midn_a1_a21 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn41 int_zn A1 midn_a1_a21 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn5 midn_a1_a2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn4 int_zn A1 midn_a1_a2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn3 X int_zn VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmn0 int_zn B VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmp4 VDD A2 midp_a1a2_b VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp3 X int_zn VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp1 VDD A1 midp_a1a2_b VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp0 midp_a1a2_b B int_zn VBP p08 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_AO21_4




.subckt SAEDRVT14_AO21B_0P5 VDD VSS VBP VBN X A1 A2 B
Mxmn4 X B midn_a_b1nrb2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn3 midn_a_b1nrb2 b1nrb2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn1 b1nrb2 A1 midn_b1_b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 midn_b1_b2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp4 X b1nrb2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp3 X B VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp1 b1nrb2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 b1nrb2 A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO21B_0P5




.subckt SAEDRVT14_AO21B_1 VDD VSS VBP VBN X A1 A2 B
Mxmnbuf2 X d1g2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmnbuf1 d1g2 x1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn4 x1 B midn_a_b1nrb2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 midn_a_b1nrb2 b1nrb2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn1 b1nrb2 A1 midn_b1_b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 midn_b1_b2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmpbuf2 X d1g2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmpbuf1 d1g2 x1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp4 x1 b1nrb2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp3 x1 B VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp1 b1nrb2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 b1nrb2 A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AO21B_1




.subckt SAEDRVT14_AO21B_2 VDD VSS VBP VBN X A1 A2 B
Mxmnbuf2 X d1g2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmnbuf1 d1g2 x1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn41 x1 B midn_a_b1nrb21 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn31 midn_a_b1nrb21 b1nrb2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn4 x1 B midn_a_b1nrb2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 midn_a_b1nrb2 b1nrb2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn1 b1nrb2 A1 midn_b1_b2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 midn_b1_b2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmpbuf2 X d1g2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmpbuf1 d1g2 x1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp4 x1 b1nrb2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp3 x1 B VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp1 b1nrb2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp0 b1nrb2 A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AO21B_2




.subckt SAEDRVT14_AO21B_4 VDD VSS VBP VBN X A1 A2 B
Mxmnbuf2 X d1g2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmnbuf1 d1g2 x1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn43 x1 B midn_a_b1nrb2_3 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn42 x1 B midn_a_b1nrb2_2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn41 x1 B midn_a_b1nrb2_1 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn33 midn_a_b1nrb2_3 b1nrb2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn32 midn_a_b1nrb2_2 b1nrb2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn31 midn_a_b1nrb2_1 b1nrb2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn4 x1 B midn_a_b1nrb2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 midn_a_b1nrb2 b1nrb2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn1 b1nrb2 A1 midn_b1_b2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 midn_b1_b2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmpbuf2 X d1g2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmpbuf1 d1g2 x1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp4 x1 b1nrb2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp3 x1 B VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp1 b1nrb2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp0 b1nrb2 A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AO21B_4




.subckt SAEDRVT14_AO21_ECO_1 VDD VSS VBP VBN X A1 A2 B
Mxmn5 midn_a1_a2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn4 int_zn A1 midn_a1_a2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 int_zn B VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp4 int_zn A2 midp_a1a2_b VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp3 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 int_zn A1 midp_a1a2_b VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp0 midp_a1a2_b B VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AO21_ECO_1




.subckt SAEDRVT14_AO21_U_0P5 vdd vss vbp vbn x a1 a2 b
xmn5 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 int_zn b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 vdd a2 midp_a1a2_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 vdd a1 midp_a1a2_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 midp_a1a2_b b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO21_U_0P5




.subckt SAEDRVT14_AO22_0P5 vdd vss vbp vbn x a1 a2 b1 b2
xmn8 int_zn b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn7 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn6 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp7 int_zn a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 int_zn a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 midp_a1a2_b1b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 midp_a1a2_b1b2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AO22_0P5




.subckt SAEDRVT14_AO22_0P75 vdd vss vbp vbn x a1 a2 b1 b2
xmn8 int_zn b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn7 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn6 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp7 int_zn a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 int_zn a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 midp_a1a2_b1b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 midp_a1a2_b1b2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AO22_0P75




.subckt SAEDRVT14_AO221_0P5 vdd vss vbp vbn x a1 a2 b1 b2 c
xmn10 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn9 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn8 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn7 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn6 int_zn b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 int_zn c vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp9 midp_a1a2_b1b2 b2 midp_b1b2_c vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp8 vdd a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp7 vdd a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp6 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 midp_a1a2_b1b2 b1 midp_b1b2_c vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_b1b2_c c int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AO221_0P5




.subckt SAEDRVT14_AO221_1 vdd vss vbp vbn x a1 a2 b1 b2 c
xmn10 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn9 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn8 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn7 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn6 int_zn b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn3 int_zn c vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp9 midp_a1a2_b1b2 b2 midp_b1b2_c vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp8 vdd a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp7 vdd a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp6 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 midp_a1a2_b1b2 b1 midp_b1b2_c vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_b1b2_c c int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AO221_1




.subckt SAEDRVT14_AO221_2 vdd vss vbp vbn x a1 a2 b1 b2 c
xmn10 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=2 nfin=2
xmn9 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=2 nfin=3
xmn8 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=2 nfin=3
xmn7 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn6 int_zn b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=2 nfin=3
xmn3 int_zn c vss vbn n08_rev l=0.014u nf=1 m=2 nfin=3
xmp9 midp_a1a2_b1b2 b2 midp_b1b2_c vbp p08_rev l=0.014u nf=1 m=2 nfin=3
xmp8 vdd a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=2 nfin=3
xmp7 vdd a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=2 nfin=3
xmp6 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp1 midp_a1a2_b1b2 b1 midp_b1b2_c vbp p08_rev l=0.014u nf=1 m=2 nfin=3
xmp0 midp_b1b2_c c int_zn vbp p08_rev l=0.014u nf=1 m=2 nfin=3
.ends SAEDRVT14_AO221_2




.subckt SAEDRVT14_AO221_4 vdd vss vbp vbn x a1 a2 b1 b2 c
xmn101 int_zn a1 midn_a1_a21 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn91 midn_a1_a21 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn81 midn_b1_b21 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn61 int_zn b1 midn_b1_b21 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn10 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn9 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn8 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn7 x int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn6 int_zn b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 int_zn c vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp6_3 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp6_2 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp6_1 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp9 midp_a1a2_b1b2 b2 midp_b1b2_c vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp8 vdd a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp7 vdd a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp6 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 midp_a1a2_b1b2 b1 midp_b1b2_c vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp0 midp_b1b2_c c int_zn vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_AO221_4




.subckt SAEDRVT14_AO22_1 vdd vss vbp vbn x a1 a2 b1 b2
xmn8 int_zn b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn7 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn6 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp7 int_zn a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 int_zn a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 midp_a1a2_b1b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 midp_a1a2_b1b2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AO22_1




.subckt SAEDRVT14_AO222_1 vdd vss vbp vbn x a1 a2 b1 b2 c1 c2
xmn13 midn_c1_c2 c2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 int_zn c1 midn_c1_c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn11 int_zn b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn10 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn9 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn8 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn6 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp13 midp_b1b2_c1c2 c2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp12 midp_a1a2_b1b2 b2 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp11 int_zn a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp10 int_zn a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp9 midp_a1a2_b1b2 b1 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp8 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_b1b2_c1c2 c1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AO222_1




.subckt SAEDRVT14_AO222_2 vdd vss vbp vbn x a1 a2 b1 b2 c1 c2
xmn13 midn_c1_c2 c2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn12 int_zn c1 midn_c1_c2 vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn11 int_zn b1 midn_b1_b2 vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn10 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn9 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn8 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn6 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp13 midp_b1b2_c1c2 c2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp12 midp_a1a2_b1b2 b2 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp11 int_zn a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp10 int_zn a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp9 midp_a1a2_b1b2 b1 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp8 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 midp_b1b2_c1c2 c1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_AO222_2




.subckt SAEDRVT14_AO222_4 vdd vss vbp vbn x a1 a2 b1 b2 c1 c2
xmn13 midn_c1_c2 c2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn12 int_zn c1 midn_c1_c2 vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmn11 int_zn b1 midn_b1_b2 vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn10 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn9 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmn8 x int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn6 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmp13 midp_b1b2_c1c2 c2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp12 midp_a1a2_b1b2 b2 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp11 int_zn a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmp10 int_zn a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmp9 midp_a1a2_b1b2 b1 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp8 x int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 midp_b1b2_c1c2 c1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_AO222_4




.subckt SAEDRVT14_AO22_2 vdd vss vbp vbn x a1 a2 b1 b2
xmn8 int_zn b1 midn_b1_b2 vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn7 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn6 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp7 int_zn a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp6 int_zn a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp5 midp_a1a2_b1b2 b2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp4 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a1a2_b1b2 b1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_AO22_2




.subckt SAEDRVT14_AO222_U_0P5 vdd vss vbp vbn x a1 a2 b1 b2 c1 c2
xmn13 midn_c1_c2 c2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 int_zn c1 midn_c1_c2 vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn11 int_zn b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn10 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn9 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn8 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn6 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp13 midp_b1b2_c1c2 c2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp12 midp_a1a2_b1b2 b2 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp11 int_zn a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp10 int_zn a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp9 midp_a1a2_b1b2 b1 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp8 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_b1b2_c1c2 c1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AO222_U_0P5




.subckt SAEDRVT14_AO22_4 vdd vss vbp vbn x a1 a2 b1 b2
xmn8 int_zn b1 midn_b1_b2 vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn7 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn6 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn5 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn4 int_zn a1 midn_a1_a2 vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp7 int_zn a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp6 int_zn a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp5 midp_a1a2_b1b2 b2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp4 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 midp_a1a2_b1b2 b1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
.ends SAEDRVT14_AO22_4




.subckt SAEDRVT14_AO2BB2_0P5 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 x1 a2 midn_a1a2_b1nrb2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x1 a1 midn_a1a2_b1nrb2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 midn_a1a2_b1nrb2 b1nrb2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 b1nrb2 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 midp_b1_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 x1 b1nrb2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 b1nrb2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 b1nrb2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO2BB2_0P5




.subckt SAEDRVT14_AO2BB2_1 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 x1 a2 midn_a1a2_b1nrb2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x1 a1 midn_a1a2_b1nrb2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 midn_a1a2_b1nrb2 b1nrb2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 b1nrb2 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 midp_b1_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 x1 b1nrb2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 b1nrb2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 b1nrb2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO2BB2_1




.subckt SAEDRVT14_AO2BB2_2 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 x1 a2 midn_a1a2_b1nrb2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x1 a1 midn_a1a2_b1nrb2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 midn_a1a2_b1nrb2 b1nrb2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 b1nrb2 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 midp_b1_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 x1 b1nrb2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 b1nrb2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 b1nrb2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO2BB2_2




.subckt SAEDRVT14_AO2BB2_4 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 x1 a2 midn_a1a2_b1nrb2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x1 a1 midn_a1a2_b1nrb2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 midn_a1a2_b1nrb2 b1nrb2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 b1nrb2 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 midp_b1_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 x1 b1nrb2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 b1nrb2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 b1nrb2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO2BB2_4




.subckt SAEDRVT14_AO2BB2_V1_0P5 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 net13 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 net13 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x1 net17 net13 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 net19 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 net17 b1 net19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 net17 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 net17 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 x1 a1 net18 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 net18 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO2BB2_V1_0P5




.subckt SAEDRVT14_AO2BB2_V1_0P75 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 net13 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 net13 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x1 net17 net13 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 net19 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 net17 b1 net19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 net17 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 net17 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 x1 a1 net18 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 net18 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO2BB2_V1_0P75




.subckt SAEDRVT14_AO2BB2_V1_1 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 net13 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 net13 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x1 net17 net13 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 net19 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 net17 b1 net19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 net17 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 net17 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 x1 a1 net18 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 net18 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO2BB2_V1_1




.subckt SAEDRVT14_AO2BB2_V1_2 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 net13 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 net13 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x1 net17 net13 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 net19 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 net17 b1 net19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 net17 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 net17 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 x1 a1 net18 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 net18 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO2BB2_V1_2




.subckt SAEDRVT14_AO2BB2_V1_4 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 net13 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 net13 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x1 net17 net13 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 net19 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 net17 b1 net19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 net17 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 net17 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 x1 a1 net18 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 net18 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO2BB2_V1_4




.subckt SAEDRVT14_AO31_1 vdd vss vbp vbn x a1 a2 a3 b
xmn7 midn_a2_a3 a3 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn6 net8 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 x net8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn4 midn_a1_a2 a2 midn_a2_a3 vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn1 net8 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp6 int_zn a3 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp5 int_zn a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 int_zn a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 net8 b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AO31_1




.subckt SAEDRVT14_AO31_2 vdd vss vbp vbn x a1 a2 a3 b
xmn7 midn_a2_a3 a3 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmn6 net8 b vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn5 x net8 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn4 midn_a1_a2 a2 midn_a2_a3 vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn1 net8 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp6 int_zn a3 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 int_zn a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp4 x net8 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 int_zn a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp0 net8 b int_zn vbp p08_rev l=0.014u nf=5 m=1 nfin=2
.ends SAEDRVT14_AO31_2




.subckt SAEDRVT14_AO31_4 vdd vss vbp vbn x a1 a2 a3 b
xmn41 midn_a1_a21 a2 midn_a2_a3 vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn11 net8 a1 midn_a1_a21 vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn7 midn_a2_a3 a3 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn6 net8 b vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmn5 x net8 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=3
xmn4 midn_a1_a2 a2 midn_a2_a3 vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn1 net8 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp6 int_zn a3 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp5 int_zn a2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp4 x net8 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmp1 int_zn a1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp0 net8 b int_zn vbp p08_rev l=0.014u nf=5 m=1 nfin=4
.ends SAEDRVT14_AO31_4




.subckt SAEDRVT14_AO31_U_0P5 vdd vss vbp vbn x a1 a2 a3 b
xmn7 midn_a2_a3 a3 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn6 net8 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 x net8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn4 midn_a1_a2 a2 midn_a2_a3 vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 net8 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmp6 int_zn a3 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp5 int_zn a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp4 x net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 int_zn a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 net8 b int_zn vbp p08_rev l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_AO31_U_0P5




.subckt SAEDRVT14_AO32_1 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmn10 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn9 midn_a1_a2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn8 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn7 int_zn a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn6 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 int_zn b1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp9 int_zn b1 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp8 int_zn b2 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp7 midp_a1a2_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 midp_a1a2_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a1a2_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO32_1




.subckt SAEDRVT14_AO32_2 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmn10 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn9 midn_a1_a2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn8 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn7 int_zn a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn6 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn4 int_zn b1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp9 int_zn b1 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp8 int_zn b2 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp7 midp_a1a2_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 midp_a1a2_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 midp_a1a2_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO32_2




.subckt SAEDRVT14_AO32_4 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn9 midn_a1_a2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn8 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn7 int_zn a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn6 x1 int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 int_zn b1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp9 int_zn b1 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp8 int_zn b2 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp7 midp_a1a2_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 midp_a1a2_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 x1 int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a1a2_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO32_4




.subckt SAEDRVT14_AO32_U_0P5 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmn10 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn9 midn_a1_a2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn8 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn7 int_zn a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn6 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 int_zn b1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp9 int_zn b1 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp8 int_zn b2 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp7 midp_a1a2_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 midp_a1a2_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 midp_a1a2_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO32_U_0P5




.subckt SAEDRVT14_AO33_1 vdd vss vbp vbn x a1 a2 a3 b1 b2 b3
xn12 int_zn b1 midn_b1_b2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn11 midn_b1_b2 b2 midn_b2_b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn10 midn_b2_b3 b3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn9 midn_a2_a3 a3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn8 midn_a1_a2 a2 midn_a2_a3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn7 x int_zn vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn4 int_zn a1 midn_a1_a2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp11 midp_a1a2a3_b1b2b3 b2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp10 midp_a1a2a3_b1b2b3 b3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp9 int_zn a3 midp_a1a2a3_b1b2b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp8 int_zn a2 midp_a1a2a3_b1b2b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp7 int_zn a1 midp_a1a2a3_b1b2b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp6 x int_zn vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 midp_a1a2a3_b1b2b3 b1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO33_1




.subckt SAEDRVT14_AO33_2 vdd vss vbp vbn x a1 a2 a3 b1 b2 b3
xn12 int_zn b1 midn_b1_b2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn11 midn_b1_b2 b2 midn_b2_b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn10 midn_b2_b3 b3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn9 midn_a2_a3 a3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn8 midn_a1_a2 a2 midn_a2_a3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn7 x int_zn vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn4 int_zn a1 midn_a1_a2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp11 midp_a1a2a3_b1b2b3 b2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp10 midp_a1a2a3_b1b2b3 b3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp9 int_zn a3 midp_a1a2a3_b1b2b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp8 int_zn a2 midp_a1a2a3_b1b2b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp7 int_zn a1 midp_a1a2a3_b1b2b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp6 x int_zn vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp1 midp_a1a2a3_b1b2b3 b1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO33_2




.subckt SAEDRVT14_AO33_4 vdd vss vbp vbn x a1 a2 a3 b1 b2 b3
xn12 int_zn b1 midn_b1_b2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn11 midn_b1_b2 b2 midn_b2_b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn10 midn_b2_b3 b3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn9 midn_a2_a3 a3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn8 midn_a1_a2 a2 midn_a2_a3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn7 x int_zn vss vbn n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 int_zn a1 midn_a1_a2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp11 midp_a1a2a3_b1b2b3 b2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp10 midp_a1a2a3_b1b2b3 b3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp9 int_zn a3 midp_a1a2a3_b1b2b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp8 int_zn a2 midp_a1a2a3_b1b2b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp7 int_zn a1 midp_a1a2a3_b1b2b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp6 x int_zn vdd vbp p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp1 midp_a1a2a3_b1b2b3 b1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO33_4




.subckt SAEDRVT14_AO33_U_0P5 vdd vss vbp vbn x a1 a2 a3 b1 b2 b3
xn12 int_zn b1 midn_b1_b2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn11 midn_b1_b2 b2 midn_b2_b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn10 midn_b2_b3 b3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn9 midn_a2_a3 a3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn8 midn_a1_a2 a2 midn_a2_a3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn7 x int_zn vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn4 int_zn a1 midn_a1_a2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp11 midp_a1a2a3_b1b2b3 b2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp10 midp_a1a2a3_b1b2b3 b3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp9 int_zn a3 midp_a1a2a3_b1b2b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp8 int_zn a2 midp_a1a2a3_b1b2b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp7 int_zn a1 midp_a1a2a3_b1b2b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp6 x int_zn vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 midp_a1a2a3_b1b2b3 b1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AO33_U_0P5




.subckt SAEDRVT14_AOBUF_IW_0P75 vdd vss x a vddr
xmn1 x int_zn vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 int_zn a vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x int_zn vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 int_zn a vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOBUF_IW_0P75




.subckt SAEDRVT14_AOBUF_IW_1P5 vdd vss x a vddr
xmn1 x int_zn vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 int_zn a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x int_zn vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 int_zn a vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOBUF_IW_1P5




.subckt SAEDRVT14_AOBUF_IW_3 vdd vss x a vddr
xmn1 x int_zn vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 int_zn a vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x int_zn vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 int_zn a vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOBUF_IW_3




.subckt SAEDRVT14_AOBUF_IW_6 vdd vss x a vddr
xmn1 x int_zn vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 int_zn a vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x int_zn vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 int_zn a vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOBUF_IW_6




.subckt SAEDRVT14_AOELVLUNOR_V2_10 a en vddi vdd vddr vss x
xm9 x net40 vss vss n08_rev l=0.014u nf=5 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=2
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddr vddr p08_rev l=0.014u nf=5 m=1 nfin=4
xm6 net40 net36 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddi vddi p08_rev l=0.014u nf=2 m=1 nfin=4
xm4 net36 en net17 vddi p08_rev l=0.014u nf=3 m=1 nfin=4
xm3 net17 net27 vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOELVLUNOR_V2_10




.subckt SAEDRVT14_AOELVLUNOR_V2_12 a en vddi vdd vddr vss x
xm9 x net40 vss vss n08_rev l=0.014u nf=6 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=2
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddr vddr p08_rev l=0.014u nf=6 m=1 nfin=4
xm6 net40 net36 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddi vddi p08_rev l=0.014u nf=2 m=1 nfin=4
xm4 net36 en net17 vddi p08_rev l=0.014u nf=3 m=1 nfin=4
xm3 net17 net27 vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOELVLUNOR_V2_12




.subckt SAEDRVT14_AOELVLUNOR_V2_1 a en vddi vdd vddr vss x
xm9 x net40 vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=3
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=3
xm6 net40 net36 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddi vddi p08_rev l=0.014u nf=2 m=1 nfin=3
xm4 net36 en net17 vddi p08_rev l=0.014u nf=3 m=1 nfin=3
xm3 net17 net27 vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOELVLUNOR_V2_1




.subckt SAEDRVT14_AOELVLUNOR_V2_2 a en vddi vdd vddr vss x
xm9 x net40 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=2
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm6 net40 net36 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddi vddi p08_rev l=0.014u nf=2 m=1 nfin=4
xm4 net36 en net17 vddi p08_rev l=0.014u nf=3 m=1 nfin=4
xm3 net17 net27 vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOELVLUNOR_V2_2




.subckt SAEDRVT14_AOELVLUNOR_V2_3 a en vddi vdd vddr vss x
xm9 x net40 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=2
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=3
xm6 net40 net36 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddi vddi p08_rev l=0.014u nf=2 m=1 nfin=4
xm4 net36 en net17 vddi p08_rev l=0.014u nf=3 m=1 nfin=4
xm3 net17 net27 vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOELVLUNOR_V2_3




.subckt SAEDRVT14_AOELVLUNOR_V2_4 a en vddi vdd vddr vss x
xm9 x net40 vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=2
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddr vddr p08_rev l=0.014u nf=3 m=1 nfin=3
xm6 net40 net36 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddi vddi p08_rev l=0.014u nf=2 m=1 nfin=4
xm4 net36 en net17 vddi p08_rev l=0.014u nf=3 m=1 nfin=4
xm3 net17 net27 vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOELVLUNOR_V2_4




.subckt SAEDRVT14_AOELVLUNOR_V2_6 a en vddi vdd vddr vss x
xm9 x net40 vss vss n08_rev l=0.014u nf=3 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=2
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddr vddr p08_rev l=0.014u nf=3 m=1 nfin=4
xm6 net40 net36 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddi vddi p08_rev l=0.014u nf=2 m=1 nfin=4
xm4 net36 en net17 vddi p08_rev l=0.014u nf=3 m=1 nfin=4
xm3 net17 net27 vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOELVLUNOR_V2_6




.subckt SAEDRVT14_AOELVLUNOR_V2_8 a en vddi vdd vddr vss x
xm9 x net40 vss vss n08_rev l=0.014u nf=4 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=2
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddr vddr p08_rev l=0.014u nf=4 m=1 nfin=4
xm6 net40 net36 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddi vddi p08_rev l=0.014u nf=2 m=1 nfin=4
xm4 net36 en net17 vddi p08_rev l=0.014u nf=3 m=1 nfin=4
xm3 net17 net27 vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOELVLUNOR_V2_8




.subckt SAEDRVT14_AOI21_0P5 vdd vss vbp vbn x a1 a2 b
xmn2 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 x b midp_a_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b1b2 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_a_b1b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOI21_0P5




.subckt SAEDRVT14_AOI21_0P75 vdd vss vbp vbn x a1 a2 b
xmn2 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 x b midp_a_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_a_b1b2 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_a_b1b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI21_0P75




.subckt SAEDRVT14_AOI211_0P5 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x1 b1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 midn_c1_c2 a2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmn1 x1 a1 midn_c1_c2 vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmn0 x1 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_a_b b2 midp_b_c1c2 vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp2 x1 b1 midp_a_b vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp1 midp_b_c1c2 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 midp_b_c1c2 a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_AOI211_0P5




.subckt SAEDRVT14_AOI211_1 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x1 b1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 midn_c1_c2 a2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn1 x1 a1 midn_c1_c2 vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn0 x1 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_a_b b2 midp_b_c1c2 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp2 x1 b1 midp_a_b vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 midp_b_c1c2 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_b_c1c2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI211_1




.subckt SAEDRVT14_AOI211_2 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2_2 midn_c1_c2_2 a2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn1_2 x1 a1 midn_c1_c2_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 x1 b1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 midn_c1_c2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 a1 midn_c1_c2 vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn0 x1 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3_2 midp_a_b_2 b2 midp_b_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2_2 x1 b1 midp_a_b_2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 midp_a_b b2 midp_b_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 b1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_b_c1c2 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_b_c1c2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI211_2




.subckt SAEDRVT14_AOI211_4 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2_4 midn_c1_c2_4 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2_3 midn_c1_c2_3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2_2 midn_c1_c2_2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1_4 x1 a1 midn_c1_c2_4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1_3 x1 a1 midn_c1_c2_3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1_2 x1 a1 midn_c1_c2_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 x1 b1 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn2 midn_c1_c2 a2 vss vbn n08_rev l=0.014u nf=7 m=1 nfin=4
xmn1 x1 a1 midn_c1_c2 vbn n08_rev l=0.014u nf=7 m=1 nfin=4
xmn0 x1 b2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3_4 midp_a_b_4 b2 midp_b_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3_3 midp_a_b_3 b2 midp_b_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3_2 midp_a_b_2 b2 midp_b_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2_4 x1 b1 midp_a_b_4 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2_3 x1 b1 midp_a_b_3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2_2 x1 b1 midp_a_b_2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 midp_a_b b2 midp_b_c1c2 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp2 x1 b1 midp_a_b vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 midp_b_c1c2 a1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp0 midp_b_c1c2 a2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_AOI211_4




.subckt SAEDRVT14_AOI21_1P5 vdd vss vbp vbn x a1 a2 b
xmn21 midn_b1_b21 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn11 x a1 midn_b1_b21 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x b vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp2 x b midp_a_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 midp_a_b1b2 a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp0 midp_a_b1b2 a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_AOI21_1P5




.subckt SAEDRVT14_AOI21_1 vdd vss vbp vbn x a1 a2 b
xmn2 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 x b midp_a_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b1b2 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_a_b1b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI21_1




.subckt SAEDRVT14_AOI21_2 vdd vss vbp vbn x a1 a2 b
xmn21 midn_b1_b21 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn11 x a1 midn_b1_b21 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x b vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp2 x b midp_a_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 midp_a_b1b2 a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp0 midp_a_b1b2 a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_AOI21_2




.subckt SAEDRVT14_AOI21_3 vdd vss vbp vbn x a1 a2 b
xmn2 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn0 x b vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmp2 x b midp_a_b1b2 vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 midp_a_b1b2 a1 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp0 midp_a_b1b2 a2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_AOI21_3




.subckt SAEDRVT14_AOI21_4 vdd vss vbp vbn x a1 a2 b
xmn2 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn0 x b vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmp2 x b midp_a_b1b2 vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 midp_a_b1b2 a1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp0 midp_a_b1b2 a2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_AOI21_4




.subckt SAEDRVT14_AOI21_6 vdd vss vbp vbn x a1 a2 b
xmn2 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn0 x b vss vbn n08_rev l=0.014u nf=6 m=1 nfin=2
xmp2 x b midp_a_b1b2 vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmp1 midp_a_b1b2 a1 vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmp0 midp_a_b1b2 a2 vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
.ends SAEDRVT14_AOI21_6




.subckt SAEDRVT14_AOI21_8 vdd vss vbp vbn x a1 a2 b
xmn2 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmn0 x b vss vbn n08_rev l=0.014u nf=8 m=1 nfin=2
xmp2 x b midp_a_b1b2 vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmp1 midp_a_b1b2 a1 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmp0 midp_a_b1b2 a2 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
.ends SAEDRVT14_AOI21_8




.subckt SAEDRVT14_AOI21_ECO_1 vdd vss vbp vbn x a1 a2 b
xmn2 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 x b midp_a_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b1b2 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_a_b1b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI21_ECO_1




.subckt SAEDRVT14_AOI21_V1_4 vdd vss vbp vbn x a1 a2 b
xmn2 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn0 x b vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmp2 midp_a_b1b2 b vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 x a1 midp_a_b1b2 vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp0 x a2 midp_a_b1b2 vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_AOI21_V1_4




.subckt SAEDRVT14_AOI21_V1_6 vdd vss vbp vbn x a1 a2 b
xmn2 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn0 x b vss vbn n08_rev l=0.014u nf=6 m=1 nfin=2
xmp2 midp_a_b1b2 b vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmp1 x a1 midp_a_b1b2 vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmp0 x a2 midp_a_b1b2 vbp p08_rev l=0.014u nf=6 m=1 nfin=4
.ends SAEDRVT14_AOI21_V1_6




.subckt SAEDRVT14_AOI21_V1_8 vdd vss vbp vbn x a1 a2 b
xmn2 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=8 m=1 nfin=3
xmn0 x b vss vbn n08_rev l=0.014u nf=8 m=1 nfin=2
xmp2 midp_a_b1b2 b vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmp1 x a1 midp_a_b1b2 vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmp0 x a2 midp_a_b1b2 vbp p08_rev l=0.014u nf=8 m=1 nfin=4
.ends SAEDRVT14_AOI21_V1_8




.subckt SAEDRVT14_AOI221_0P5 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 x1 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 x1 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 x1 a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_a1a2_b1b2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 midp_a1a2_b1b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOI221_0P5




.subckt SAEDRVT14_AOI22_0P75 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 x1 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn3 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x1 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x1 a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a1a2_b1b2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_a1a2_b1b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOI22_0P75




.subckt SAEDRVT14_AOI221_0P5 vdd vss vbp vbn x a1 a2 b1 b2 c
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 x1 a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x1 c vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 midn_c1_c2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 x1 b1 midn_c1_c2 vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 midp_a_b1b2 a1 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 midp_a_b1b2 a2 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 x1 c midp_a_b1b2 vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 midp_b1b2_c1c2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 midp_b1b2_c1c2 b2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_AOI221_0P5




.subckt SAEDRVT14_AOI221_1 vdd vss vbp vbn x a1 a2 b1 b2 c
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 x1 a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 x1 c vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 midn_c1_c2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 b1 midn_c1_c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 midp_a_b1b2 a1 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp4 midp_a_b1b2 a2 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 c midp_a_b1b2 vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 midp_b1b2_c1c2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_b1b2_c1c2 b2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_AOI221_1




.subckt SAEDRVT14_AOI221_2 vdd vss vbp vbn x a1 a2 b1 b2 c
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn51 x1 a1 midn_b1_b21 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn41 midn_b1_b21 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn21 midn_c1_c21 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn11 x1 b1 midn_c1_c21 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 x1 a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 x1 c vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 midn_c1_c2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 b1 midn_c1_c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 midp_a_b1b2 a1 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp4 midp_a_b1b2 a2 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp2 x1 c midp_a_b1b2 vbp p08_rev l=0.014u nf=5 m=1 nfin=4
xmp1 midp_b1b2_c1c2 b1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp0 midp_b1b2_c1c2 b2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_AOI221_2




.subckt SAEDRVT14_AOI221_4 vdd vss vbp vbn x a1 a2 b1 b2 c
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn53 x1 a1 midn_b1_b23 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn52 x1 a1 midn_b1_b22 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn51 x1 a1 midn_b1_b21 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn43 midn_b1_b23 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn42 midn_b1_b22 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn41 midn_b1_b21 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn23 midn_c1_c23 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn22 midn_c1_c22 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn21 midn_c1_c21 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn13 x1 b1 midn_c1_c23 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 x1 b1 midn_c1_c22 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn11 x1 b1 midn_c1_c21 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 x1 a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 midn_b1_b2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 x1 c vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 midn_c1_c2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 b1 midn_c1_c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 midp_a_b1b2 a1 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp4 midp_a_b1b2 a2 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=5 m=1 nfin=4
xmp2 x1 c midp_a_b1b2 vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 midp_b1b2_c1c2 b1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp0 midp_b1b2_c1c2 b2 vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=4
.ends SAEDRVT14_AOI221_4




.subckt SAEDRVT14_AOI22_1P5 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 x1 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn2 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp1 midp_a1a2_b1b2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_a1a2_b1b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI22_1P5




.subckt SAEDRVT14_AOI22_1 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 x1 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a1a2_b1b2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_a1a2_b1b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI22_1




.subckt SAEDRVT14_AOI222_0P5 vdd vss vbp vbn x a1 a2 b1 b2 c1 c2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn7 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn6 x1 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 x1 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 midn_c1_c2 c2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 x1 c1 midn_c1_c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp7 x1 a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp6 x1 a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 midp_a1a2_b1b2 b1 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 midp_a1a2_b1b2 b2 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_b1b2_c1c2 c1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 midp_b1b2_c1c2 c2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOI222_0P5




.subckt SAEDRVT14_AOI222_1 vdd vss vbp vbn x a1 a2 b1 b2 c1 c2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn7 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn6 x1 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn5 x1 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 midn_c1_c2 c2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 c1 midn_c1_c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp7 x1 a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp6 x1 a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp5 midp_a1a2_b1b2 b1 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 midp_a1a2_b1b2 b2 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_b1b2_c1c2 c1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_b1b2_c1c2 c2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI222_1




.subckt SAEDRVT14_AOI222_2 vdd vss vbp vbn x a1 a2 b1 b2 c1 c2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn7 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn6 x1 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn5 x1 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn2 midn_c1_c2 c2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 c1 midn_c1_c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp7 x1 a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp6 x1 a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp5 midp_a1a2_b1b2 b1 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 midp_a1a2_b1b2 b2 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp1 midp_b1b2_c1c2 c1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_b1b2_c1c2 c2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI222_2




.subckt SAEDRVT14_AOI222_4 vdd vss vbp vbn x a1 a2 b1 b2 c1 c2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn7 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn6 x1 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn5 x1 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn2 midn_c1_c2 c2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 c1 midn_c1_c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp7 x1 a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp6 x1 a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp5 midp_a1a2_b1b2 b1 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 midp_a1a2_b1b2 b2 midp_b1b2_c1c2 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp1 midp_b1b2_c1c2 c1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_b1b2_c1c2 c2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI222_4




.subckt SAEDRVT14_AOI222_2 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 x1 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn2 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp1 midp_a1a2_b1b2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_a1a2_b1b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI222_2




.subckt SAEDRVT14_AOI22_3 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 x1 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn2 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp1 midp_a1a2_b1b2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_a1a2_b1b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI22_3




.subckt SAEDRVT14_AOI22_4 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 x1 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn2 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp1 midp_a1a2_b1b2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_a1a2_b1b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI22_4




.subckt SAEDRVT14_AOI22_6 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 x1 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn2 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp1 midp_a1a2_b1b2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_a1a2_b1b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI22_6




.subckt SAEDRVT14_AOI22_ECO_1 vdd vss vbp vbn x a1 a2 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn4 x1 a1 midn_a1_a2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 midn_a1_a2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 midn_b1_b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x1 b1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 x1 a1 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 a2 midp_a1a2_b1b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a1a2_b1b2 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_a1a2_b1b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI22_ECO_1




.subckt SAEDRVT14_AOI31_0P5 vdd vss vbp vbn x a1 a2 a3 b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x1 a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x1 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_a_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 x1 b midp_a_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 midp_a_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOI31_0P5




.subckt SAEDRVT14_AOI31_0P75 vdd vss vbp vbn x a1 a2 a3 b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x1 a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 x1 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_a_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x1 b midp_a_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 midp_a_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOI31_0P75




.subckt SAEDRVT14_AOI311_0P5 vdd vss vbp vbn x a1 a2 a3 b1 b2
xn4 midn_c2_c3 a3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn3 x1 b1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 midn_c1_c2 a2 midn_c2_c3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn1 x1 a1 midn_c1_c2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn0 x1 b2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xp4 midp_b_c1c2c3 a3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 midp_a_b b2 midp_b_c1c2c3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x1 b1 midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 midp_b_c1c2c3 a1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 midp_b_c1c2c3 a2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOI311_0P5




.subckt SAEDRVT14_AOI311_0P75 vdd vss vbp vbn x a1 a2 a3 b1 b2
xn4 midn_c2_c3 a3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn3 x1 b1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 midn_c1_c2 a2 midn_c2_c3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn1 x1 a1 midn_c1_c2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn0 x1 b2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xp4 midp_b_c1c2c3 a3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 midp_a_b b2 midp_b_c1c2c3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x1 b1 midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 midp_b_c1c2c3 a1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 midp_b_c1c2c3 a2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOI311_0P75




.subckt SAEDRVT14_AOI311_1 vdd vss vbp vbn x a1 a2 a3 b1 b2
xn4 midn_c2_c3 a3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn3 x1 b1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 midn_c1_c2 a2 midn_c2_c3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn1 x1 a1 midn_c1_c2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn0 x1 b2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xp4 midp_b_c1c2c3 a3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 midp_a_b b2 midp_b_c1c2c3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x1 b1 midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 midp_b_c1c2c3 a1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 midp_b_c1c2c3 a2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOI311_1




.subckt SAEDRVT14_AOI311_2 vdd vss vbp vbn x a1 a2 a3 b1 b2
xn4 midn_c2_c3 a3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn3 x1 b1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 midn_c1_c2 a2 midn_c2_c3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn1 x1 a1 midn_c1_c2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn0 x1 b2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xp4 midp_b_c1c2c3 a3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 midp_a_b b2 midp_b_c1c2c3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x1 b1 midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 midp_b_c1c2c3 a1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 midp_b_c1c2c3 a2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOI311_2




.subckt SAEDRVT14_AOI311_4 vdd vss vbp vbn x a1 a2 a3 b1 b2
xn4 midn_c2_c3 a3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn3 x1 b1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 midn_c1_c2 a2 midn_c2_c3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn1 x1 a1 midn_c1_c2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn0 x1 b2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xp4 midp_b_c1c2c3 a3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 midp_a_b b2 midp_b_c1c2c3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x1 b1 midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 midp_b_c1c2c3 a1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 midp_b_c1c2c3 a2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOI311_4




.subckt SAEDRVT14_AOI31_1 vdd vss vbp vbn x a1 a2 a3 b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x1 a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 x1 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_a_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x1 b midp_a_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 midp_a_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOI31_1




.subckt SAEDRVT14_AOI31_2 vdd vss vbp vbn x a1 a2 a3 b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x1 a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 x1 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_a_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x1 b midp_a_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 midp_a_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOI31_2




.subckt SAEDRVT14_AOI31_4 vdd vss vbp vbn x a1 a2 a3 b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x1 a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 x1 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_a_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x1 b midp_a_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 midp_a_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOI31_4




.subckt SAEDRVT14_AOI31_ECO_1 vdd vss vbp vbn x a1 a2 a3 b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 a1 midn_b1_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x1 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_a_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 b midp_a_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_a_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOI31_ECO_1




.subckt SAEDRVT14_AOI32_0P5 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmn5 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=3
xmn4 x b1 midn_a1_a2 vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmn3 midn_a1_a2 b2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmn2 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=5 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=5 m=1 nfin=3
xmp4 midp_a1a2_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x b1 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp2 x b2 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp1 midp_a1a2_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 midp_a1a2_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOI32_0P5




.subckt SAEDRVT14_AOI32_0P75 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmn5 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn4 x b1 midn_a1_a2 vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmn3 midn_a1_a2 b2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmn2 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=7 m=1 nfin=3
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=7 m=1 nfin=3
xmp4 midp_a1a2_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 x b1 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x b2 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp1 midp_a1a2_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_a1a2_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOI32_0P75




.subckt SAEDRVT14_AOI32_1 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmn5 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn4 x b1 midn_a1_a2 vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn3 midn_a1_a2 b2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn2 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=7 m=1 nfin=4
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=7 m=1 nfin=4
xmp4 midp_a1a2_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 x b1 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x b2 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 midp_a1a2_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_a1a2_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI32_1




.subckt SAEDRVT14_AOI32_2 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmn2_2 midn_b1_b2_2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1_2 x a1 midn_b1_b2_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmn4 x b1 midn_a1_a2 vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn3 midn_a1_a2 b2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn2 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmp4 midp_a1a2_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 x b1 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x b2 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a1a2_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_a1a2_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI32_2




.subckt SAEDRVT14_AOI32_4 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmn2_4 midn_b1_b2_4 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2_3 midn_b1_b2_3 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2_2 midn_b1_b2_2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1_4 x a1 midn_b1_b2_4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1_3 x a1 midn_b1_b2_3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1_2 x a1 midn_b1_b2_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 midn_b2_b3 a3 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmn4 x b1 midn_a1_a2 vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn3 midn_a1_a2 b2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn2 midn_b1_b2 a2 midn_b2_b3 vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmn1 x a1 midn_b1_b2 vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmp4 midp_a1a2_b1b2b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 x b1 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp2 x b2 midp_a1a2_b1b2b3 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 midp_a1a2_b1b2b3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_a1a2_b1b2b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI32_4




.subckt SAEDRVT14_AOI33_0P5 vdd vss vbp vbn x a1 a2 a3 b1 b2 b3
xmn6 midn_a2_a3 a3 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn5 midn_b2_b3 b3 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=3
xmn4 x a1 midn_a1_a2 vbn n08_rev l=0.014u nf=5 m=1 nfin=3
xmn3 midn_a1_a2 a2 midn_a2_a3 vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn2 midn_b1_b2 b2 midn_b2_b3 vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn1 x b1 midn_b1_b2 vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmp5 x a3 midp_a1a2a3_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp4 midp_a1a2a3_b1b2b3 b3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x a1 midp_a1a2a3_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x a2 midp_a1a2a3_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_a1a2a3_b1b2b3 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 midp_a1a2a3_b1b2b3 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOI33_0P5




.subckt SAEDRVT14_AOI33_0P75 vdd vss vbp vbn x a1 a2 a3 b1 b2 b3
xmn6 midn_a2_a3 a3 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn5 midn_b2_b3 b3 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn4 x a1 midn_a1_a2 vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn3 midn_a1_a2 a2 midn_a2_a3 vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn2 midn_b1_b2 b2 midn_b2_b3 vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn1 x b1 midn_b1_b2 vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmp5 x a3 midp_a1a2a3_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp4 midp_a1a2a3_b1b2b3 b3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 x a1 midp_a1a2a3_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x a2 midp_a1a2a3_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_a1a2a3_b1b2b3 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_a1a2a3_b1b2b3 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOI33_0P75




.subckt SAEDRVT14_AOI33_1 vdd vss vbp vbn x a1 a2 a3 b1 b2 b3
xmn6 midn_a2_a3 a3 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn5 midn_b2_b3 b3 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn4 x a1 midn_a1_a2 vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn3 midn_a1_a2 a2 midn_a2_a3 vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn2 midn_b1_b2 b2 midn_b2_b3 vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn1 x b1 midn_b1_b2 vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmp5 x a3 midp_a1a2a3_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 midp_a1a2a3_b1b2b3 b3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 x a1 midp_a1a2a3_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x a2 midp_a1a2a3_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a1a2a3_b1b2b3 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_a1a2a3_b1b2b3 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI33_1




.subckt SAEDRVT14_AOI33_2 vdd vss vbp vbn x a1 a2 a3 b1 b2 b3
xmn41 x a1 midn_a1_a21 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn31 midn_a1_a21 a2 midn_a2_a3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn21 midn_b1_b21 b2 midn_b2_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn11 x b1 midn_b1_b21 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn6 midn_a2_a3 a3 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmn5 midn_b2_b3 b3 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmn4 x a1 midn_a1_a2 vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmn3 midn_a1_a2 a2 midn_a2_a3 vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmn2 midn_b1_b2 b2 midn_b2_b3 vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmn1 x b1 midn_b1_b2 vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmp5 x a3 midp_a1a2a3_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 midp_a1a2a3_b1b2b3 b3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 x a1 midp_a1a2a3_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x a2 midp_a1a2a3_b1b2b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a1a2a3_b1b2b3 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_a1a2a3_b1b2b3 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOI33_2




.subckt SAEDRVT14_AOLVLUBUFE0_IY2V1_8 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE0_IY2V1_8




.subckt SAEDRVT14_AOINV_IW_0P5 vdd vss x a vddr
xmmn0 x a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xmmp0 x a vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOINV_IW_0P5




.subckt SAEDRVT14_AOINV_IW_1 vdd vss x a vddr
xmmn0 x a vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xmmp0 x a vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOINV_IW_1




.subckt SAEDRVT14_AOINV_IW_2 vdd vss x a vddr
xmmn0 x a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmmp0 x a vddr vdd p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_AOINV_IW_2




.subckt SAEDRVT14_AOINV_IW_4 vdd vss x a vddr
xmmn0 x a vss vss n08_rev l=0.014u nf=4 m=1 nfin=3
xmmp0 x a vddr vdd p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_AOINV_IW_4




.subckt SAEDRVT14_AOINV_IW_6 vdd vss x a vddr
xmmn0 x a vss vss n08_rev l=0.014u nf=6 m=1 nfin=3
xmmp0 x a vddr vdd p08_rev l=0.014u nf=6 m=1 nfin=4
.ends SAEDRVT14_AOINV_IW_6




.subckt SAEDRVT14_AOLVLUBUFE0_IY2_10 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE0_IY2_10




.subckt SAEDRVT14_AOLVLUBUFE0_IY2_12 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE0_IY2_12




.subckt SAEDRVT14_AOLVLUBUFE0_IY2_1 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUFE0_IY2_1




.subckt SAEDRVT14_AOLVLUBUFE0_IY2_2 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUFE0_IY2_2




.subckt SAEDRVT14_AOLVLUBUFE0_IY2_3 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUFE0_IY2_3




.subckt SAEDRVT14_AOLVLUBUFE0_IY2_4 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE0_IY2_4




.subckt SAEDRVT14_AOLVLUBUFE0_IY2_6 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE0_IY2_6




.subckt SAEDRVT14_AOLVLUBUFE0_IY2_8 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE0_IY2_8




.subckt SAEDRVT14_AOLVLUBUFE0_IY2V1_10 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE0_IY2V1_10




.subckt SAEDRVT14_AOLVLUBUFE0_IY2V1_12 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE0_IY2V1_12




.subckt SAEDRVT14_AOLVLUBUFE0_IY2V1_1 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUFE0_IY2V1_1




.subckt SAEDRVT14_AOLVLUBUFE0_IY2V1_2 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=2 m=2 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE0_IY2V1_2




.subckt SAEDRVT14_AOLVLUBUFE0_IY2V1_3 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE0_IY2V1_3




.subckt SAEDRVT14_AOLVLUBUFE0_IY2V1_4 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE0_IY2V1_4




.subckt SAEDRVT14_AOLVLUBUFE0_IY2V1_6 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE0_IY2V1_6




.subckt SAEDRVT14_AOLVLUBUFE0_IY2V1_8 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE0_IY2V1_8


SAEDRVT14_AOLVLUBUF_E1_IY2_10

.subckt SAEDRVT14_AOLVLUBUF_E1_IY2_10 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUF_E1_IY2_10




.subckt SAEDRVT14_AOLVLUBUFE1_IY2_10 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE1_IY2_10




.subckt SAEDRVT14_AOLVLUBUF_E1_IY2_12 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUF_E1_IY2_12




.subckt SAEDRVT14_AOLVLUBUFE1_IY2_12 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE1_IY2_12




.subckt SAEDRVT14_AOLVLUBUF_E1_IY2_1 vss vddi x a en vddr
xn5 x net16 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_E1_IY2_1




.subckt SAEDRVT14_AOLVLUBUFE1_IY2_1 vss x a en vddl vddr
xn5 x net16 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUFE1_IY2_1




.subckt SAEDRVT14_AOLVLUBUF_E1_IY2_2 vss vddi x a en vddr
xn5 x net16 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_E1_IY2_2




.subckt SAEDRVT14_AOLVLUBUFE1_IY2_2 vss x a en vddl vddr
xn5 x net16 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUFE1_IY2_2




.subckt SAEDRVT14_AOLVLUBUF_E1_IY2_3 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_E1_IY2_3




.subckt SAEDRVT14_AOLVLUBUFE1_IY2_3 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUFE1_IY2_3




.subckt SAEDRVT14_AOLVLUBUF_E1_IY2_4 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_E1_IY2_4




.subckt SAEDRVT14_AOLVLUBUFE1_IY2_4 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUFE1_IY2_4




.subckt SAEDRVT14_AOLVLUBUF_E1_IY2_6 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_E1_IY2_6




.subckt SAEDRVT14_AOLVLUBUFE1_IY2_6 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUFE1_IY2_6




.subckt SAEDRVT14_AOLVLUBUF_E1_IY2_8 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOLVLUBUF_E1_IY2_8




.subckt SAEDRVT14_AOLVLUBUFE1_IY2_8 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOLVLUBUFE1_IY2_8




.subckt SAEDRVT14_AOLVLUBUF_E1_IY2V1_10 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUF_E1_IY2V1_10




.subckt SAEDRVT14_AOLVLUBUFE1_IY2V1_10 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE1_IY2V1_10




.subckt SAEDRVT14_AOLVLUBUF_E1_IY2V1_12 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUF_E1_IY2V1_12




.subckt SAEDRVT14_AOLVLUBUFE1_IY2V1_12 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_AOLVLUBUFE1_IY2V1_12




.subckt SAEDRVT14_AOLVLUBUF_E1_IY2V1_1 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_E1_IY2V1_1




.subckt SAEDRVT14_AOLVLUBUFE1_IY2V1_1 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUFE1_IY2V1_1




.subckt SAEDRVT14_BUF_PECO_4 a vbn vbp vddr vss x
xn1 x int_zn vss vbn n08_rev2 l=0.014u nf=4 m=1 nfin=3
xn0 int_zn a vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=3
xp1 x int_zn vddr vbp p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp0 int_zn a vddr vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_BUF_PECO_4




.subckt SAEDRVT14_AOLVLUBUFE1_IY2V1_2 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUFE1_IY2V1_2




.subckt SAEDRVT14_AOLVLUBUF_E1_IY2V1_3 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_E1_IY2V1_3




.subckt SAEDRVT14_AOLVLUBUFE1_IY2V1_3 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUFE1_IY2V1_3




.subckt SAEDRVT14_AOLVLUBUF_E1_IY2V1_4 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_E1_IY2V1_4




.subckt SAEDRVT14_AOLVLUBUFE1_IY2V1_4 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUFE1_IY2V1_4




.subckt SAEDRVT14_AOLVLUBUF_E1_IY2V1_6 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_E1_IY2V1_4




.subckt SAEDRVT14_AOLVLUBUFE1_IY2V1_6 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUFE1_IY2V1_6




.subckt SAEDRVT14_AOLVLUBUF_E1_IY2V1_8 vddr vss vddi x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOLVLUBUF_E1_IY2V1_8




.subckt SAEDRVT14_AOLVLUBUFE1_IY2V1_8 vddr vss x a en vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddr vddr p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 net_025 vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_AOLVLUBUFE1_IY2V1_8




.subckt SAEDRVT14_AOLVLUBUF_IY2V1_10 vddr vss x a vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=9 m=1 nfin=4
xp4 x net14 vddr vddr p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp3 net14 net1 vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_IY2V1_10




.subckt SAEDRVT14_AOLVLUBUF_IY2V1_12 vddr vss x a vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=9 m=1 nfin=4
xp4 x net14 vddr vddr p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp3 net14 net1 vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_IY2V1_12




.subckt SAEDRVT14_AOLVLUBUF_IY2V1_1 vddr vss x a vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=7 m=1 nfin=4
xp4 x net14 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net14 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net1 net2 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_IY2V1_1




.subckt SAEDRVT14_AOLVLUBUF_IY2V1_2 vddr vss x a vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=7 m=1 nfin=4
xp4 x net14 vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net14 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net1 net2 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_IY2V1_2




.subckt SAEDRVT14_AOLVLUBUF_IY2V1_3 vddr vss x a vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=7 m=1 nfin=4
xp4 x net14 vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net14 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net1 net2 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_IY2V1_3




.subckt SAEDRVT14_AOLVLUBUF_IY2V1_4 vddr vss x a vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=7 m=1 nfin=4
xp4 x net14 vddr vddr p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp3 net14 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net1 net2 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_IY2V1_4




.subckt SAEDRVT14_AOLVLUBUF_IY2V1_6 vddr vss x a vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=9 m=1 nfin=4
xp4 x net14 vddr vddr p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp3 net14 net1 vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp2 net1 net2 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_IY2V1_6




.subckt SAEDRVT14_AOLVLUBUF_IY2V1_8 vddr vss x a vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=9 m=1 nfin=4
xp4 x net14 vddr vddr p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp3 net14 net1 vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp2 net1 net2 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOLVLUBUF_IY2V1_8




.subckt SAEDRVT14_AOTIE0_IW vdd vddr vss x
xmn0 x net16 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 net16 net16 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOTIE0_IW




.subckt SAEDRVT14_AOTIE1_IW vdd vddr vss x
xmn0 net19 net19 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 x net19 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_AOTIE1_IW




.subckt SAEDRVT14_BUF_10 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=10 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=10 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_BUF_10



.subckt SAEDRVT14_BUF_12 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=12 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=12 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_BUF_12




.subckt SAEDRVT14_BUF_16 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=16 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=16 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=4
.ends SAEDRVT14_BUF_16




.subckt SAEDRVT14_BUF_1P5 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_BUF_1P5




.subckt SAEDRVT14_BUF_1 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_BUF_1




.subckt SAEDRVT14_BUF_20 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=20 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=20 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
.ends SAEDRVT14_BUF_20




.subckt SAEDRVT14_BUF_2 vdd vss vbp vbn x a
xmmn2 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn1 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmp2 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp1 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_BUF_2




.subckt SAEDRVT14_BUF_3 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_BUF_3




.subckt SAEDRVT14_BUF_4 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_BUF_4




.subckt SAEDRVT14_BUF_6 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_BUF_6




.subckt SAEDRVT14_BUF_8 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_BUF_8




.subckt SAEDRVT14_BUF_CDC_2 vdd vss vbp vbn x a
xmmn2 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn1 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmp2 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp1 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_BUF_CDC_2




.subckt SAEDRVT14_BUF_CDC_4 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_BUF_CDC_4




.subckt SAEDRVT14_BUF_ECO_1 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_BUF_ECO_1




.subckt SAEDRVT14_BUF_ECO_2 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_BUF_ECO_2




.subckt SAEDRVT14_BUF_ECO_3 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_BUF_ECO_3




.subckt SAEDRVT14_BUF_ECO_4 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_BUF_ECO_4




.subckt SAEDRVT14_BUF_ECO_6 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_BUF_ECO_6




.subckt SAEDRVT14_BUF_ECO_7 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=7 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=7 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_BUF_ECO_7




.subckt SAEDRVT14_BUF_ECO_8 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_BUF_ECO_8




.subckt SAEDRVT14_BUF_PECO_12 A VBN VBP VDDR VSS X
Mxn1 X int_zn VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxn0 int_zn A VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxp1 X int_zn VDDR VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxp0 int_zn A VDDR VBP p08 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_BUF_PECO_12




.subckt SAEDRVT14_BUF_PECO_1 a vbn vbp vdd vddr vss x
xp1 x int_zn vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp0 int_zn a vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp1 net14 net14 net14 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xn1 x int_zn vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn0 int_zn a vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xmn1 net14 net14 net14 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_BUF_PECO_1




.subckt SAEDRVT14_BUF_PECO_2 a vbn vbp vddr vss x
xn1 x int_zn vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=3
xn0 int_zn a vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp1 x int_zn vddr vbp p08_rev2 l=0.014u nf=2 m=2 nfin=4
xp0 int_zn a vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_BUF_PECO_2




.subckt SAEDRVT14_BUF_PECO_4 A VBN VBP VDDR VSS X
Mxn1 X int_zn VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxn0 int_zn A VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxp1 X int_zn VDDR VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxp0 int_zn A VDDR VBP p08 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_BUF_PECO_4




.subckt SAEDRVT14_BUF_PECO_8 a vbn vbp vddr vss x
xn1 x int_zn vss vbn n08_rev2 l=0.014u nf=4 m=1 nfin=3
xn0 int_zn a vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=3
xp1 x int_zn vddr vbp p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp0 int_zn a vddr vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_BUF_PECO_8




.subckt SAEDRVT14_BUF_PS_0P75 a vbn vbp vddr vss x
xn1 x int_zn vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn0 int_zn a vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp1 x int_zn vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp0 int_zn a vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_BUF_PS_0P75




.subckt SAEDRVT14_BUF_PS_1P5 vdd vss vddr x a
xn1 x int_zn vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=3
xn0 int_zn a vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp1 x int_zn vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=3
xp0 int_zn a vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_BUF_PS_1P5




.subckt SAEDRVT14_BUF_PS_3 vdd vss vddr x a
xn1 x int_zn vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=3
xn0 int_zn a vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=3
xp1 x int_zn vddr vddr p08_rev2 l=0.014u nf=4 m=1 nfin=3
xp0 int_zn a vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_BUF_PS_3




.subckt SAEDRVT14_BUF_PS_6 vdd vss vddr x a
xn1 x int_zn vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=3
xn0 int_zn a vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=3
xp1 x int_zn vddr vddr p08_rev2 l=0.014u nf=8 m=1 nfin=3
xp0 int_zn a vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=3
.ends SAEDRVT14_BUF_PS_6




.subckt SAEDRVT14_BUF_S_0P5 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_BUF_S_0P5




.subckt SAEDRVT14_BUF_S_0P75 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_BUF_S_0P75




.subckt SAEDRVT14_BUF_S_10 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=10 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=10 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_BUF_S_10




.subckt SAEDRVT14_BUF_UCDC_0P5 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_BUF_UCDC_0P5




.subckt SAEDRVT14_BUF_S_16 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=16 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=16 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=4
.ends SAEDRVT14_BUF_S_16




.subckt SAEDRVT14_BUF_S_1P5 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=1 m=2 nfin=3
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=2 nfin=3
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_BUF_S_1P5




.subckt SAEDRVT14_BUF_S_1 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_BUF_S_1




.subckt SAEDRVT14_BUF_S_20 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=20 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=20 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
.ends SAEDRVT14_BUF_S_20




.subckt SAEDRVT14_BUF_S_2 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_BUF_S_2




.subckt SAEDRVT14_BUF_S_3 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_BUF_S_3




.subckt SAEDRVT14_BUF_S_4 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_BUF_S_4




.subckt SAEDRVT14_BUF_S_6 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_BUF_S_6




.subckt SAEDRVT14_BUF_S_8 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_BUF_S_8




.subckt SAEDRVT14_BUF_U_0P5 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_BUF_U_0P5




.subckt SAEDRVT14_BUF_U_0P75 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_BUF_U_0P75




.subckt SAEDRVT14_BUF_UCDC_0P5 VDD VSS VBP VBN X A
Mxmn1 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn0 int_zn A VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp1 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 int_zn A VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_BUF_UCDC_0P5




.subckt SAEDRVT14_BUF_UCDC_1 vdd vss vbp vbn x a
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 int_zn a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 int_zn a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_BUF_UCDC_1




.subckt SAEDRVT14_CAPB2 vdd vss
.ends SAEDRVT14_CAPB2




.subckt SAEDRVT14_CAPB3 vdd vss
.ends SAEDRVT14_CAPB3



.subckt SAEDRVT14_CAPBC8 vdd vss
.ends SAEDRVT14_CAPBC8




.subckt SAEDRVT14_CAPBIN13 vdd vss
.ends SAEDRVT14_CAPBIN13




.subckt SAEDRVT14_CAPBTAP6 vdd vss
.ends SAEDRVT14_CAPBTAP6




.subckt SAEDRVT14_CAPLR8 vdd vss vbp vbn
.ends SAEDRVT14_CAPLR8




.subckt SAEDRVT14_CAPSPACER1 VDD VSS VBP VBN
.ends SAEDRVT14_CAPSPACER1




.subckt SAEDRVT14_CAPT2 vdd vss
.ends SAEDRVT14_CAPT2




.subckt SAEDRVT14_CAPT3 vdd vss
.ends SAEDRVT14_CAPT3




.subckt SAEDRVT14_CAPTC8 vdd vss
.ends SAEDRVT14_CAPTC8




.subckt SAEDRVT14_CAPTIN13 vdd vss
.ends SAEDRVT14_CAPTIN13




.subckt SAEDRVT14_CAPTTAP6 vdd vss
.ends SAEDRVT14_CAPTTAP6




.subckt SAEDRVT14_CAPTTAPP6 vdd vss vddr
.ends SAEDRVT14_CAPTTAPP6




.subckt SAEDRVT14_CKGTNLT_V5_12 vdd vss vbp vbn q ck en se
xmn24 nmose_nr_te se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 zn net013 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn16 zn ck vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn14 q zn vss vbn n08_rev l=0.014u nf=12 m=1 nfin=4
xmn10 nmose_nr_te en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn10 net013 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmose_nr_te ckbb i1 vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn12 i1 ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp23 pmose_nr_te se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 net021 net013 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp19 zn ck net021 vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp11 q zn vdd vbp p08_rev l=0.014u nf=12 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp10 net013 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp21 i1 ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckb pmose_nr_te vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_CKGTNLT_V5_12




.subckt SAEDRVT14_CKGTNLT_V5_1 vdd vss vbp vbn q ck en se
xmn24 nmose_nr_te se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 zn net013 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn16 zn ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn14 q zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn10 nmose_nr_te en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn10 net013 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmose_nr_te ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 pmose_nr_te se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 net018 net013 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp19 zn ck net018 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp11 q zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp10 net013 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp21 i1 ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckb pmose_nr_te vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKGTNLT_V5_1




.subckt SAEDRVT14_CKGTNLT_V5_2 vdd vss vbp vbn q ck en se
xmn24 nmose_nr_te se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 zn net013 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn16 zn ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn14 q zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn10 nmose_nr_te en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn10 net013 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmose_nr_te ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 pmose_nr_te se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 net019 net013 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp19 zn ck net019 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp11 q zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp10 net013 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp21 i1 ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckb pmose_nr_te vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKGTNLT_V5_2




.subckt SAEDRVT14_CKGTNLT_V5_3 vdd vss vbp vbn q ck en se
xmn24 nmose_nr_te se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 zn net013 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn16 zn ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn14 q zn vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn10 nmose_nr_te en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn10 net013 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmose_nr_te ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 pmose_nr_te se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 net019 net013 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp19 zn ck net019 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp11 q zn vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp10 net013 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp21 i1 ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckb pmose_nr_te vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKGTNLT_V5_3




.subckt SAEDRVT14_CKGTNLT_V5_4 vdd vss vbp vbn q ck en se
xmn24 nmose_nr_te se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 zn net013 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn16 zn ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn14 q zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn10 nmose_nr_te en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn10 net013 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmose_nr_te ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 pmose_nr_te se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 net019 net013 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp19 zn ck net019 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp11 q zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp10 net013 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp21 i1 ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckb pmose_nr_te vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKGTNLT_V5_4




.subckt SAEDRVT14_CKGTNLT_V5_5 vdd vss vbp vbn q ck en se
xmn24 nmose_nr_te se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 zn net013 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn16 zn ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn14 q zn vss vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmn10 nmose_nr_te en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn10 net013 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmose_nr_te ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 i1 ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp23 pmose_nr_te se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 net019 net013 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp19 zn ck net019 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp11 q zn vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp10 net013 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp21 i1 ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckb pmose_nr_te vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_CKGTNLT_V5_5




.subckt SAEDRVT14_CKGTNLT_V5_6 vdd vss vbp vbn q ck se e
xmn24 nmose_nr_te se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 zn net013 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn16 zn ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn14 q zn vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn10 nmose_nr_te e vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn10 net013 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmose_nr_te ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 i1 ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp23 pmose_nr_te se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 e vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 net019 net013 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp19 zn ck net019 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp11 q zn vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp10 net013 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp21 i1 ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckb pmose_nr_te vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_CKGTNLT_V5_6




.subckt SAEDRVT14_CKGTNLT_V5_8 vdd vss vbp vbn q ck en se
xmn24 nmose_nr_te se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 zn net013 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmn16 zn ck vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmn14 q zn vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmn10 nmose_nr_te en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn10 net013 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmose_nr_te ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 i1 ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp23 pmose_nr_te se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 net018 net013 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp19 zn ck net018 vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp11 q zn vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp10 net013 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp21 i1 ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckb pmose_nr_te vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_CKGTNLT_V5_8




.subckt SAEDRVT14_CKGTPLT_V5_12 vdd vss vbp vbn q ck en se
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fn13 i31#2fmidn_en_ck3 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn12 i31#2fmidn_en_ck2 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn11 i31#2fmidn_en_ck1 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn03 zn ck i31#2fmidn_en_ck3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn02 zn ck i31#2fmidn_en_ck2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn01 zn ck i31#2fmidn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn2 q zn vss vbn n08_rev l=0.014u nf=12 m=1 nfin=4
xmi31#2fn1 i31#2fmidn_en_ck i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn0 zn ck i31#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp23 net014 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fp2 q zn vdd vbp p08_rev l=0.014u nf=12 m=1 nfin=4
xmi31#2fp1 zn ck vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmi31#2fp0 zn i2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net014 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_CKGTPLT_V5_12




.subckt SAEDRVT14_CKGTPLT_V5_16 vdd vss vbp vbn q ck en se
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fn13 i31#2fmidn_en_ck3 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn12 i31#2fmidn_en_ck2 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn11 i31#2fmidn_en_ck1 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn03 zn ck i31#2fmidn_en_ck3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn02 zn ck i31#2fmidn_en_ck2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn01 zn ck i31#2fmidn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn2 q zn vss vbn n08_rev l=0.014u nf=16 m=1 nfin=4
xmi31#2fn1 i31#2fmidn_en_ck i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn0 zn ck i31#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp23 net014 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fp2 q zn vdd vbp p08_rev l=0.014u nf=16 m=1 nfin=4
xmi31#2fp1 zn ck vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmi31#2fp0 zn i2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net014 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_CKGTPLT_V5_16




.subckt SAEDRVT14_CKGTPLT_V5_1 vdd vss vbp vbn q ck en se
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fn2 q zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn1 i31#2fmidn_en_ck i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fn0 zn ck i31#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 net014 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fp2 q zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fp1 zn ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fp0 zn i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net014 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKGTPLT_V5_1




.subckt SAEDRVT14_CKGTPLT_V5_20 vdd vss vbp vbn q ck en se
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fn14 i31#2fmidn_en_ck4 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn13 i31#2fmidn_en_ck3 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn12 i31#2fmidn_en_ck2 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn11 i31#2fmidn_en_ck1 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn04 zn ck i31#2fmidn_en_ck4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn03 zn ck i31#2fmidn_en_ck3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn02 zn ck i31#2fmidn_en_ck2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn01 zn ck i31#2fmidn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn2 q zn vss vbn n08_rev l=0.014u nf=20 m=1 nfin=4
xmi31#2fn1 i31#2fmidn_en_ck i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn0 zn ck i31#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp23 net014 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fp2 q zn vdd vbp p08_rev l=0.014u nf=20 m=1 nfin=4
xmi31#2fp1 zn ck vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=3
xmi31#2fp0 zn i2 vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=3
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net014 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_CKGTPLT_V5_20




.subckt SAEDRVT14_CKGTPLT_V5_24 vdd vss vbp vbn q ck en se
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fn15 i31#2fmidn_en_ck5 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn14 i31#2fmidn_en_ck4 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn13 i31#2fmidn_en_ck3 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn12 i31#2fmidn_en_ck2 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn11 i31#2fmidn_en_ck1 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn05 zn ck i31#2fmidn_en_ck5 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn04 zn ck i31#2fmidn_en_ck4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn03 zn ck i31#2fmidn_en_ck3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn02 zn ck i31#2fmidn_en_ck2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn01 zn ck i31#2fmidn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn2 q zn vss vbn n08_rev l=0.014u nf=24 m=1 nfin=4
xmi31#2fn1 i31#2fmidn_en_ck i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn0 zn ck i31#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp23 net014 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fp2 q zn vdd vbp p08_rev l=0.014u nf=24 m=1 nfin=4
xmi31#2fp1 zn ck vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=3
xmi31#2fp0 zn i2 vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=3
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net014 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_CKGTPLT_V5_24




.subckt SAEDRVT14_CKGTPLT_V5_2 vdd vss vbp vbn q ck en se
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fn2 q zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi31#2fn1 i31#2fmidn_en_ck i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fn0 zn ck i31#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 net014 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fp2 q zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi31#2fp1 zn ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fp0 zn i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net014 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKGTPLT_V5_2




.subckt SAEDRVT14_CKGTPLT_V5_3 vdd vss vbp vbn q ck en se
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fn2 q zn vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmi31#2fn1 i31#2fmidn_en_ck i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn0 zn ck i31#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 net014 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fp2 q zn vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmi31#2fp1 zn ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fp0 zn i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net014 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKGTPLT_V5_3




.subckt SAEDRVT14_CKGTPLT_V5_4 vdd vss vbp vbn q ck en se
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fn11 i31#2fmidn_en_ck1 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fn01 zn ck i31#2fmidn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fn2 q zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi31#2fn1 i31#2fmidn_en_ck i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fn0 zn ck i31#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 net014 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi31#2fp2 q zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi31#2fp1 zn ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi31#2fp0 zn i2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net014 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKGTPLT_V5_4




.subckt SAEDRVT14_CKGTPLT_V5_5 vdd vss vbp vbn q ck en se
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fn11 i31#2fmidn_en_ck1 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fn01 zn ck i31#2fmidn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fn2 q zn vss vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmi31#2fn1 i31#2fmidn_en_ck i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fn0 zn ck i31#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp23 net014 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fp2 q zn vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=4
xmi31#2fp1 zn ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi31#2fp0 zn i2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net014 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_CKGTPLT_V5_5




.subckt SAEDRVT14_CKGTPLT_V5_6 vdd vss vbp vbn q ck en se
xmn24 nmose_nr_te se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 zn net013 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn16 zn ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn14 q zn vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn10 nmose_nr_te en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn10 net013 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmose_nr_te ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 i1 ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp23 pmose_nr_te se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 net019 net013 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp19 zn ck net019 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp11 q zn vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp10 net013 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp21 i1 ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckb pmose_nr_te vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_CKGTPLT_V5_6




.subckt SAEDRVT14_CKGTPLT_V5_8 vdd vss vbp vbn q ck en se
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fn12 i31#2fmidn_en_ck2 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn11 i31#2fmidn_en_ck1 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn02 zn ck i31#2fmidn_en_ck2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn01 zn ck i31#2fmidn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn2 q zn vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmi31#2fn1 i31#2fmidn_en_ck i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi31#2fn0 zn ck i31#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp23 net014 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi31#2fp2 q zn vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmi31#2fp1 zn ck vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmi31#2fp0 zn i2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net014 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_CKGTPLT_V5_8




.subckt SAEDRVT14_CKGTPL_V5_0P5 vdd vss vbp vbn q ck en
xmi1#2fn2 q int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn1 i1#2fmidn_en_ck net9 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn0 int_zn ck i1#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn24 i0#2fnet12 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 i0#2fckbb i0#2fckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi2#2fn0 net9 i0#2fi1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fn23 i0#2fi1#2fnet61 i0#2fi2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fn20 i0#2fnet12 i0#2fckb i0#2fi1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fn12 i0#2fi1 i0#2fckbb i0#2fi1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fn10 i0#2fi2 i0#2fi1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp2 q int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp1 int_zn ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 int_zn net9 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp23 i0#2fnet13 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 i0#2fckbb i0#2fckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi2#2fp1 net9 i0#2fi1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fp21 i0#2fi1 i0#2fckb i0#2fi1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fp18 i0#2fi1 i0#2fckbb i0#2fnet13 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fp9 i0#2fi1#2fnet98 i0#2fi2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fp8 i0#2fi2 i0#2fi1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKGTPL_V5_0P5




.subckt SAEDRVT14_CKGTPL_V5_1 vdd vss vbp vbn q ck en
xmi1#2fn2 q int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 i1#2fmidn_en_ck net9 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 int_zn ck i1#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn24 i0#2fnet12 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn1 i0#2fckbb i0#2fckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi2#2fn0 net9 i0#2fi1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi1#2fn23 i0#2fi1#2fnet61 i0#2fi2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fn20 i0#2fnet12 i0#2fckb i0#2fi1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fn12 i0#2fi1 i0#2fckbb i0#2fi1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fn10 i0#2fi2 i0#2fi1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp2 q int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 int_zn ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 int_zn net9 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp23 i0#2fnet13 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp1 i0#2fckbb i0#2fckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi2#2fp1 net9 i0#2fi1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi1#2fp21 i0#2fi1 i0#2fckb i0#2fi1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fp18 i0#2fi1 i0#2fckbb i0#2fnet13 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fp9 i0#2fi1#2fnet98 i0#2fi2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fp8 i0#2fi2 i0#2fi1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKGTPL_V5_1




.subckt SAEDRVT14_CKGTPL_V5_2 vdd vss vbp vbn q ck en
xmi1#2fn2 q int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 i1#2fmidn_en_ck net9 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 int_zn ck i1#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn24 i0#2fnet12 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn1 i0#2fckbb i0#2fckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi2#2fn0 net9 i0#2fi1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi1#2fn23 i0#2fi1#2fnet61 i0#2fi2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fn20 i0#2fnet12 i0#2fckb i0#2fi1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fn12 i0#2fi1 i0#2fckbb i0#2fi1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fn10 i0#2fi2 i0#2fi1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp2 q int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 int_zn ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 int_zn net9 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp23 i0#2fnet13 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp1 i0#2fckbb i0#2fckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi2#2fp1 net9 i0#2fi1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi1#2fp21 i0#2fi1 i0#2fckb i0#2fi1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fp18 i0#2fi1 i0#2fckbb i0#2fnet13 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fp9 i0#2fi1#2fnet98 i0#2fi2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fp8 i0#2fi2 i0#2fi1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKGTPL_V5_2




.subckt SAEDRVT14_CKGTPL_V5_4 vdd vss vbp vbn q ck en
xmi1#2fn2 q int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 i1#2fmidn_en_ck net9 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 int_zn ck i1#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn24 i0#2fnet12 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn1 i0#2fckbb i0#2fckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi2#2fn0 net9 i0#2fi1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi1#2fn23 i0#2fi1#2fnet61 i0#2fi2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fn20 i0#2fnet12 i0#2fckb i0#2fi1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fn12 i0#2fi1 i0#2fckbb i0#2fi1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fn10 i0#2fi2 i0#2fi1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp2 q int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 int_zn ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 int_zn net9 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp23 i0#2fnet13 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp1 i0#2fckbb i0#2fckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi2#2fp1 net9 i0#2fi1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi1#2fp21 i0#2fi1 i0#2fckb i0#2fi1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fp18 i0#2fi1 i0#2fckbb i0#2fnet13 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fp9 i0#2fi1#2fnet98 i0#2fi2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi1#2fp8 i0#2fi2 i0#2fi1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKGTPL_V5_4




.subckt SAEDRVT14_CKINVGTPLT_V7_1 vdd vss vbp vbn qb ck en se
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 net43 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn16 qb ck net43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 net016 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 qb i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp19 qb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net016 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKINVGTPLT_V7_1




.subckt SAEDRVT14_CKINVGTPLT_V7_2 vdd vss vbp vbn qb ck en se
xmn171 net431 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn161 qb ck net431 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 net43 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn16 qb ck net43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 net016 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 qb i2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp19 qb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net016 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKINVGTPLT_V7_2




.subckt SAEDRVT14_CKINVGTPLT_V7_3 vdd vss vbp vbn qb ck en se
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 net43 i2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmn16 qb ck net43 vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 net016 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 qb i2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=2
xmp19 qb ck vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net016 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKINVGTPLT_V7_3




.subckt SAEDRVT14_CKINVGTPLT_V7_4 vdd vss vbp vbn qb ck en se
xmn173 net433 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn172 net432 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn171 net431 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn163 qb ck net433 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn162 qb ck net432 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn161 qb ck net431 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 net43 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn16 qb ck net43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 net016 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 qb i2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmp19 qb ck vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net016 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKINVGTPLT_V7_4




.subckt SAEDRVT14_CKINVGTPLT_V7_5 vdd vss vbp vbn qb ck en se
xmn174 net434 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn173 net433 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn172 net432 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn171 net431 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn164 qb ck net434 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn163 qb ck net433 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn162 qb ck net432 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn161 qb ck net431 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 net43 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn16 qb ck net43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 net016 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 qb i2 vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=2
xmp19 qb ck vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net016 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKINVGTPLT_V7_5




.subckt SAEDRVT14_CKINVGTPLT_V7_6 vdd vss vbp vbn qb ck en se
xmn175 net435 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn174 net434 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn173 net433 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn172 net432 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn171 net431 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn165 qb ck net435 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn164 qb ck net434 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn163 qb ck net433 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn162 qb ck net432 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn161 qb ck net431 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 net43 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn16 qb ck net43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 net016 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 qb i2 vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=2
xmp19 qb ck vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net016 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKINVGTPLT_V7_6




.subckt SAEDRVT14_CKINVGTPLT_V7_8 vdd vss vbp vbn qb ck en se
xmn177 net437 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn176 net436 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn175 net435 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn174 net434 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn173 net433 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn172 net432 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn171 net431 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn167 qb ck net437 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn166 qb ck net436 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn165 qb ck net435 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn164 qb ck net434 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn163 qb ck net433 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn162 qb ck net432 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn161 qb ck net431 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn24 net06 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn17 net43 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn16 qb ck net43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn10 net06 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn23 i1#2fnet61 i2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 net06 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 i1 ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 i2 i1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 net016 se net42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp22 net42 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 qb i2 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=2
xmp19 qb ck vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp21 i1 ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 i1 ckbb net016 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKINVGTPLT_V7_8




.subckt SAEDRVT14_CKSPLT_1 vdd vss vbp vbn ckout ckoutb ck
xmn27 net28 net28 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn22 ckout net7 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn21 net7 ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn20 net31 net29 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn14 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 net014 net010 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 net010 ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn4 ckoutb qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn3 net30 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn2 ckb net014 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn1 ckbb net010 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn0 net31 ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp27 net29 net29 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp20 ckout net7 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp19 net7 ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp18 net30 net28 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp12 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 net014 net010 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 net010 ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp4 ckoutb qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp3 qf ckbb net30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp2 ckb net014 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 ckbb net010 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp0 qf ckb net31 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_CKSPLT_1




.subckt SAEDRVT14_CKSPLT_8 vdd vss vbp vbn ckout ckoutb ck
xmn27 net28 net28 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn22 ckout net7 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn21 net7 ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn20 net31 net29 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn14 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 net014 net010 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn0 net010 ck vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmmn4 ckoutb qf_x vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmmn3 net30 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn2 ckb net014 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn1 ckbb net010 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn0 net31 ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp27 net29 net29 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp20 ckout net7 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp19 net7 ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp18 net30 net28 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp12 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 net014 net010 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp0 net010 ck vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmmp4 ckoutb qf_x vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmmp3 qf ckbb net30 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp2 ckb net014 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 ckbb net010 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 qf ckb net31 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_CKSPLT_8




.subckt SAEDRVT14_DCAP_ECO_12 vdd vss vbp vbn
xmn1 vss net10 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 net8 net10 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn1 vdd net8 vdd vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp1 vdd net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 net10 net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp1 vss net10 vss vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_DCAP_ECO_12




.subckt SAEDRVT14_DCAP_ECO_15 vdd vss vbp vbn
xmn1 vss net10 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn0 net8 net10 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn1 vdd net8 vdd vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp1 vdd net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 net10 net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp1 vss net10 vss vbp p08_rev l=0.014u nf=3 m=1 nfin=2
.ends SAEDRVT14_DCAP_ECO_15




.subckt SAEDRVT14_DCAP_ECO_18 vdd vss vbp vbn
xmn1 vss net10 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn0 net8 net10 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn1 vdd net8 vdd vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmp1 vdd net8 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp0 net10 net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp1 vss net10 vss vbp p08_rev l=0.014u nf=3 m=1 nfin=2
.ends SAEDRVT14_DCAP_ECO_18




.subckt SAEDRVT14_DCAP_ECO_6 vdd vss vbp vbn
xmn0 net8 net10 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn1 vdd net8 vdd vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 net10 net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp1 vss net10 vss vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_DCAP_ECO_6




.subckt SAEDRVT14_DCAP_ECO_9 vdd vss vbp vbn
xmn1 vss net10 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 net8 net10 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn1 vdd net8 vdd vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 net10 net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp1 vss net10 vss vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_DCAP_ECO_9




.subckt SAEDRVT14_DCAP_PV1ECO_12 vdd vss vddr
xn0 net8 net10 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn2 vss net10 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 vddr net8 vddr vss n08_rev l=0.014u nf=2 m=1 nfin=4
xp0 net10 net8 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp2 vddr net8 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 vss net10 vss vddr p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_DCAP_PV1ECO_12




.subckt SAEDRVT14_DCAP_PV1ECO_15 vdd vss vddr
xn0 net8 net10 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn2 vss net10 vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 vddr net8 vddr vss n08_rev l=0.014u nf=2 m=1 nfin=4
xp0 net10 net8 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp2 vddr net8 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 vss net10 vss vddr p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_DCAP_PV1ECO_15




.subckt SAEDRVT14_DCAP_PV1ECO_18 vdd vss vddr
xn0 net8 net10 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn2 vss net10 vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 vddr net8 vddr vss n08_rev l=0.014u nf=3 m=1 nfin=4
xp0 net10 net8 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp2 vddr net8 vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 vss net10 vss vddr p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_DCAP_PV1ECO_18




.subckt SAEDRVT14_DCAP_PV1ECO_6 vdd vss vddr
xn0 net8 net10 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn1 vddr net8 vddr vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp0 net10 net8 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp1 vss net10 vss vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_DCAP_PV1ECO_6




.subckt SAEDRVT14_DCAP_PV1ECO_9 vdd vss vddr
xn0 net8 net10 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn2 vss net10 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 vddr net8 vddr vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp0 net10 net8 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp1 vss net10 vss vddr p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_DCAP_PV1ECO_9




.subckt SAEDRVT14_DCAP_PV3_3 vdd vss vddr
xmn1 net3 net3 net3 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 net3 net3 net3 vss n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_DCAP_PV3_3




.subckt SAEDRVT14_DCAP_V4_16 vdd vss vbp vbn
xmp0 net10 net8 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmmp3 vdd net10 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmn1 vdd net8 vdd vbp p08_rev l=0.014u nf=10 m=1 nfin=2
xmn0 net8 net10 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmmp1 vss net10 vss vbn n08_rev l=0.014u nf=10 m=1 nfin=2
xmmn3 vss net8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_DCAP_V4_16




.subckt SAEDRVT14_DCAP_V4_32 vdd vss vbp vbn
xmp0 net10 net8 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=2
xmmp3 vdd net10 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmn1 vdd net8 vdd vbp p08_rev l=0.014u nf=22 m=1 nfin=2
xmn0 net8 net10 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=2
xmmp1 vss net10 vss vbn n08_rev l=0.014u nf=22 m=1 nfin=2
xmmn3 vss net8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_DCAP_V4_32




.subckt SAEDRVT14_DCAP_V4_5 vdd vss vbp vbn
xmp0 net10 net8 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmmp3 vdd net10 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmn1 vdd net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 net8 net10 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmmp1 vss net10 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn4 vss net8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_DCAP_V4_5




.subckt SAEDRVT14_DCAP_V4_64 vdd vss vbp vbn
xmp0 net10 net8 vdd vbp p08_rev l=0.014u nf=16 m=1 nfin=2
xmmp3 vdd net10 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmn1 vdd net8 vdd vbp p08_rev l=0.014u nf=46 m=1 nfin=2
xmn0 net8 net10 vss vbn n08_rev l=0.014u nf=16 m=1 nfin=2
xmmp1 vss net10 vss vbn n08_rev l=0.014u nf=46 m=1 nfin=2
xmmn3 vss net8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_DCAP_V4_64




.subckt SAEDRVT14_DCAP_V4_8 vdd vss vbp vbn
xmp0 net10 net8 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmmp3 vdd net10 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmn1 vdd net8 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmn0 net8 net10 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmmp1 vss net10 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmmn4 vss net8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_DCAP_V4_8




.subckt SAEDRVT14_DEL_L4D100_1 vdd vss vbp vbn x a
xn18 net22 net_n1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn11 x n3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net_n1 a vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn1 n3 net_n2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 net_n2 net_n1 net22 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xp18 net27 net_n1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp11 x n3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net_n1 a vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 n3 net_n2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net_n2 net_n1 net27 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_DEL_L4D100_1




.subckt SAEDRVT14_DEL_L4D100_2 vdd vss vbp vbn x a
xn18 net22 net_n1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn11 x n3 vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net_n1 a vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn1 n3 net_n2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 net_n2 net_n1 net22 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xp18 net27 net_n1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp11 x n3 vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp2 net_n1 a vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 n3 net_n2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net_n2 net_n1 net27 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_DEL_L4D100_2




.subckt SAEDRVT14_DEL_PR2V2_1 a vbn vbp vdd vddr vss x
xp18 net14 a vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp11 x n1 net010 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp0 n1 a net14 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp2 net010 n1 vddr vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xn18 net13 a vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn11 x n1 net09 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 n1 a net13 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn2 net09 n1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_DEL_PR2V2_1




.subckt SAEDRVT14_DELPROGS4_12 vdd vss vbp vbn x a s0 s1 s2 s3
xmi22#2fn1 net10 net11 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi21#2fn1 net8 net12 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi20#2fn1 net9 net13 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi19#2fn1 net13 net14 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi18#2fn1 i18#2fmidn_en_ck net10 vss vbn n08_rev l=0.014u nf=12 m=1 nfin=4
xmi18#2fn0 x net15 i18#2fmidn_en_ck vbn n08_rev l=0.014u nf=12 m=1 nfin=4
xmi17#2fn1 i17#2fmidn_en_ck net8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi17#2fn0 net11 net16 i17#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fn1 i16#2fmidn_en_ck net9 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fn0 net12 net17 i16#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi15#2fn11 i15#2fmidn_en_ck1 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn01 net15 a i15#2fmidn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn1 i15#2fmidn_en_ck s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn0 net15 a i15#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi14#2fn1 i14#2fmidn_en_ck s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi14#2fn0 net16 a i14#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi13#2fn1 i13#2fmidn_en_ck s2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi13#2fn0 net17 a i13#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi12#2fn1 i12#2fmidn_en_ck s3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi12#2fn0 net14 a i12#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi22#2fp1 net10 net11 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi21#2fp1 net8 net12 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi20#2fp1 net9 net13 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi19#2fp1 net13 net14 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi18#2fp1 x net15 vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmi18#2fp0 x net10 vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmi17#2fp1 net11 net16 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi17#2fp0 net11 net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fp1 net12 net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fp0 net12 net9 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi15#2fp1 net15 a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi15#2fp0 net15 s0 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi14#2fp1 net16 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi14#2fp0 net16 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi13#2fp1 net17 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi13#2fp0 net17 s2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi12#2fp1 net14 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi12#2fp0 net14 s3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_DELPROGS4_12




.subckt SAEDRVT14_DELPROGS4_16 vdd vss vbp vbn x a s0 s1 s2 s3
xmi22#2fn1 net10 net11 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi21#2fn1 net8 net12 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi20#2fn1 net9 net13 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi19#2fn1 net13 net14 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi18#2fn1 i18#2fmidn_en_ck net10 vss vbn n08_rev l=0.014u nf=16 m=1 nfin=4
xmi18#2fn0 x net15 i18#2fmidn_en_ck vbn n08_rev l=0.014u nf=16 m=1 nfin=4
xmi17#2fn1 i17#2fmidn_en_ck net8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi17#2fn0 net11 net16 i17#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fn1 i16#2fmidn_en_ck net9 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fn0 net12 net17 i16#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi15#2fn11 i15#2fmidn_en_ck1 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn01 net15 a i15#2fmidn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn1 i15#2fmidn_en_ck s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn0 net15 a i15#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi14#2fn1 i14#2fmidn_en_ck s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi14#2fn0 net16 a i14#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi13#2fn1 i13#2fmidn_en_ck s2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi13#2fn0 net17 a i13#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi12#2fn1 i12#2fmidn_en_ck s3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi12#2fn0 net14 a i12#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi22#2fp1 net10 net11 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi21#2fp1 net8 net12 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi20#2fp1 net9 net13 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi19#2fp1 net13 net14 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi18#2fp1 x net15 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmi18#2fp0 x net10 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmi17#2fp1 net11 net16 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi17#2fp0 net11 net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fp1 net12 net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fp0 net12 net9 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi15#2fp1 net15 a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi15#2fp0 net15 s0 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi14#2fp1 net16 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi14#2fp0 net16 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi13#2fp1 net17 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi13#2fp0 net17 s2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi12#2fp1 net14 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi12#2fp0 net14 s3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_DELPROGS4_16




.subckt SAEDRVT14_DELPROGS4_4 vdd vss vbp vbn x a s0 s1 s2 s3
xmi22#2fn1 net10 net11 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi21#2fn1 net8 net12 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi20#2fn1 net9 net13 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi19#2fn1 net13 net14 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi18#2fn1 i18#2fmidn_en_ck net10 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi18#2fn0 x net15 i18#2fmidn_en_ck vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmi17#2fn1 i17#2fmidn_en_ck net8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi17#2fn0 net11 net16 i17#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fn1 i16#2fmidn_en_ck net9 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fn0 net12 net17 i16#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi15#2fn11 i15#2fmidn_en_ck1 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn01 net15 a i15#2fmidn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn1 i15#2fmidn_en_ck s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn0 net15 a i15#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi14#2fn1 i14#2fmidn_en_ck s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi14#2fn0 net16 a i14#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi13#2fn1 i13#2fmidn_en_ck s2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi13#2fn0 net17 a i13#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi12#2fn1 i12#2fmidn_en_ck s3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi12#2fn0 net14 a i12#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi22#2fp1 net10 net11 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi21#2fp1 net8 net12 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi20#2fp1 net9 net13 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi19#2fp1 net13 net14 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi18#2fp1 x net15 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi18#2fp0 x net10 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi17#2fp1 net11 net16 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi17#2fp0 net11 net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fp1 net12 net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fp0 net12 net9 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi15#2fp1 net15 a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi15#2fp0 net15 s0 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi14#2fp1 net16 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi14#2fp0 net16 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi13#2fp1 net17 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi13#2fp0 net17 s2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi12#2fp1 net14 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi12#2fp0 net14 s3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_DELPROGS4_4




.subckt SAEDRVT14_DELPROGS4_6 vdd vss vbp vbn x a s0 s1 s2 s3
xmi22#2fn1 net10 net11 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi21#2fn1 net8 net12 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi20#2fn1 net9 net13 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi19#2fn1 net13 net14 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi18#2fn1 i18#2fmidn_en_ck net10 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmi18#2fn0 x net15 i18#2fmidn_en_ck vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmi17#2fn1 i17#2fmidn_en_ck net8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi17#2fn0 net11 net16 i17#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fn1 i16#2fmidn_en_ck net9 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fn0 net12 net17 i16#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi15#2fn11 i15#2fmidn_en_ck1 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn01 net15 a i15#2fmidn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn1 i15#2fmidn_en_ck s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn0 net15 a i15#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi14#2fn1 i14#2fmidn_en_ck s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi14#2fn0 net16 a i14#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi13#2fn1 i13#2fmidn_en_ck s2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi13#2fn0 net17 a i13#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi12#2fn1 i12#2fmidn_en_ck s3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi12#2fn0 net14 a i12#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi22#2fp1 net10 net11 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi21#2fp1 net8 net12 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi20#2fp1 net9 net13 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi19#2fp1 net13 net14 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi18#2fp1 x net15 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmi18#2fp0 x net10 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmi17#2fp1 net11 net16 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi17#2fp0 net11 net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fp1 net12 net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fp0 net12 net9 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi15#2fp1 net15 a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi15#2fp0 net15 s0 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi14#2fp1 net16 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi14#2fp0 net16 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi13#2fp1 net17 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi13#2fp0 net17 s2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi12#2fp1 net14 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi12#2fp0 net14 s3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_DELPROGS4_6




.subckt SAEDRVT14_DELPROGS4_8 vdd vss vbp vbn x a s0 s1 s2 s3
xmi22#2fn1 net10 net11 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi21#2fn1 net8 net12 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi20#2fn1 net9 net13 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi19#2fn1 net13 net14 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi18#2fn1 i18#2fmidn_en_ck net10 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmi18#2fn0 x net15 i18#2fmidn_en_ck vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmi17#2fn1 i17#2fmidn_en_ck net8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi17#2fn0 net11 net16 i17#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fn1 i16#2fmidn_en_ck net9 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fn0 net12 net17 i16#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi15#2fn11 i15#2fmidn_en_ck1 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn01 net15 a i15#2fmidn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn1 i15#2fmidn_en_ck s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi15#2fn0 net15 a i15#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi14#2fn1 i14#2fmidn_en_ck s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi14#2fn0 net16 a i14#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi13#2fn1 i13#2fmidn_en_ck s2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi13#2fn0 net17 a i13#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi12#2fn1 i12#2fmidn_en_ck s3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi12#2fn0 net14 a i12#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi22#2fp1 net10 net11 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi21#2fp1 net8 net12 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi20#2fp1 net9 net13 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi19#2fp1 net13 net14 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi18#2fp1 x net15 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi18#2fp0 x net10 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi17#2fp1 net11 net16 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi17#2fp0 net11 net8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fp1 net12 net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fp0 net12 net9 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi15#2fp1 net15 a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi15#2fp0 net15 s0 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi14#2fp1 net16 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi14#2fp0 net16 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi13#2fp1 net17 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi13#2fp0 net17 s2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi12#2fp1 net14 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi12#2fp0 net14 s3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_DELPROGS4_8




.subckt SAEDRVT14_DELPROGS4_Y2_24 vdd vss vbp vbn x a s0 s1 s2 s3
xmi22#2fn1 net10 net11 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmi21#2fn1 net8 net12 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi20#2fn1 net9 net13 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi19#2fn1 net13 net14 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi18#2fn1 i18#2fmidn_en_ck net10 vss vbn n08_rev l=0.014u nf=22 m=1 nfin=4
xmi18#2fn0 x net15 i18#2fmidn_en_ck vbn n08_rev l=0.014u nf=22 m=1 nfin=4
xmi17#2fn11 i17#2fmidn_en_ck1 net8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi17#2fn01 net11 net16 i17#2fmidn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi17#2fn1 i17#2fmidn_en_ck net8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi17#2fn0 net11 net16 i17#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi16#2fn1 i16#2fmidn_en_ck net9 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fn0 net12 net17 i16#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi15#2fn1 i15#2fmidn_en_ck s0 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi15#2fn0 net15 a i15#2fmidn_en_ck vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi14#2fn1 i14#2fmidn_en_ck s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi14#2fn0 net16 a i14#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi13#2fn1 i13#2fmidn_en_ck s2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi13#2fn0 net17 a i13#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi12#2fn1 i12#2fmidn_en_ck s3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi12#2fn0 net14 a i12#2fmidn_en_ck vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi22#2fp1 net10 net11 vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=4
xmi21#2fp1 net8 net12 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi20#2fp1 net9 net13 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi19#2fp1 net13 net14 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi18#2fp1 x net15 vdd vbp p08_rev l=0.014u nf=12 m=1 nfin=4
xmi18#2fp0 x net10 vdd vbp p08_rev l=0.014u nf=12 m=1 nfin=4
xmi17#2fp1 net11 net16 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi17#2fp0 net11 net8 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi16#2fp1 net12 net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi16#2fp0 net12 net9 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi15#2fp1 net15 a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi15#2fp0 net15 s0 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi14#2fp1 net16 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi14#2fp0 net16 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi13#2fp1 net17 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi13#2fp0 net17 s2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi12#2fp1 net14 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi12#2fp0 net14 s3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_DELPROGS4_Y2_24




.subckt SAEDRVT14_DELPROGS9_V1_4 vdd vss vbp vbn x a s0 s1 s2 s3 s4 s5 s6 s7 s8
xmi9#2fn4 i9#2fnet60 net97 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi9#2fn3 i9#2fnet44 i9#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi9#2fn2 net103 i9#2fnet60 i9#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi9#2fn1 i9#2fnet52 s2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi9#2fn0 i9#2fnet80 net118 i9#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi8#2fn4 i8#2fnet60 net91 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi8#2fn3 i8#2fnet44 i8#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi8#2fn2 net97 i8#2fnet60 i8#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi8#2fn1 i8#2fnet52 s3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi8#2fn0 i8#2fnet80 net118 i8#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi7#2fn4 i7#2fnet60 net85 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi7#2fn3 i7#2fnet44 i7#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi7#2fn2 net91 i7#2fnet60 i7#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi7#2fn1 i7#2fnet52 s4 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi7#2fn0 i7#2fnet80 net118 i7#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi6#2fn4 i6#2fnet60 net79 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi6#2fn3 i6#2fnet44 i6#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi6#2fn2 net85 i6#2fnet60 i6#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi6#2fn1 i6#2fnet52 s5 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi6#2fn0 i6#2fnet80 net118 i6#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi5#2fn4 i5#2fnet60 net73 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi5#2fn3 i5#2fnet44 i5#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi5#2fn2 net79 i5#2fnet60 i5#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi5#2fn1 i5#2fnet52 s6 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi5#2fn0 i5#2fnet80 net118 i5#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi4#2fn4 i4#2fnet60 net67 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi4#2fn3 i4#2fnet44 i4#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi4#2fn2 net73 i4#2fnet60 i4#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi4#2fn1 i4#2fnet52 s7 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi4#2fn0 i4#2fnet80 net118 i4#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi3#2fn4 i3#2fnet60 net126 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn3 i3#2fnet44 i3#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi3#2fn2 net67 i3#2fnet60 i3#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi3#2fn1 i3#2fnet52 s8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fn0 i3#2fnet80 net118 i3#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 net126 i2#2fnet17 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi11#2fn4 i11#2fnet60 net109 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi11#2fn3 i11#2fnet44 i11#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi11#2fn2 net115 i11#2fnet60 i11#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi11#2fn1 i11#2fnet52 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi11#2fn0 i11#2fnet80 net118 i11#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi10#2fn4 i10#2fnet60 net103 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi10#2fn3 i10#2fnet44 i10#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi10#2fn2 net109 i10#2fnet60 i10#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi10#2fn1 i10#2fnet52 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi10#2fn0 i10#2fnet80 net118 i10#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 x net115 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn1 net118 a vss vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmi9#2fp4 i9#2fnet60 net97 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi9#2fp3 net103 i9#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi9#2fp2 net103 i9#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi9#2fp1 i9#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi9#2fp0 i9#2fnet80 s2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi8#2fp4 i8#2fnet60 net91 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi8#2fp3 net97 i8#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi8#2fp2 net97 i8#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi8#2fp1 i8#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi8#2fp0 i8#2fnet80 s3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi7#2fp4 i7#2fnet60 net85 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi7#2fp3 net91 i7#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi7#2fp2 net91 i7#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi7#2fp1 i7#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi7#2fp0 i7#2fnet80 s4 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi6#2fp4 i6#2fnet60 net79 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi6#2fp3 net85 i6#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi6#2fp2 net85 i6#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi6#2fp1 i6#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi6#2fp0 i6#2fnet80 s5 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi5#2fp4 i5#2fnet60 net73 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi5#2fp3 net79 i5#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi5#2fp2 net79 i5#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi5#2fp1 i5#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi5#2fp0 i5#2fnet80 s6 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi4#2fp4 i4#2fnet60 net67 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi4#2fp3 net73 i4#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi4#2fp2 net73 i4#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi4#2fp1 i4#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi4#2fp0 i4#2fnet80 s7 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fp4 i3#2fnet60 net126 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp3 net67 i3#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp2 net67 i3#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 i3#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp0 i3#2fnet80 s8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp0 i2#2fnet17 i2#2fnet17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi11#2fp4 i11#2fnet60 net109 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi11#2fp3 net115 i11#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi11#2fp2 net115 i11#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi11#2fp1 i11#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi11#2fp0 i11#2fnet80 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi10#2fp4 i10#2fnet60 net103 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi10#2fp3 net109 i10#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi10#2fp2 net109 i10#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi10#2fp1 i10#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi10#2fp0 i10#2fnet80 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp1 x net115 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmi0#2fp1 net118 a vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_DELPROGS9_V1_4




.subckt SAEDRVT14_DELPROGS9_V2_4 vdd vss vbp vbn x a s0 s1 s2 s3 s4 s5 s6 s7 s8
xmi9#2fn10 net103 i9#2fnet025 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi9#2fn9 i9#2fnet025 i9#2fnet022 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi9#2fn4 i9#2fnet60 net97 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi9#2fn3 i9#2fnet44 i9#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi9#2fn2 i9#2fnet022 i9#2fnet60 i9#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi9#2fn1 i9#2fnet52 s2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi9#2fn0 i9#2fnet80 net118 i9#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi8#2fn10 net97 i8#2fnet025 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi8#2fn9 i8#2fnet025 i8#2fnet022 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi8#2fn4 i8#2fnet60 net91 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi8#2fn3 i8#2fnet44 i8#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi8#2fn2 i8#2fnet022 i8#2fnet60 i8#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi8#2fn1 i8#2fnet52 s3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi8#2fn0 i8#2fnet80 net118 i8#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi7#2fn10 net91 i7#2fnet025 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi7#2fn9 i7#2fnet025 i7#2fnet022 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi7#2fn4 i7#2fnet60 net85 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi7#2fn3 i7#2fnet44 i7#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi7#2fn2 i7#2fnet022 i7#2fnet60 i7#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi7#2fn1 i7#2fnet52 s4 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi7#2fn0 i7#2fnet80 net118 i7#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi6#2fn10 net85 i6#2fnet025 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi6#2fn9 i6#2fnet025 i6#2fnet022 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi6#2fn4 i6#2fnet60 net79 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi6#2fn3 i6#2fnet44 i6#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi6#2fn2 i6#2fnet022 i6#2fnet60 i6#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi6#2fn1 i6#2fnet52 s5 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi6#2fn0 i6#2fnet80 net118 i6#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi5#2fn10 net79 i5#2fnet025 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi5#2fn9 i5#2fnet025 i5#2fnet022 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi5#2fn4 i5#2fnet60 net73 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi5#2fn3 i5#2fnet44 i5#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi5#2fn2 i5#2fnet022 i5#2fnet60 i5#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi5#2fn1 i5#2fnet52 s6 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi5#2fn0 i5#2fnet80 net118 i5#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi4#2fn10 net73 i4#2fnet025 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi4#2fn9 i4#2fnet025 i4#2fnet022 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi4#2fn4 i4#2fnet60 net67 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi4#2fn3 i4#2fnet44 i4#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi4#2fn2 i4#2fnet022 i4#2fnet60 i4#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi4#2fn1 i4#2fnet52 s7 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi4#2fn0 i4#2fnet80 net118 i4#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi3#2fn10 net67 i3#2fnet025 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fn9 i3#2fnet025 i3#2fnet022 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fn4 i3#2fnet60 net126 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi3#2fn3 i3#2fnet44 i3#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi3#2fn2 i3#2fnet022 i3#2fnet60 i3#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi3#2fn1 i3#2fnet52 s8 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fn0 i3#2fnet80 net118 i3#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 net126 i2#2fnet17 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi11#2fn4 i11#2fnet60 net109 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi11#2fn3 i11#2fnet44 i11#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi11#2fn2 net115 i11#2fnet60 i11#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi11#2fn1 i11#2fnet52 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi11#2fn0 i11#2fnet80 net118 i11#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi10#2fn10 net109 i10#2fnet025 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi10#2fn9 i10#2fnet025 i10#2fnet022 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi10#2fn4 i10#2fnet60 net103 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi10#2fn3 i10#2fnet44 i10#2fnet80 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi10#2fn2 i10#2fnet022 i10#2fnet60 i10#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi10#2fn1 i10#2fnet52 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi10#2fn0 i10#2fnet80 net118 i10#2fnet52 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 x net115 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn1 net118 a vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmi9#2fp10 net103 i9#2fnet025 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi9#2fp9 i9#2fnet025 i9#2fnet022 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi9#2fp4 i9#2fnet60 net97 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi9#2fp3 i9#2fnet022 i9#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi9#2fp2 i9#2fnet022 i9#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi9#2fp1 i9#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi9#2fp0 i9#2fnet80 s2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi8#2fp10 net97 i8#2fnet025 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi8#2fp9 i8#2fnet025 i8#2fnet022 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi8#2fp4 i8#2fnet60 net91 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi8#2fp3 i8#2fnet022 i8#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi8#2fp2 i8#2fnet022 i8#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi8#2fp1 i8#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi8#2fp0 i8#2fnet80 s3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi7#2fp10 net91 i7#2fnet025 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi7#2fp9 i7#2fnet025 i7#2fnet022 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi7#2fp4 i7#2fnet60 net85 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi7#2fp3 i7#2fnet022 i7#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi7#2fp2 i7#2fnet022 i7#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi7#2fp1 i7#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi7#2fp0 i7#2fnet80 s4 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi6#2fp10 net85 i6#2fnet025 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi6#2fp9 i6#2fnet025 i6#2fnet022 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi6#2fp4 i6#2fnet60 net79 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi6#2fp3 i6#2fnet022 i6#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi6#2fp2 i6#2fnet022 i6#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi6#2fp1 i6#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi6#2fp0 i6#2fnet80 s5 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi5#2fp10 net79 i5#2fnet025 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi5#2fp9 i5#2fnet025 i5#2fnet022 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi5#2fp4 i5#2fnet60 net73 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi5#2fp3 i5#2fnet022 i5#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi5#2fp2 i5#2fnet022 i5#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi5#2fp1 i5#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi5#2fp0 i5#2fnet80 s6 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi4#2fp10 net73 i4#2fnet025 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi4#2fp9 i4#2fnet025 i4#2fnet022 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi4#2fp4 i4#2fnet60 net67 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi4#2fp3 i4#2fnet022 i4#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi4#2fp2 i4#2fnet022 i4#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi4#2fp1 i4#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi4#2fp0 i4#2fnet80 s7 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp10 net67 i3#2fnet025 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fp9 i3#2fnet025 i3#2fnet022 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fp4 i3#2fnet60 net126 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi3#2fp3 i3#2fnet022 i3#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi3#2fp2 i3#2fnet022 i3#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi3#2fp1 i3#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi3#2fp0 i3#2fnet80 s8 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp0 i2#2fnet17 i2#2fnet17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi11#2fp4 i11#2fnet60 net109 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi11#2fp3 net115 i11#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi11#2fp2 net115 i11#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi11#2fp1 i11#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi11#2fp0 i11#2fnet80 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi10#2fp10 net109 i10#2fnet025 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi10#2fp9 i10#2fnet025 i10#2fnet022 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi10#2fp4 i10#2fnet60 net103 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi10#2fp3 i10#2fnet022 i10#2fnet60 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi10#2fp2 i10#2fnet022 i10#2fnet80 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi10#2fp1 i10#2fnet80 net118 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi10#2fp0 i10#2fnet80 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp1 x net115 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmi0#2fp1 net118 a vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_DELPROGS9_V2_4




.subckt SAEDRVT14_DEL_R2V1_1 a vbn vbp vdd vss x
xmp18 net14 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp11 x n1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 n1 a net14 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 net13 a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn11 x n1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 n1 a net13 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_DEL_R2V1_1




.subckt SAEDRVT14_DEL_R2V1_2 a vbn vbp vdd vss x
xmp18 net14 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp11 x n1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp0 n1 a net14 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 net13 a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn11 x n1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn0 n1 a net13 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_DEL_R2V1_2




.subckt SAEDRVT14_DEL_R2V2_1 vdd vss vbp vbn x a
xmn18 net15 a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 net18 net_n1 vss vbn n08_rev l=0.014u nf=1 m=2 nfin=4
xmn1 x net_n1 net18 vbn n08_rev l=0.014u nf=1 m=2 nfin=4
xmn0 net_n1 a net15 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp18 net16 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 net17 net_n1 vdd vbp p08_rev l=0.014u nf=1 m=2 nfin=4
xmp1 x net_n1 net17 vbp p08_rev l=0.014u nf=1 m=2 nfin=4
xmp0 net_n1 a net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_DEL_R2V2_1




.subckt SAEDRVT14_DEL_R2V2_2 vdd vss vbp vbn x a
xmn18 net15 a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 net18 net_n1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 x net_n1 net18 vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn0 net_n1 a net15 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp18 net16 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 net17 net_n1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x net_n1 net17 vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp0 net_n1 a net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_DEL_R2V2_2




.subckt SAEDRVT14_DEL_R2V3_1 vdd vss vbp vbn x a
xmn18 net15 a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 net18 net_n1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x net_n1 net18 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 net04 a net15 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn3 net_n1 a net04 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp18 net16 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 net17 net_n1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x net_n1 net17 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 net04 a net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmmp3 net_n1 a net04 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_DEL_R2V3_1




.subckt SAEDRVT14_DEL_R2V3_2 vdd vss vbp vbn x a
xmn21 net181 net_n1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn18 net15 a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn11 x net_n1 net181 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 net18 net_n1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x net_n1 net18 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 net04 a net15 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn3 net_n1 a net04 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp21 net171 net_n1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp18 net16 a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp11 x net_n1 net171 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 net17 net_n1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x net_n1 net17 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 net04 a net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp3 net_n1 a net04 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_DEL_R2V3_2




.subckt SAEDRVT14_ELVLDNOR_V2_10 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=6 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xm2 net36 net27 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddl vddl p08_rev l=0.014u nf=6 m=1 nfin=4
xm6 net40 net36 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=3
xm5 net27 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
xm4 net36 en net17 vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm3 net17 net27 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ELVLDNOR_V2_10




.subckt SAEDRVT14_ELVLDNOR_V2_12 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=7 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xm2 net36 net27 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddl vddl p08_rev l=0.014u nf=7 m=1 nfin=4
xm6 net40 net36 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=3
xm5 net27 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
xm4 net36 en net17 vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm3 net17 net27 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ELVLDNOR_V2_12




.subckt SAEDRVT14_ELVLDNOR_V2_1 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xm7 net40 net36 vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xm2 net36 net27 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=3
xm6 net40 net36 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=3
xm5 net27 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm4 net36 en net17 vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm3 net17 net27 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ELVLDNOR_V2_1




.subckt SAEDRVT14_ELVLDNOR_V2_2 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm7 net40 net36 vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xm2 net36 net27 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=3
xm6 net40 net36 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=3
xm5 net27 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm4 net36 en net17 vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm3 net17 net27 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ELVLDNOR_V2_2




.subckt SAEDRVT14_ELVLDNOR_V2_3 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm2 net36 net27 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xm6 net40 net36 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=3
xm5 net27 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm4 net36 en net17 vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm3 net17 net27 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ELVLDNOR_V2_3




.subckt SAEDRVT14_ELVLDNOR_V2_4 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=3 m=1 nfin=3
xm7 net40 net36 vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xm2 net36 net27 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddl vddl p08_rev l=0.014u nf=3 m=1 nfin=3
xm6 net40 net36 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=3
xm5 net27 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm4 net36 en net17 vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm3 net17 net27 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ELVLDNOR_V2_4




.subckt SAEDRVT14_ELVLDNOR_V2_6 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=4 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xm2 net36 net27 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddl vddl p08_rev l=0.014u nf=4 m=1 nfin=4
xm6 net40 net36 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=3
xm5 net27 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
xm4 net36 en net17 vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm3 net17 net27 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ELVLDNOR_V2_6




.subckt SAEDRVT14_ELVLDNOR_V2_8 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=5 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xm2 net36 net27 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddl vddl p08_rev l=0.014u nf=5 m=1 nfin=4
xm6 net40 net36 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=3
xm5 net27 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
xm4 net36 en net17 vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm3 net17 net27 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ELVLDNOR_V2_8




.subckt SAEDRVT14_ELVLUNOR_V2_10 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=5 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=2
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddh vddh p08_rev l=0.014u nf=5 m=1 nfin=4
xm6 net40 net36 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xm4 net36 en net17 vddl p08_rev l=0.014u nf=3 m=1 nfin=4
xm3 net17 net27 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ELVLUNOR_V2_10




.subckt SAEDRVT14_ELVLUNOR_V2_12 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=6 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=2
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddh vddh p08_rev l=0.014u nf=6 m=1 nfin=4
xm6 net40 net36 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xm4 net36 en net17 vddl p08_rev l=0.014u nf=3 m=1 nfin=4
xm3 net17 net27 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ELVLUNOR_V2_12




.subckt SAEDRVT14_ELVLUNOR_V2_1 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=3 nfin=3
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
xm6 net40 net36 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=3
xm4 net36 en net17 vddl p08_rev l=0.014u nf=3 m=1 nfin=3
xm3 net17 net27 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ELVLUNOR_V2_1




.subckt SAEDRVT14_ELVLUNOR_V2_2 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=2
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
xm6 net40 net36 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xm4 net36 en net17 vddl p08_rev l=0.014u nf=3 m=1 nfin=4
xm3 net17 net27 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ELVLUNOR_V2_2




.subckt SAEDRVT14_ELVLUNOR_V2_3 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=2
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xm6 net40 net36 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xm4 net36 en net17 vddl p08_rev l=0.014u nf=3 m=1 nfin=4
xm3 net17 net27 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ELVLUNOR_V2_3




.subckt SAEDRVT14_ELVLUNOR_V2_4 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=2
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddh vddh p08_rev l=0.014u nf=3 m=1 nfin=3
xm6 net40 net36 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xm4 net36 en net17 vddl p08_rev l=0.014u nf=3 m=1 nfin=4
xm3 net17 net27 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ELVLUNOR_V2_4




.subckt SAEDRVT14_ELVLUNOR_V2_6 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=3 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=2
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddh vddh p08_rev l=0.014u nf=3 m=1 nfin=4
xm6 net40 net36 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xm4 net36 en net17 vddl p08_rev l=0.014u nf=3 m=1 nfin=4
xm3 net17 net27 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ELVLUNOR_V2_6




.subckt SAEDRVT14_ELVLUNOR_V2_8 a en vss x vddh vddl
xm9 x net40 vss vss n08_rev l=0.014u nf=4 m=1 nfin=4
xm7 net40 net36 vss vss n08_rev l=0.014u nf=3 m=1 nfin=2
xm2 net36 net27 vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xm1 net36 en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 net27 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 x net40 vddh vddh p08_rev l=0.014u nf=4 m=1 nfin=4
xm6 net40 net36 vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 net27 a vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xm4 net36 en net17 vddl p08_rev l=0.014u nf=3 m=1 nfin=4
xm3 net17 net27 vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ELVLUNOR_V2_8




.subckt SAEDRVT14_EN2_0P5 vdd vss vbp vbn x a1 a2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi0#2fn3 i0#2fi0#2fbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fi0#2fn1 i0#2fi0#2fbbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fi0#2fp3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 a1 i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_EN2_0P5




.subckt SAEDRVT14_EN2_1P5 vdd vss vbp vbn x a1 a2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi0#2fi0#2fndummy vss a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn3 i0#2fi0#2fbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn1 i0#2fi0#2fbbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fi0#2fp3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 a1 i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_EN2_1P5




.subckt SAEDRVT14_EN2_1 vdd vss vbp vbn x a1 a2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi0#2fn3 i0#2fi0#2fbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi0#2fi0#2fn1 i0#2fi0#2fbbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 a1 i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_EN2_1




.subckt SAEDRVT14_EN2_2 vdd vss vbp vbn x a1 a2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn5 vss a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn3 i0#2fi0#2fbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn1 i0#2fi0#2fbbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 a1 i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_EN2_2




.subckt SAEDRVT14_EN2_3 vdd vss vbp vbn x a1 a2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmi0#2fi0#2fndummy vss a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn3 i0#2fi0#2fbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn1 i0#2fi0#2fbbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmi0#2fi0#2fp3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 a1 i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_EN2_3




.subckt SAEDRVT14_EN2_4 vdd vss vbp vbn x a1 a2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn4 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fi0#2fn3 i0#2fi0#2fbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fi0#2fn1 i0#2fi0#2fbbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp4 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fi0#2fp3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fi0#2fp1 i0#2fi0#2fnet17 a1 i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp0 i0#2fi0#2fnet17 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_EN2_4




.subckt SAEDRVT14_EN2_ECO_1 vdd vss vbp vbn x a1 a2
xmn5 ab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 bb a1 int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 bb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 bbb ab int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 bbb bb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp5 ab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 bb ab int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 bb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 net21 a1 int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 net21 bb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_EN2_ECO_1




.subckt SAEDRVT14_EN2_V1_0P75 vdd vss vbp vbn x a1 a2
xn5 x1 a2 midn_a1a2_b1nrb2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn3 x1 a1 midn_a1a2_b1nrb2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 midn_a1a2_b1nrb2 b1nrb2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn1 midn_b1_b2 a2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn0 b1nrb2 a1 midn_b1_b2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 midp_b1_b2 a2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp4 x1 b1nrb2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 x1 a1 midp_b1_b2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 b1nrb2 a1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp0 b1nrb2 a2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_EN2_V1_0P75




.subckt SAEDRVT14_EN2_V1_1P5 vdd vss vbp vbn x a1 a2
xn5 x1 a2 midn_a1a2_b1nrb2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn3 x1 a1 midn_a1a2_b1nrb2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 midn_a1a2_b1nrb2 b1nrb2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn1 midn_b1_b2 a2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn0 b1nrb2 a1 midn_b1_b2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 midp_b1_b2 a2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp4 x1 b1nrb2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 x1 a1 midp_b1_b2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 b1nrb2 a1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp0 b1nrb2 a2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_EN2_V1_1P5




.subckt SAEDRVT14_EN3_1 vdd vss vbp vbn x a1 a2 a3
xmmn12 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn11 c_xn_b c_xr_b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn10 bb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn3 i1#2fbb c_xr_b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn2 i1#2fbb a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn1 i1#2fbbb c_xn_b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 i1#2fbbb i1#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fbb a2 c_xr_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn2 i0#2fbb a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn1 i0#2fbbb bb c_xr_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 i0#2fbbb i0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmp12 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp11 c_xn_b c_xr_b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp10 bb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp3 i1#2fbb c_xn_b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp2 i1#2fbb a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp1 i1#2fnet21 c_xr_b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 i1#2fnet21 i1#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fbb bb c_xr_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fbb a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp1 i0#2fnet21 a2 c_xr_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet21 i0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_EN3_1




.subckt SAEDRVT14_EN3_2 vdd vss vbp vbn x a1 a2 a3
xmmn12 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn11 c_xn_b c_xr_b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn10 bb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn3 i1#2fbb c_xr_b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn2 i1#2fbb a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 i1#2fbbb c_xn_b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn0 i1#2fbbb i1#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn3 i0#2fbb a2 c_xr_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn2 i0#2fbb a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn1 i0#2fbbb bb c_xr_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 i0#2fbbb i0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpdummy vdd a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp12 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp11 c_xn_b c_xr_b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp10 bb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp3 i1#2fbb c_xn_b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp2 i1#2fbb a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 i1#2fnet21 c_xr_b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp0 i1#2fnet21 i1#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fbb bb c_xr_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fbb a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp1 i0#2fnet21 a2 c_xr_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet21 i0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_EN3_2




.subckt SAEDRVT14_EN3_3 vdd vss vbp vbn x a1 a2 a3
xmmn12 x int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmmn11 c_xn_b c_xr_b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn10 bb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn3 i1#2fbb c_xr_b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn2 i1#2fbb a1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 i1#2fbbb c_xn_b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn0 i1#2fbbb i1#2fbb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn3 i0#2fbb a2 c_xr_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn2 i0#2fbb a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1 i0#2fbbb bb c_xr_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 i0#2fbbb i0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmp13 vdd a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp12 x int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmmp11 c_xn_b c_xr_b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp10 bb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp3 i1#2fbb c_xn_b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp2 i1#2fbb a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 i1#2fnet21 c_xr_b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp0 i1#2fnet21 i1#2fbb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp3 i0#2fbb bb c_xr_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 i0#2fbb a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1 i0#2fnet21 a2 c_xr_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0 i0#2fnet21 i0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_EN3_3




.subckt SAEDRVT14_EN3_U_0P5 vdd vss vbp vbn x a1 a2 a3
xmmn12 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn11 net8 net1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn10 bb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn3 net3 net1 int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn2 net3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn1 net4 net8 int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 net4 net3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 net2 a2 net1 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn2 net2 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn1 net6 bb net1 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 net6 net2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmp12 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp11 net8 net1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp10 bb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp3 net3 net8 int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp2 net3 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp1 net5 net1 int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 net5 net3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 net2 bb net1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 net2 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp1 net7 a2 net1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 net7 net2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_EN3_U_0P5




.subckt SAEDRVT14_EN4_2 vdd vss vbp vbn x a1 a2 a3 a4
xn10 x int_zn vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn9 a_xr_b c_xn_d int_zn vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn8 a_xn_b c_xr_d int_zn vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn5 ab a1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn4 a_xn_b a_xr_b vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn16 c_xn_d c_xr_d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn15 cb a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xi1#2fn3 i1#2fbb a3 c_xr_d vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn2 i1#2fbb a4 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn1 i1#2fbbb cb c_xr_d vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn0 i1#2fbbb i1#2fbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn3 i0#2fbb a1 a_xr_b vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn2 i0#2fbb a2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn1 i0#2fbbb ab a_xr_b vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn0 i0#2fbbb i0#2fbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xp12 a_xr_b c_xr_d int_zn vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp11 a_xn_b c_xn_d int_zn vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp9 x int_zn vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp5 ab a1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp4 a_xn_b a_xr_b vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp16 c_xn_d c_xr_d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp15 cb a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xi1#2fp3 i1#2fbb cb c_xr_d vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp2 i1#2fbb a4 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp1 i1#2fnet21 a3 c_xr_d vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp0 i1#2fnet21 i1#2fbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp3 i0#2fbb ab a_xr_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp2 i0#2fbb a2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp1 i0#2fnet21 a1 a_xr_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp0 i0#2fnet21 i0#2fbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
.ends SAEDRVT14_EN4_2




.subckt SAEDRVT14_FDN_V2_4 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet030 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xqn7 qn qf vss vbn n08 l=0.014u nf=4 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_FDN_V2_4



.subckt SAEDRVT14_FDN8_V2_4 ck d1 d2 d3 d4 d5 d6 d7 do q1 q2 q3 q4 q5 q6 q7 qn1 qn2 qn3 qn4 qn5 qn6 qn7 qno qo vbn vbp vdd vss
xi5 vdd vss vbp vbn q7 qn7 ck d7 SAEDRVT14_FDN_V2_4
xi4 vdd vss vbp vbn q6 qn6 ck d6 SAEDRVT14_FDN_V2_4
xi3 vdd vss vbp vbn q5 qn5 ck d5 SAEDRVT14_FDN_V2_4
xi2 vdd vss vbp vbn q4 qn4 ck d4 SAEDRVT14_FDN_V2_4
xi1 vdd vss vbp vbn q3 qn3 ck d3 SAEDRVT14_FDN_V2_4
xi0 vdd vss vbp vbn q2 qn2 ck d2 SAEDRVT14_FDN_V2_4
xsaedrvt14_fdn8_v2_4 vdd vss vbp vbn q1 qn1 ck d1 SAEDRVT14_FDN_V2_4
xhdbsvt14_fdn2_v2_2_0 vdd vss vbp vbn qo qno ck do SAEDRVT14_FDN_V2_4
.ends SAEDRVT14_FDN8_V2_4




.subckt SAEDRVT14_EN4_M_1 vdd vss vbp vbn x a1 a2 a3 a4
xmn10 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn9 a_xr_b c_xn_d int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn8 a_xn_b c_xr_d int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 ab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 a_xn_b a_xr_b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn16 c_xn_d c_xr_d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn15 cb a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn3 i1#2fbb a3 c_xr_d vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn2 i1#2fbb a4 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 i1#2fbbb cb c_xr_d vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn0 i1#2fbbb i1#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fbb a1 a_xr_b vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fbb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1 i0#2fbbb ab a_xr_b vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fbbb i0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp12 a_xr_b c_xr_d int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp11 a_xn_b c_xn_d int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp9 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp5 ab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 a_xn_b a_xr_b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp16 c_xn_d c_xr_d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp15 cb a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp3 i1#2fbb cb c_xr_d vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp2 i1#2fbb a4 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 i1#2fnet21 a3 c_xr_d vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 i1#2fnet21 i1#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fbb ab a_xr_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fbb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1 i0#2fnet21 a1 a_xr_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp0 i0#2fnet21 i0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_EN4_M_1




.subckt SAEDRVT14_EN4_U_0P5 vdd vss vbp vbn x a1 a2 a3 a4
xn10 x int_zn vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn9 a_xr_b c_xn_d int_zn vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn8 a_xn_b c_xr_d int_zn vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn5 ab a1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn4 a_xn_b a_xr_b vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xmn16 c_xn_d c_xr_d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn15 cb a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xi1#2fn3 i1#2fbb a3 c_xr_d vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn2 i1#2fbb a4 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn1 i1#2fbbb cb c_xr_d vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn0 i1#2fbbb i1#2fbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn3 i0#2fbb a1 a_xr_b vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn2 i0#2fbb a2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn1 i0#2fbbb ab a_xr_b vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn0 i0#2fbbb i0#2fbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xp12 a_xr_b c_xr_d int_zn vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp11 a_xn_b c_xn_d int_zn vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp9 x int_zn vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp5 ab a1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp4 a_xn_b a_xr_b vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xmp16 c_xn_d c_xr_d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp15 cb a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xi1#2fp3 i1#2fbb cb c_xr_d vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp2 i1#2fbb a4 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp1 i1#2fnet21 a3 c_xr_d vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp0 i1#2fnet21 i1#2fbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp3 i0#2fbb ab a_xr_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp2 i0#2fbb a2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp1 i0#2fnet21 a1 a_xr_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp0 i0#2fnet21 i0#2fbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
.ends SAEDRVT14_EN4_U_0P5




.subckt SAEDRVT14_EO2_0P5 vdd vss vbp vbn x a1 a2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fn3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fn1 i0#2fi0#2fbbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fp3 i0#2fi0#2fbb a1 i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_EO2_0P5




.subckt SAEDRVT14_EO2_1P5 vdd vss vbp vbn x a1 a2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi0#2fi0#2fndummy vss a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn1 i0#2fi0#2fbbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi0#2fi0#2fp3 i0#2fi0#2fbb a1 i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_EO2_1P5




.subckt SAEDRVT14_EO2_1 vdd vss vbp vbn x a1 a2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fn1 i0#2fi0#2fbbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp3 i0#2fi0#2fbb a1 i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_EO2_1




.subckt SAEDRVT14_EO2_2 vdd vss vbp vbn x a1 a2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fi0#2fndummy vss a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn1 i0#2fi0#2fbbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fi0#2fp3 i0#2fi0#2fbb a1 i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_EO2_2




.subckt SAEDRVT14_EO2_3 vdd vss vbp vbn x a1 a2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmi0#2fi0#2fndummy vss a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn1 i0#2fi0#2fbbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmi0#2fi0#2fp3 i0#2fi0#2fbb a1 i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_EO2_3




.subckt SAEDRVT14_EO2_4 vdd vss vbp vbn x a1 a2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fi0#2fn3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn1 i0#2fi0#2fbbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fi0#2fp3 i0#2fi0#2fbb a1 i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_EO2_4




.subckt SAEDRVT14_EO2_ECO_1 vdd vss vbp vbn x a1 a2
xmn8 x int_zn yn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn7 yn int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn6 int_zn x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 ab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 x1 int_zn1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 int_zn1 ab bb vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 bb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 int_zn1 a1 bbb vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 bbb bb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp8 x int_zn yp vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp7 yp int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp6 int_zn x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 ab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 x1 int_zn1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 int_zn1 a1 bb vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 bb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 int_zn1 ab net28 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 net28 bb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_EO2_ECO_1




.subckt SAEDRVT14_EO2_MM_0P5 vdd vss vbp vbn x a1 a2
xmn8 x int_zn yn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn7 yn int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn6 int_zn x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 x1 i0#2fint_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn1 i0#2fi0#2fbbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp8 x int_zn yp vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp7 yp int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp6 int_zn x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 x1 i0#2fint_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi0#2fp3 i0#2fi0#2fbb a1 i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_EO2_MM_0P5




.subckt SAEDRVT14_EO2_MM_1 vdd vss vbp vbn x a1 a2
xmn8 x int_zn yn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn7 yn int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn6 int_zn x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 x1 i0#2fint_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fn1 i0#2fi0#2fbbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp8 x int_zn yp vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp7 yp int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp6 int_zn x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 x1 i0#2fint_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fi0#2fp3 i0#2fi0#2fbb a1 i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_EO2_MM_1




.subckt SAEDRVT14_EO2_MM_2 vdd vss vbp vbn x a1 a2
xmn8 x int_zn yn vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn7 yn int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn6 int_zn x1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn4 x1 i0#2fint_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fi0#2fn3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fi0#2fn1 i0#2fi0#2fbbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmp8 x int_zn yp vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp7 yp int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp6 int_zn x1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp4 x1 i0#2fint_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi0#2fi0#2fp3 i0#2fi0#2fbb a1 i0#2fint_zn vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_EO2_MM_2




.subckt SAEDRVT14_EO2_MM_4 vdd vss vbp vbn x a1 a2
xmn8 x int_zn yn vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn7 yn int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn6 int_zn x1 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmi0#2fn5 i0#2fab a1 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmi0#2fn4 x1 i0#2fint_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fi0#2fn3 i0#2fi0#2fbb i0#2fab i0#2fint_zn vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmi0#2fi0#2fn2 i0#2fi0#2fbb a2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fi0#2fn1 i0#2fi0#2fbbb a1 i0#2fint_zn vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmi0#2fi0#2fn0 i0#2fi0#2fbbb i0#2fi0#2fbb vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmp8 x int_zn yp vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp7 yp int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp6 int_zn x1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmi0#2fp5 i0#2fab a1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmi0#2fp4 x1 i0#2fint_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmi0#2fi0#2fp3 i0#2fi0#2fbb a1 i0#2fint_zn vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmi0#2fi0#2fp2 i0#2fi0#2fbb a2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fi0#2fp1 i0#2fi0#2fnet21 i0#2fab i0#2fint_zn vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fi0#2fp0 i0#2fi0#2fnet21 i0#2fi0#2fbb vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_EO2_MM_4




.subckt SAEDRVT14_EO2_V1_0P75 vdd vss vbp vbn x a1 a2
xn5 midn_a1_a2 a2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn4 x b1ndb2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn3 x a1 midn_a1_a2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn1 b1ndb2 a1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 b1ndb2 a2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp5 x a2 midp_a1a2_b1ndb2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 x a1 midp_a1a2_b1ndb2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 midp_a1a2_b1ndb2 b1ndb2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 midp_b1_b2 a2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp0 b1ndb2 a1 midp_b1_b2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_EO2_V1_0P75




.subckt SAEDRVT14_EO2_V1_1P5 vdd vss vbp vbn x a1 a2
xn51 midn_a1_a21 a2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn31 x a1 midn_a1_a21 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn5 midn_a1_a2 a2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn4 x b1ndb2 vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=2
xn3 x a1 midn_a1_a2 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn1 b1ndb2 a1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 b1ndb2 a2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp5 x a2 midp_a1a2_b1ndb2 vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 x a1 midp_a1a2_b1ndb2 vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp2 midp_a1a2_b1ndb2 b1ndb2 vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp1 midp_b1_b2 a2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp0 b1ndb2 a1 midp_b1_b2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_EO2_V1_1P5




.subckt SAEDRVT14_EO3_0P5 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn12 x1 int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn11 c_xr_b c_xn_b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn10 bb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn3 i1#2fbb c_xn_b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn2 i1#2fbb a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn1 i1#2fbbb c_xr_b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn0 i1#2fbbb i1#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fbb bb c_xn_b vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fbb a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 i0#2fbbb a2 c_xn_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 i0#2fbbb i0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmmp12 x1 int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp11 c_xr_b c_xn_b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp10 bb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp3 i1#2fbb c_xr_b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp2 i1#2fbb a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp1 i1#2fnet21 c_xn_b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 i1#2fnet21 i1#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fbb a2 c_xn_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fbb a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 i0#2fnet21 bb c_xn_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet21 i0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_EO3_0P5




.subckt SAEDRVT14_EO3_1 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn12 x1 int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn11 c_xr_b c_xn_b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn10 bb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn3 i1#2fbb c_xn_b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn2 i1#2fbb a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn1 i1#2fbbb c_xr_b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn0 i1#2fbbb i1#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fbb bb c_xn_b vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fbb a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 i0#2fbbb a2 c_xn_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 i0#2fbbb i0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmmp12 x1 int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp11 c_xr_b c_xn_b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp10 bb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp3 i1#2fbb c_xr_b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp2 i1#2fbb a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp1 i1#2fnet21 c_xn_b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 i1#2fnet21 i1#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fbb a2 c_xn_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fbb a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 i0#2fnet21 bb c_xn_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet21 i0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_EO3_1




.subckt SAEDRVT14_EO3_2 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn12 x1 int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn11 c_xr_b c_xn_b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn10 bb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn3 i1#2fbb c_xn_b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn2 i1#2fbb a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn1 i1#2fbbb c_xr_b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn0 i1#2fbbb i1#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fbb bb c_xn_b vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fbb a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 i0#2fbbb a2 c_xn_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 i0#2fbbb i0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmmp12 x1 int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp11 c_xr_b c_xn_b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp10 bb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp3 i1#2fbb c_xr_b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp2 i1#2fbb a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp1 i1#2fnet21 c_xn_b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 i1#2fnet21 i1#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fbb a2 c_xn_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fbb a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 i0#2fnet21 bb c_xn_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet21 i0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_EO3_2




.subckt SAEDRVT14_EO3_4 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn12 x1 int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn11 c_xr_b c_xn_b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn10 bb a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn3 i1#2fbb c_xn_b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn2 i1#2fbb a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn1 i1#2fbbb c_xr_b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn0 i1#2fbbb i1#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fbb bb c_xn_b vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fbb a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 i0#2fbbb a2 c_xn_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 i0#2fbbb i0#2fbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmmp12 x1 int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp11 c_xr_b c_xn_b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp10 bb a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp3 i1#2fbb c_xr_b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp2 i1#2fbb a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp1 i1#2fnet21 c_xn_b int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 i1#2fnet21 i1#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fbb a2 c_xn_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fbb a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 i0#2fnet21 bb c_xn_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet21 i0#2fbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_EO3_4




.subckt SAEDRVT14_EO4_1 vdd vss vbp vbn x a1 a2 a3 a4
xn10 x int_zn vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn9 a_xn_b c_xn_d int_zn vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn8 a_xr_b c_xr_d int_zn vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn5 ab a1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn4 a_xn_b a_xr_b vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xmn16 c_xn_d c_xr_d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn15 cb a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xi1#2fn3 i1#2fbb a3 c_xr_d vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn2 i1#2fbb a4 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn1 i1#2fbbb cb c_xr_d vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn0 i1#2fbbb i1#2fbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn3 i0#2fbb a1 a_xr_b vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn2 i0#2fbb a2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn1 i0#2fbbb ab a_xr_b vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn0 i0#2fbbb i0#2fbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xp12 a_xn_b c_xr_d int_zn vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp11 a_xr_b c_xn_d int_zn vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp9 x int_zn vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp5 ab a1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp4 a_xn_b a_xr_b vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xmp16 c_xn_d c_xr_d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp15 cb a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xi1#2fp3 i1#2fbb cb c_xr_d vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp2 i1#2fbb a4 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp1 i1#2fnet21 a3 c_xr_d vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp0 i1#2fnet21 i1#2fbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp3 i0#2fbb ab a_xr_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp2 i0#2fbb a2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp1 i0#2fnet21 a1 a_xr_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp0 i0#2fnet21 i0#2fbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
.ends SAEDRVT14_EO4_1




.subckt SAEDRVT14_EO4_2 vdd vss vbp vbn x a1 a2 a3 a4
xn10 x int_zn vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn9 a_xn_b c_xn_d int_zn vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn8 a_xr_b c_xr_d int_zn vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn5 ab a1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn4 a_xn_b a_xr_b vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xmn16 c_xn_d c_xr_d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn15 cb a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xi1#2fn3 i1#2fbb a3 c_xr_d vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn2 i1#2fbb a4 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn1 i1#2fbbb cb c_xr_d vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn0 i1#2fbbb i1#2fbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn3 i0#2fbb a1 a_xr_b vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn2 i0#2fbb a2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn1 i0#2fbbb ab a_xr_b vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn0 i0#2fbbb i0#2fbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xp12 a_xn_b c_xr_d int_zn vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp11 a_xr_b c_xn_d int_zn vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp9 x int_zn vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp5 ab a1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp4 a_xn_b a_xr_b vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xmp16 c_xn_d c_xr_d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp15 cb a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xi1#2fp3 i1#2fbb cb c_xr_d vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp2 i1#2fbb a4 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp1 i1#2fnet21 a3 c_xr_d vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp0 i1#2fnet21 i1#2fbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp3 i0#2fbb ab a_xr_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp2 i0#2fbb a2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp1 i0#2fnet21 a1 a_xr_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp0 i0#2fnet21 i0#2fbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_EO4_2




.subckt SAEDRVT14_EO4_4 vdd vss vbp vbn x a1 a2 a3 a4
xn10 x int_zn vss vbn n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn9 a_xn_b c_xn_d int_zn vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn8 a_xr_b c_xr_d int_zn vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn5 ab a1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn4 a_xn_b a_xr_b vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xmn16 c_xn_d c_xr_d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn15 cb a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xi1#2fn3 i1#2fbb a3 c_xr_d vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn2 i1#2fbb a4 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn1 i1#2fbbb cb c_xr_d vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn0 i1#2fbbb i1#2fbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn3 i0#2fbb a1 a_xr_b vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn2 i0#2fbb a2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn1 i0#2fbbb ab a_xr_b vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn0 i0#2fbbb i0#2fbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xp12 a_xn_b c_xr_d int_zn vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp11 a_xr_b c_xn_d int_zn vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp9 x int_zn vdd vbp p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp5 ab a1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp4 a_xn_b a_xr_b vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xmp16 c_xn_d c_xr_d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp15 cb a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xi1#2fp3 i1#2fbb cb c_xr_d vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp2 i1#2fbb a4 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp1 i1#2fnet21 a3 c_xr_d vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp0 i1#2fnet21 i1#2fbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp3 i0#2fbb ab a_xr_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp2 i0#2fbb a2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp1 i0#2fnet21 a1 a_xr_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp0 i0#2fnet21 i0#2fbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_EO4_4




.subckt SAEDRVT14_EO4_U_0P5 vdd vss vbp vbn x a1 a2 a3 a4
xn10 x1 int_zn1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn9 a_xn_b c_xn_d int_zn1 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn8 a_xr_b c_xr_d int_zn1 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn5 ab a1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn4 a_xn_b a_xr_b vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=3
xmn16 c_xn_d c_xr_d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn15 cb a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn8 x int_zn yn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn7 yn int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn6 int_zn x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xi1#2fn3 i1#2fbb a3 c_xr_d vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn2 i1#2fbb a4 vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=3   
xi1#2fn1 i1#2fbbb cb c_xr_d vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn0 i1#2fbbb i1#2fbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn3 i0#2fbb a1 a_xr_b vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn2 i0#2fbb a2 vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=3   
xi0#2fn1 i0#2fbbb ab a_xr_b vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn0 i0#2fbbb i0#2fbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xp12 a_xn_b c_xr_d int_zn1 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp11 a_xr_b c_xn_d int_zn1 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp9 x1 int_zn1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp5 ab a1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp4 a_xn_b a_xr_b vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=3
xmp16 c_xn_d c_xr_d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp15 cb a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp8 x int_zn yp vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp7 yp int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp6 int_zn x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xi1#2fp3 i1#2fbb cb c_xr_d vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp2 i1#2fbb a4 vdd vbp p08_rev3 l=0.014u nf=2 m=1 nfin=3   
xi1#2fp1 i1#2fnet21 a3 c_xr_d vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp0 i1#2fnet21 i1#2fbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp3 i0#2fbb ab a_xr_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp2 i0#2fbb a2 vdd vbp p08_rev3 l=0.014u nf=2 m=1 nfin=3   
xi0#2fp1 i0#2fnet21 a1 a_xr_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp0 i0#2fnet21 i0#2fbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
.ends SAEDRVT14_EO4_U_0P5


SAEDRVT14_FDN_V2_0P5

.subckt SAEDRVT14_FDN_V2_0P5 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDN_V2_0P5

.subckt SAEDRVT14_FDN2_V2_0P5 vdd vss vbp vbn q0 q1 qn1 ck d0 d1 qno
xhdbsvt14_fdn2_v2_0p5_1 vdd vss vbp vbn q1 qn1 ck d1 SAEDRVT14_FDN_V2_0P5
xhdbsvt14_fdn2_v2_0p5_0 vdd vss vbp vbn q0 qno ck d0 SAEDRVT14_FDN_V2_0P5
.ends SAEDRVT14_FDN2_V2_0P5




.subckt SAEDRVT14_FDN_V2_1 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FDN_V2_1



.subckt SAEDRVT14_FDN2_V2_1 vdd vss vbp vbn q0 q1 qn0 qn1 ck d0 d1
xi1 vdd vss vbp vbn q1 qn1 ck d1 SAEDRVT14_FDN_V2_1
xi0 vdd vss vbp vbn q0 qn0 ck d0 SAEDRVT14_FDN_V2_1
.ends SAEDRVT14_FDN2_V2_1




.subckt SAEDRVT14_FDN_V2_1 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet027 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_FDN_V2_1

.subckt SAEDRVT14_FDN2_V2_2 vdd vss vbp vbn q0 q1 qn0 qn1 ck d0 d1
xi1 vdd vss vbp vbn q1 qn1 ck d1 SAEDRVT14_FDN_V2_1
xi0 vdd vss vbp vbn q0 qn0 ck d0 SAEDRVT14_FDN_V2_1
.ends SAEDRVT14_FDN2_V2_2




.subckt SAEDRVT14_FDN_V2_4 vdd vss vbp vbn q qn ck d
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xqn7 qn qf vss vbn n08 l=0.014u nf=4 m=1 nfin=4
xmibase#2fn0 ibase#2fnet030 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn6 mq_x ckbb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp4 mq_x ckb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FDN_V2_4

.subckt SAEDRVT14_FDN2_V2_4 vdd vss vbp vbn q0 q1 qn0 qn1 ck d1 do
xhdbsvt14_fdn2_v2_2_1 vdd vss vbp vbn q1 qn1 ck d1 SAEDRVT14_FDN_V2_4
xhdbsvt14_fdn2_v2_2_0 vdd vss vbp vbn q0 qn0 ck do SAEDRVT14_FDN_V2_4
.ends SAEDRVT14_FDN2_V2_4




.subckt SAEDRVT14_FDN_V2_0P5 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDN_V2_0P5

.subckt SAEDRVT14_FDN4_V2_0P5 vdd vss vbp vbn q1 qn0 qn1 ck d0 d1 d2 d3 q2 q3 qn2 qn3 qo
xi3 vdd vss vbp vbn q3 qn3 ck d3 SAEDRVT14_FDN_V2_0P5
xi2 vdd vss vbp vbn q2 qn2 ck d2 SAEDRVT14_FDN_V2_0P5
xhdbsvt14_fdsaedrvt14_fdn4_v2_0p5n2_v2_0p5_1 vdd vss vbp vbn q1 qn1 ck d1 SAEDRVT14_FDN_V2_0P5
xsaedrvt14_fdn4_v2_0p5 vdd vss vbp vbn qo qn0 ck d0 SAEDRVT14_FDN_V2_0P5
.ends SAEDRVT14_FDN4_V2_0P5




.subckt SAEDRVT14_FDN_V2_1 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FDN_V2_1

.subckt SAEDRVT14_FDN4_V2_1 vdd vss vbp vbn q0 q1 qn0 qn1 ck d0 d1 d2 d3 q2 q3 qn2 qn3
xi1 vdd vss vbp vbn q3 qn3 ck d3 SAEDRVT14_FDN_V2_1
xi0 vdd vss vbp vbn q2 qn2 ck d2 SAEDRVT14_FDN_V2_1
xsaedrvt14_fdn4_v2_1 vdd vss vbp vbn q1 qn1 ck d1 SAEDRVT14_FDN_V2_1
xhdbsvt14_fdn2_v2_1_0 vdd vss vbp vbn q0 qn0 ck d0 SAEDRVT14_FDN_V2_1
.ends SAEDRVT14_FDN4_V2_1




.subckt SAEDRVT14_FDN_V2_2 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xm0 ibase#2fnet030 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_FDN_V2_2

.subckt SAEDRVT14_FDN4_V2_2 vdd vss vbp vbn q0 q1 qn0 qn1 ck d0 d1 d2 d3 q2 q3 qn2 qn3
xi6 vdd vss vbp vbn q0 qn0 ck d0 SAEDRVT14_FDN_V2_2
xi7 vdd vss vbp vbn q1 qn1 ck d1 SAEDRVT14_FDN_V2_2
xi8 vdd vss vbp vbn q2 qn2 ck d2 SAEDRVT14_FDN_V2_2
xi9 vdd vss vbp vbn q3 qn3 ck d3 SAEDRVT14_FDN_V2_2
.ends SAEDRVT14_FDN4_V2_2




.subckt SAEDRVT14_FDN_V2_4 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet030 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xqn7 qn qf vss vbn n08 l=0.014u nf=4 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_FDN_V2_4

.subckt SAEDRVT14_FDN4_V2_4 ck d0 d1 d2 d3 q0 q1 q2 q3 qn0 qn1 qn2 qn3 vbn vbp vdd vss
xi5 vdd vss vbp vbn q3 qn3 ck d3 SAEDRVT14_FDN_V2_4
xi4 vdd vss vbp vbn q2 qn2 ck d2 SAEDRVT14_FDN_V2_4
xi3 vdd vss vbp vbn q1 qn1 ck d1 SAEDRVT14_FDN_V2_4
xi2 vdd vss vbp vbn q0 qn0 ck d0 SAEDRVT14_FDN_V2_4
.ends SAEDRVT14_FDN4_V2_4




.subckt SAEDRVT14_FDN_V2_0P5 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDN_V2_0P5

.subckt SAEDRVT14_FDN8_V2_0P5 vdd vss vbp vbn q0 q1 qn0 qn1 ck d0 d1 d2 d3 d4 d5 d6 d7 q2 q3 q4 q5 q6 q7 qn2 qn3 qn4 qn5 qn6 qn7
xi6 vdd vss vbp vbn q0 qn0 ck d0 SAEDRVT14_FDN_V2_0P5
xi7 vdd vss vbp vbn q1 qn1 ck d1 SAEDRVT14_FDN_V2_0P5
xi8 vdd vss vbp vbn q2 qn2 ck d2 SAEDRVT14_FDN_V2_0P5
xi9 vdd vss vbp vbn q3 qn3 ck d3 SAEDRVT14_FDN_V2_0P5
xi10 vdd vss vbp vbn q4 qn4 ck d4 SAEDRVT14_FDN_V2_0P5
xi11 vdd vss vbp vbn q5 qn5 ck d5 SAEDRVT14_FDN_V2_0P5
xi12 vdd vss vbp vbn q6 qn6 ck d6 SAEDRVT14_FDN_V2_0P5
xi13 vdd vss vbp vbn q7 qn7 ck d7 SAEDRVT14_FDN_V2_0P5
.ends SAEDRVT14_FDN8_V2_0P5




.subckt SAEDRVT14_FDN_V2_1 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FDN_V2_1

.subckt SAEDRVT14_FDN8_V2_1 vdd vss vbp vbn q1 qn1 ck d1 d2 d3 d4 d5 d6 d7 do q2 q3 q4 q5 q6 q7 qn2 qn3 qn4 qn5 qn6 qn7 qno qo
xi5 vdd vss vbp vbn q7 qn7 ck d7 SAEDRVT14_FDN_V2_1
xi4 vdd vss vbp vbn q6 qn6 ck d6 SAEDRVT14_FDN_V2_1
xi3 vdd vss vbp vbn q5 qn5 ck d5 SAEDRVT14_FDN_V2_1
xi2 vdd vss vbp vbn q4 qn4 ck d4 SAEDRVT14_FDN_V2_1
xio vdd vss vbp vbn q3 qn3 ck d3 SAEDRVT14_FDN_V2_1
xi0 vdd vss vbp vbn q2 qn2 ck d2 SAEDRVT14_FDN_V2_1
xsaedrvt14_fdn8_v2_1 vdd vss vbp vbn q1 qn1 ck d1 SAEDRVT14_FDN_V2_1
xhdbsvt14_fdn2_v2_1_0 vdd vss vbp vbn qo qno ck do SAEDRVT14_FDN_V2_1
.ends SAEDRVT14_FDN8_V2_1




.subckt SAEDRVT14_FDN_V2_2 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xm0 ibase#2fnet030 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_FDN_V2_2

.subckt SAEDRVT14_FDN8_V2_2 vdd vss vbp vbn q0 q1 qn0 qn1 ck d0 d1 d2 d3 d4 d5 d6 d7 q2 q3 q4 q5 q6 q7 qn2 qn3 qn4 qn5 qn6 qn7
xi5 vdd vss vbp vbn q7 qn7 ck d7 SAEDRVT14_FDN_V2_2
xi4 vdd vss vbp vbn q6 qn6 ck d6 SAEDRVT14_FDN_V2_2
xi3 vdd vss vbp vbn q5 qn5 ck d5 SAEDRVT14_FDN_V2_2
xi2 vdd vss vbp vbn q4 qn4 ck d4 SAEDRVT14_FDN_V2_2
xi1 vdd vss vbp vbn q3 qn3 ck d3 SAEDRVT14_FDN_V2_2
xi0 vdd vss vbp vbn q2 qn2 ck d2 SAEDRVT14_FDN_V2_2
xhdbsvt14_fdn2_v2_2_1 vdd vss vbp vbn q1 qn1 ck d1 SAEDRVT14_FDN_V2_2
xhdbsvt14_fdn2_v2_2_0 vdd vss vbp vbn q0 qn0 ck d0 SAEDRVT14_FDN_V2_2
.ends SAEDRVT14_FDN8_V2_2




.subckt SAEDRVT14_FDN8_V2_4 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet030 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xqn7 qn qf vss vbn n08 l=0.014u nf=4 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_FDN8_V2_4

.subckt SAEDRVT14_FDN8_V2_4 ck d1 d2 d3 d4 d5 d6 d7 do q1 q2 q3 q4 q5 q6 q7 qn1 qn2 qn3 qn4 qn5 qn6 qn7 qno qo vbn vbp vdd vss
xi5 vdd vss vbp vbn q7 qn7 ck d7 SAEDRVT14_FDN_V2_4
xi4 vdd vss vbp vbn q6 qn6 ck d6 SAEDRVT14_FDN_V2_4
xi3 vdd vss vbp vbn q5 qn5 ck d5 SAEDRVT14_FDN_V2_4
xi2 vdd vss vbp vbn q4 qn4 ck d4 SAEDRVT14_FDN_V2_4
xi1 vdd vss vbp vbn q3 qn3 ck d3 SAEDRVT14_FDN_V2_4
xi0 vdd vss vbp vbn q2 qn2 ck d2 SAEDRVT14_FDN_V2_4
xsaedrvt14_fdn8_v2_4 vdd vss vbp vbn q1 qn1 ck d1 SAEDRVT14_FDN_V2_4
xhdbsvt14_fdn2_v2_2_0 vdd vss vbp vbn qo qno ck do SAEDRVT14_FDN_V2_4
.ends SAEDRVT14_FDN8_V2_4




.subckt SAEDRVT14_FDNQ_V2_8 vdd vss vbp vbn q ck d
xmn1 net17 net13 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn0 net13 ck vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmmn2 ckb net17 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn1 ckbb net13 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fsltn1 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf ckbb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fn7 mq_x d ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq_x ckb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmn17 ibase#2fnet31 ckbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmp1 net17 net13 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp0 net13 ck vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmmp2 ckb net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 ckbb net13 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fsltp1 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf ckb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp5 ibase#2fnet41 ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq_x ckbb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp17 mq_x d ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
.ends SAEDRVT14_FDNQ_V2_8




.subckt SAEDRVT14_FDNQ_V3_1 vdd vss vbp vbn q ck d
xmibase#2fsltn1 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 qf ckbb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn16 ibase#2fnet28 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn7 mq_x d ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq_x ckb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn18 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fsltp1 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf ckb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp5 ibase#2fnet41 ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp19 mq_x ckbb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp18 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp17 mq_x d ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_FDNQ_V3_1




.subckt SAEDRVT14_FDNQ_V3_2 vdd vss vbp vbn q ck d
xmibase#2fsltn1 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 qf ckbb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn16 ibase#2fnet28 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn7 mq_x d ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq_x ckb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn18 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fsltp1 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf ckb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp5 ibase#2fnet41 ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp19 mq_x ckbb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp18 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp17 mq_x d ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_FDNQ_V3_2




.subckt SAEDRVT14_FDNQ_V3_4 vdd vss vbp vbn q ck d
xmibase#2fsltn1 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf ckbb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fn7 mq_x d ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq_x ckb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmn17 ibase#2fnet31 ckbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fsltp1 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf ckb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp5 ibase#2fnet41 ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq_x ckbb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp17 mq_x d ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_FDNQ_V3_4




.subckt SAEDRVT14_FDNRBSBQ_V2_0P5 vdd vss vbp vbn q ck d rd sd
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn8 i2 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet038 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet038 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn1 i1 ckbb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 net10 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet016 ckbb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckb ibase#2fnet026 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 ibase#2fnet026 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 i98 ckbb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 ibase#2fnet026 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 i1 ckb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net11 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDNRBSBQ_V2_0P5




.subckt SAEDRVT14_FDNRBSBQ_V2_1 vdd vss vbp vbn q ck d rd sd
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn8 i2 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet038 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet038 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn1 i1 ckbb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 net10 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet016 ckbb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckb ibase#2fnet026 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 ibase#2fnet026 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 i98 ckbb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 ibase#2fnet026 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 i1 ckb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net11 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDNRBSBQ_V2_1




.subckt SAEDRVT14_FDNRBSBQ_V2_2 vdd vss vbp vbn q ck d rd sd
xmibase#2fn9_1 ibase#2fnet43_1 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn2_1 i99 i98 ibase#2fnet43_1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn8 i2 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet027 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet027 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn1 i1 ckbb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 net10 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet016 ckbb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckb ibase#2fnet026 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 ibase#2fnet026 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 i98 ckbb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 ibase#2fnet026 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 i1 ckb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net11 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDNRBSBQ_V2_2




.subckt SAEDRVT14_FDNRBSBQ_V2_4 vdd vss vbp vbn q ck d rd sd
xmibase#2fn9_1 ibase#2fnet43_1 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn2_1 i99 i98 ibase#2fnet43_1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn8 i2 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet027 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet027 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn1 i1 ckbb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 net10 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet016 ckbb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckb ibase#2fnet026 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 ibase#2fnet026 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 i98 ckbb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 ibase#2fnet026 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 i1 ckb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net11 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDNRBSBQ_V2_4




.subckt SAEDRVT14_FDN_V2_0P5 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDN_V2_0P5




.subckt SAEDRVT14_FDN_V2_1 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FDN_V2_1




.subckt SAEDRVT14_FDN_V2_2 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet030 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_FDN_V2_2




.subckt SAEDRVT14_FDN_V2_4 vdd vss vbp vbn q qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fn6 mq_x ckbb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet030 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 qn qf vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fp4 mq_x ckb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_FDN_V2_2




.subckt SAEDRVT14_FDPCBQ_V2_0P5 vdd vss vbp vbn q ck d rs
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net10 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 net10 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 net10 rs vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net7 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn14 i0#2fnet23 rs vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 net7 d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPCBQ_V2_0P5




.subckt SAEDRVT14_FDPCBQ_V2_1 vdd vss vbp vbn q ck d rs
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net7 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn14 i0#2fnet23 rs vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 net7 d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net10 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 net10 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 net10 rs vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPCBQ_V2_1




.subckt SAEDRVT14_FDPCBQ_V2_2 vdd vss vbp vbn q ck d rs
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net7 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn14 i0#2fnet23 rs vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 net7 d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net10 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 net10 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 net10 rs vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPCBQ_V2_2




.subckt SAEDRVT14_FDPCBQ_V2_4 vdd vss vbp vbn q ck d rs
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net10 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 net10 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 net10 rs vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fn6 mq_x ckb net7 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn14 i0#2fnet23 rs vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 net7 d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPCBQ_V2_4




.subckt SAEDRVT14_FDPCBQ_V2LP_0P5 vdd vss vbp vbn q ck d rs
xmn1 ckbb ckb vss vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq mq_x vss vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net7 vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq ckbb qf vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet23 rs vss vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 net7 d i0#2fnet23 vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net10 vbp p08_lvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf ckb mq vbp p08_lvt l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 net10 d vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 net10 rs vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPCBQ_V2LP_0P5




.subckt SAEDRVT14_FDPCBQ_V2LP_1 vdd vss vbp vbn q ck d rs
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net10 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp12 net10 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 net10 rs vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net7 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn14 i0#2fnet23 rs vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 net7 d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPCBQ_V2LP_1




.subckt SAEDRVT14_FDPCBQ_V2LP_2 vdd vss vbp vbn q ck d rs
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net10 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp12 net10 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 net10 rs vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net7 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn14 i0#2fnet23 rs vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 net7 d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPCBQ_V2LP_2




.subckt SAEDRVT14_FDPCBQ_V3_1 vdd vss vbp vbn q ck d rs
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf_x ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp1 net049 rs vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 qf_x ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn1 net049 d i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn0 i0#2fmidn_a_b rs vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FDPCBQ_V3_1




.subckt SAEDRVT14_FDPCBQ_V3_2 vdd vss vbp vbn q ck d rs
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp14 qf_x ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp1 net049 rs vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf_x ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn1 net049 d i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn0 i0#2fmidn_a_b rs vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FDPCBQ_V3_2




.subckt SAEDRVT14_FDPCBQ_V3_4 vdd vss vbp vbn q ck d rs
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp14 qf_x ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=2 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp1 net049 rs vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf_x ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn1 net049 d i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn0 i0#2fmidn_a_b rs vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FDPCBQ_V3_4




.subckt SAEDRVT14_FDPMQ_0P5 vdd vss vbp vbn q ck d0 d1 s
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 net51 net68 net53 net52 n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 net48 net67 net50 net49 n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 net45 net66 net47 net46 n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 net42 net65 net44 net43 n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 net39 net64 net41 net40 n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 net36 net63 net38 net37 n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 net33 net62 net35 net34 n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 net30 net61 net32 net31 n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 net27 net60 net29 net28 n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 i0#2fseb i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 s i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net050 s i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net050 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPMQ_0P5




.subckt SAEDRVT14_FDPMQ_1 vdd vss vbp vbn q ck d0 d1 s
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net050 s i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net050 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 i0#2fseb i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 s i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPMQ_1




.subckt SAEDRVT14_FDPMQ_2 vdd vss vbp vbn q ck d0 d1 s
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net050 s i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net050 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet030 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 i0#2fseb i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 s i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPMQ_2




.subckt SAEDRVT14_FDPMQ_4 vdd vss vbp vbn q ck d0 d1 s
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fp15 i0#2fseb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net050 s i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net050 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet030 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fn17 i0#2fseb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 i0#2fseb i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 s i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPMQ_4




.subckt SAEDRVT14_FDPQB_V2_1 vdd vss vbp vbn qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FDPQB_V2_1




.subckt SAEDRVT14_FDPQB_V2_2 vdd vss vbp vbn qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_FDPQB_V2_2




.subckt SAEDRVT14_FDPQB_V2_4 vdd vss vbp vbn qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet030 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_FDPQB_V2_4




.subckt SAEDRVT14_FDPQB_V2_8 vdd vss vbp vbn qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn0 ibase#2fnet030 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
.ends SAEDRVT14_FDPQB_V2_8




.subckt SAEDRVT14_FDPQB_V2LP_0P5 vdd vss vbp vbn qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPQB_V2LP_0P5




.subckt SAEDRVT14_FDPQB_V2LP_1 vdd vss vbp vbn qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FDPQB_V2LP_1




.subckt SAEDRVT14_FDPQB_V2LP_2 vdd vss vbp vbn qn ck d
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_FDPQB_V2LP_2




.subckt SAEDRVT14_FDPQB_V3_1 vdd vss vbp vbn qn ck d
xmibase#2fsltn1 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 qf ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn16 ibase#2fnet28 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq_x d ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq_x ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn18 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fsltp1 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq_x ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp17 mq_x d ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_FDPQB_V3_1




.subckt SAEDRVT14_FDPQB_V3_2 vdd vss vbp vbn qn ck d
xmibase#2fsltn1 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq_x d ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn20 mq_x ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fsltp1 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp15 ibase#2fnet27 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp14 qf ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq_x ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp17 mq_x d ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_FDPQB_V3_2




.subckt SAEDRVT14_FDPQB_V3_4 vdd vss vbp vbn qn ck d
xmibase#2fsltn1 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq_x d ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmn20 mq_x ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fsltp1 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp15 ibase#2fnet27 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp14 qf ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq_x ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp17 mq_x d ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_FDPQB_V3_4




.subckt SAEDRVT14_FDPQB_V3_8 vdd vss vbp vbn qn ck d
xmibase#2fsltn1 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq_x d ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmn20 mq_x ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fsltp1 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp15 ibase#2fnet27 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp14 qf ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq_x ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp17 mq_x d ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_FDPQB_V3_8




.subckt SAEDRVT14_FDPQ_V2_1 vdd vss vbp vbn q ck d
xmn1 net17 net13 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 net13 ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn2 ckb net17 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn1 ckbb net13 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltn1 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 qf ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn16 ibase#2fnet28 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn7 mq_x d ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq_x ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn18 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 net17 net13 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 net13 ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp2 ckb net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 ckbb net13 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltp1 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp19 mq_x ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp18 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp17 mq_x d ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FDPQ_V2_1




.subckt SAEDRVT14_FDPQ_V2_6 vdd vss vbp vbn q ck d
xmn20 q qf_x vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn18 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn14 d ckb mq vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn13 net31 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn12 mq ckbb net29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn11 net29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 mq_x mq vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn9 qf_x ckb net31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp18 q qf_x vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp16 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp12 mq ckbb d vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp11 net32 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp10 mq ckb net30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp9 net30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp8 mq_x mq vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=2
xmp7 qf_x ckbb net32 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_FDPQ_V2_6




.subckt SAEDRVT14_FDPQ_V2_8 vdd vss vbp vbn q ck d
xmn1 net17 net13 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn0 net13 ck vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmmn2 ckb net17 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn1 ckbb net13 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fsltn1 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fn7 mq_x d ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq_x ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmp1 net17 net13 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp0 net13 ck vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmmp2 ckb net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 ckbb net13 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fsltp1 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq_x ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp17 mq_x d ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
.ends SAEDRVT14_FDPQ_V2_8




.subckt SAEDRVT14_FDPQ_V2ECO_1 vdd vss vbp vbn q ck d
xmn13 net32 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 mq_x ckbb net34 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn11 net34 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn9 qf ckb net32 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn6 mq_x ckb net35 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 net35 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn1 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp11 net31 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp10 mq_x ckb net33 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp9 net33 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp7 qf ckbb net31 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 mq_x ckbb net36 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 net36 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FDPQ_V2ECO_1




.subckt SAEDRVT14_FDPQ_V3_1 vdd vss vbp vbn q ck d
xmibase#2fsltn1 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 qf ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn7 mq_x d ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq_x ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fsltp1 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp14 qf ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq_x ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp17 mq_x d ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_FDPQ_V3_1




.subckt SAEDRVT14_FDPQ_V3_2 vdd vss vbp vbn q ck d
xmibase#2fsltn1 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 qf ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn16 ibase#2fnet28 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn7 mq_x d ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq_x ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn18 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fsltp1 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp19 mq_x ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp18 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp17 mq_x d ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_FDPQ_V3_2




.subckt SAEDRVT14_FDPQ_V3_4 vdd vss vbp vbn q ck d
xmibase#2fsltn1 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fn7 mq_x d ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq_x ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fsltp1 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq_x ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp17 mq_x d ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_FDPQ_V3_4




.subckt SAEDRVT14_FDPRBQ_V2_0P5 vdd vss vbp vbn q ck d rd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPRBQ_V2_0P5




.subckt SAEDRVT14_FDPRBQ_V2_1 vdd vss vbp vbn q ck d rd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 net050 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPRBQ_V2_1




.subckt SAEDRVT14_FDPRBQ_V2_2 vdd vss vbp vbn q ck d rd
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp1 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn0 net050 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPRBQ_V2_2




.subckt SAEDRVT14_FDPRBQ_V2_4 vdd vss vbp vbn q ck d rd
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fp1 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fn0 net050 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPRBQ_V2_4




.subckt SAEDRVT14_FDPRBQ_V2LP_0P5 vdd vss vbp vbn q ck d rd
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPRBQ_V2LP_0P5




.subckt SAEDRVT14_FDPRBQ_V2LP_1 vdd vss vbp vbn q ck d rd
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 net050 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPRBQ_V2LP_1




.subckt SAEDRVT14_FDPRBQ_V2LP_2 vdd vss vbp vbn q ck d rd
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp1 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn0 net050 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPRBQ_V2LP_2




.subckt SAEDRVT14_FDPRBSBQ_V2_0P5 vdd vss vbp vbn q ck d rd sd
xmibase#2fp26 ibase#2fnet016 ckb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckbb ibase#2fnet026 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 ibase#2fnet026 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 i98 ckb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 ibase#2fnet026 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 i1 ckbb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net11 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn8 i2 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet038 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet038 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn1 i1 ckb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 net10 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPRBSBQ_V2_0P5




.subckt SAEDRVT14_FDPRBSBQ_V2_1 vdd vss vbp vbn q ck d rd sd
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn8 i2 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet038 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet038 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn1 i1 ckb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 net10 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet016 ckb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckbb ibase#2fnet026 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 ibase#2fnet026 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 i98 ckb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 ibase#2fnet026 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 i1 ckbb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net11 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPRBSBQ_V2_1




.subckt SAEDRVT14_FDPRBSBQ_V2_2 vdd vss vbp vbn q ck d rd sd
xmibase#2fp26 ibase#2fnet016 ckb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckbb ibase#2fnet026 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 ibase#2fnet026 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 i98 ckb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 ibase#2fnet026 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 i1 ckbb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net11 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9_1 ibase#2fnet43_1 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn2_1 i99 i98 ibase#2fnet43_1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn8 i2 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet027 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet027 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn1 i1 ckb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 net10 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPRBSBQ_V2_2




.subckt SAEDRVT14_FDPRBSBQ_V2_4 vdd vss vbp vbn q ck d rd sd
xmibase#2fn9_1 ibase#2fnet43_1 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn2_1 i99 i98 ibase#2fnet43_1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn8 i2 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet027 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet027 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn1 i1 ckb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 net10 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet016 ckb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckbb ibase#2fnet026 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 ibase#2fnet026 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 i98 ckb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 ibase#2fnet026 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 i1 ckbb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net11 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPRBSBQ_V2_4




.subckt SAEDRVT14_FDPRB_V3_2 vdd vss vbp vbn q qn ck d rd
xmibase#2fsltn1 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn32 ibase#2fnet025 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn31 ibase#2fnet025 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn30 ibase#2fnet025 reseth vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn7 mq_x d ibase#2fnet038 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn21 mq reseth vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmn20 mq_x ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet038 ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi30#2fn0 reseth rd vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi29#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fsltp1 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp31 qf ckbb ibase#2fnet025 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp30 ibase#2fnet035 reseth vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp29 ibase#2fnet025 qf_x ibase#2fnet035 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp5 ibase#2fnet037 ckbb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp21 ibase#2fnet033 reseth vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq_x ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq mq_x ibase#2fnet033 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp17 mq_x d ibase#2fnet037 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi30#2fp1 reseth rd vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi29#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_FDPRB_V3_2




.subckt SAEDRVT14_FDPSBQ_0P5 vdd vss vbp vbn q ck d sd
xmibase#2fp23 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp22 ibase#2fnet025 ckbb qf vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp20 mq sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp19 ibase#2fnet025 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet025 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp10 mq_x ckb ibase#2fnet31 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet31 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn25 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn24 ibase#2fnet24 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet33 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn22 mq mq_x ibase#2fnet33 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 ibase#2fnet30 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet24 qf_x ibase#2fnet30 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet32 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 net050 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPSBQ_0P5




.subckt SAEDRVT14_FDPSBQ_1 vdd vss vbp vbn q ck d sd
xmibase#2fp23 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp22 ibase#2fnet025 ckbb qf vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp20 mq sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp19 ibase#2fnet025 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet025 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp10 mq_x ckb ibase#2fnet31 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet31 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn25 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn24 ibase#2fnet24 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet33 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn22 mq mq_x ibase#2fnet33 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 ibase#2fnet30 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet24 qf_x ibase#2fnet30 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet32 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 net050 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPSBQ_1




.subckt SAEDRVT14_FDPSBQ_2 vdd vss vbp vbn q ck d sd
xmibase#2fn25 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn24 ibase#2fnet24 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet33 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn22 mq mq_x ibase#2fnet33 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 ibase#2fnet30 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn13 ibase#2fnet24 qf_x ibase#2fnet30 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn12 mq_x ckbb ibase#2fnet32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet32 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 net050 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp23 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp22 ibase#2fnet025 ckbb qf vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp20 mq sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp19 ibase#2fnet025 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp11 ibase#2fnet025 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp10 mq_x ckb ibase#2fnet31 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet31 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPSBQ_2




.subckt SAEDRVT14_FDPSBQ_4 vdd vss vbp vbn q ck d sd
xmibase#2fp23 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp22 ibase#2fnet025 ckbb qf vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp20 mq sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp19 ibase#2fnet025 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp11 ibase#2fnet025 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp10 mq_x ckb ibase#2fnet31 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet31 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn25 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn24 ibase#2fnet24 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet33 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn22 mq mq_x ibase#2fnet33 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 ibase#2fnet30 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn13 ibase#2fnet24 qf_x ibase#2fnet30 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn12 mq_x ckbb ibase#2fnet32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet32 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 net050 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPSBQ_4




.subckt SAEDRVT14_FDPSQB_2 ck d qn sd vbn vbp vdd vss
xmibase#2fp23 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp22 ibase#2fnet025 ckbb qf vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp20 mq net06 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp19 ibase#2fnet025 net06 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet025 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp10 mq_x ckb ibase#2fnet31 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet31 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi29#2fp1 net06 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net049 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn25 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn24 ibase#2fnet24 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet33 net06 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn22 mq mq_x ibase#2fnet33 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 ibase#2fnet30 net06 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet24 qf_x ibase#2fnet30 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet32 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi29#2fn0 net06 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 net050 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPSQB_2




.subckt SAEDRVT14_FDPS_V3_2 vdd vss vbp vbn q qn ck d s
xmibase#2fsltn1 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn32 ibase#2fnet025 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn31 ibase#2fnet025 qf_x ibase#2fnet031 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn30 ibase#2fnet031 set vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn7 mq_x d ibase#2fnet038 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn21_2 ibase#2fnet032_2 set vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn18_2 mq mq_x ibase#2fnet032_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn21 ibase#2fnet032 set vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn20 mq_x ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq mq_x ibase#2fnet032 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet038 ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi30#2fn0 set s vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi29#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fsltp1 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp31 qf ckbb ibase#2fnet025 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp30 ibase#2fnet025 set vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp29 ibase#2fnet025 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp5 ibase#2fnet037 ckbb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp21 mq set vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq_x ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp17 mq_x d ibase#2fnet037 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi30#2fp1 set s vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi29#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_FDPS_V3_2




.subckt SAEDRVT14_FDPSYNSBQ_V2_0P5 vdd vss vbp vbn q ck d sd
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net12 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnet011 i0#2fsnb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 net12 d i0#2fnet011 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp12 i0#2fsnb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net9 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn14 net9 i0#2fsnb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 net9 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn12 i0#2fsnb sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPSYNSBQ_V2_0P5




.subckt SAEDRVT14_FDPSYNSBQ_V2_1 vdd vss vbp vbn q ck d sd
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net12 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnet011 i0#2fsnb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 net12 d i0#2fnet011 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp12 i0#2fsnb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net9 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn14 net9 i0#2fsnb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 net9 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn12 i0#2fsnb sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPSYNSBQ_V2_1




.subckt SAEDRVT14_FDPSYNSBQ_V2_2 vdd vss vbp vbn q ck d sd
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net12 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnet011 i0#2fsnb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 net12 d i0#2fnet011 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp12 i0#2fsnb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net9 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn14 net9 i0#2fsnb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 net9 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn12 i0#2fsnb sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPSYNSBQ_V2_2




.subckt SAEDRVT14_FDPSYNSBQ_V2_4 vdd vss vbp vbn q ck d sd
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net12 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnet011 i0#2fsnb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 net12 d i0#2fnet011 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp12 i0#2fsnb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fn6 mq_x ckb net9 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn14 net9 i0#2fsnb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 net9 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn12 i0#2fsnb sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDPSYNSBQ_V2_4




.subckt SAEDRVT14_FDP_V2_0P5 VDD VSS VBP VBN Q QN CK D
Mxmn1 ckbb ckb VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 ckb CK VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn13 ibase#2fnet046 qf_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn12 mq_x ckbb ibase#2fnet048 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn11 ibase#2fnet048 mq VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn10 mq mq_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn9 qf ckb ibase#2fnet046 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn8 qf_x qf VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn6 mq_x ckb ibase#2fnet028 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn5 mq ckbb qf VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn0 ibase#2fnet028 D VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi3#2fn0 QN qf VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi2#2fn0 Q qf_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp1 ckbb ckb VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 ckb CK VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp11 ibase#2fnet045 qf_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp10 mq_x ckb ibase#2fnet047 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp9 ibase#2fnet047 mq VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp8 mq mq_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp7 qf ckbb ibase#2fnet045 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp6 qf_x qf VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp4 mq_x ckbb ibase#2fnet027 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp3 qf ckb mq VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp1 ibase#2fnet027 D VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi3#2fp1 QN qf VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi2#2fp1 Q qf_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDP_V2_0P5




.subckt SAEDRVT14_FDP_V2_1 VDD VSS VBP VBN Q QN CK D
Mxmn1 ckbb ckb VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 ckb CK VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn13 ibase#2fnet046 qf_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn12 mq_x ckbb ibase#2fnet048 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn11 ibase#2fnet048 mq VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn10 mq mq_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn9 qf ckb ibase#2fnet046 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn8 qf_x qf VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn6 mq_x ckb ibase#2fnet028 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn5 mq ckbb qf VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn0 ibase#2fnet028 D VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi3#2fn0 QN qf VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi2#2fn0 Q qf_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 ckbb ckb VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 ckb CK VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp11 ibase#2fnet045 qf_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp10 mq_x ckb ibase#2fnet047 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp9 ibase#2fnet047 mq VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp8 mq mq_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp7 qf ckbb ibase#2fnet045 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp6 qf_x qf VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp4 mq_x ckbb ibase#2fnet027 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp3 qf ckb mq VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp1 ibase#2fnet027 D VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi3#2fp1 QN qf VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi2#2fp1 Q qf_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FDP_V2_1




.subckt SAEDRVT14_FDP_V2_2 VDD VSS VBP VBN Q QN CK D
Mxmn1 ckbb ckb VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 ckb CK VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn13 ibase#2fnet046 qf_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn12 mq_x ckbb ibase#2fnet048 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn11 ibase#2fnet048 mq VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn10 mq mq_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn9 qf ckb ibase#2fnet046 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn8 qf_x qf VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmibase#2fn6 mq_x ckb ibase#2fnet030 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn5 mq ckbb qf VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn0 ibase#2fnet030 D VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi3#2fn0 QN qf VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmi2#2fn0 Q qf_x VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmp1 ckbb ckb VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 ckb CK VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp11 ibase#2fnet045 qf_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp10 mq_x ckb ibase#2fnet047 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp9 ibase#2fnet047 mq VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp8 mq mq_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp7 qf ckbb ibase#2fnet045 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp6 qf_x qf VDD VBP p08 l=0.014u nf=2 m=1 nfin=2
Mxmibase#2fp4 mq_x ckbb ibase#2fnet029 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp3 qf ckb mq VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmibase#2fp1 ibase#2fnet029 D VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi3#2fp1 QN qf VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmi2#2fp1 Q qf_x VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_FDP_V2_2




.subckt SAEDRVT14_FDP_V2_4 VDD VSS VBP VBN Q QN CK D
Mxmn1 ckbb ckb VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 ckb CK VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn13 ibase#2fnet046 qf_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn12 mq_x ckbb ibase#2fnet048 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn11 ibase#2fnet048 mq VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn10 mq mq_x VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmibase#2fn9 qf ckb ibase#2fnet046 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn8 qf_x qf VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmibase#2fn6 mq_x ckb ibase#2fnet030 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn5 mq ckbb qf VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn0 ibase#2fnet030 D VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi3#2fn0 QN qf VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmi2#2fn0 Q qf_x VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmp1 ckbb ckb VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 ckb CK VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp11 ibase#2fnet045 qf_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp10 mq_x ckb ibase#2fnet047 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp9 ibase#2fnet047 mq VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp8 mq mq_x VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmibase#2fp7 qf ckbb ibase#2fnet045 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp6 qf_x qf VDD VBP p08 l=0.014u nf=2 m=1 nfin=2
Mxmibase#2fp4 mq_x ckbb ibase#2fnet029 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp3 qf ckb mq VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmibase#2fp1 ibase#2fnet029 D VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi3#2fp1 QN qf VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmi2#2fp1 Q qf_x VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_FDP_V2_4




.subckt SAEDRVT14_FDP_V2LP_0P5 VDD VSS VBP VBN Q QN CK D
Mxmn1 ckbb ckb VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn0 ckb CK VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn13 ibase#2fnet046 qf_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn12 mq_x ckbb ibase#2fnet048 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn11 ibase#2fnet048 mq VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn10 mq mq_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn9 qf ckb ibase#2fnet046 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn8 qf_x qf VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn6 mq_x ckb ibase#2fnet028 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn5 mq ckbb qf VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn0 ibase#2fnet028 D VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi3#2fn0 QN qf VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi2#2fn0 Q qf_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp1 ckbb ckb VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 ckb CK VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp11 ibase#2fnet045 qf_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp10 mq_x ckb ibase#2fnet047 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp9 ibase#2fnet047 mq VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp8 mq mq_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp7 qf ckbb ibase#2fnet045 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp6 qf_x qf VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp4 mq_x ckbb ibase#2fnet027 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp3 qf ckb mq VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp1 ibase#2fnet027 D VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi3#2fp1 QN qf VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi2#2fp1 Q qf_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FDP_V2LP_0P5




.subckt SAEDRVT14_FDP_V2LP_1 VDD VSS VBP VBN Q QN CK D
Mxmn1 ckbb ckb VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn0 ckb CK VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn13 ibase#2fnet046 qf_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn12 mq_x ckbb ibase#2fnet048 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn11 ibase#2fnet048 mq VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn10 mq mq_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn9 qf ckb ibase#2fnet046 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn8 qf_x qf VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn6 mq_x ckb ibase#2fnet028 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn5 mq ckbb qf VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn0 ibase#2fnet028 D VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi3#2fn0 QN qf VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmi2#2fn0 Q qf_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 ckbb ckb VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 ckb CK VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp11 ibase#2fnet045 qf_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp10 mq_x ckb ibase#2fnet047 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp9 ibase#2fnet047 mq VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp8 mq mq_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp7 qf ckbb ibase#2fnet045 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp6 qf_x qf VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp4 mq_x ckbb ibase#2fnet027 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp3 qf ckb mq VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp1 ibase#2fnet027 D VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi3#2fp1 QN qf VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmi2#2fp1 Q qf_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FDP_V2LP_1




.subckt SAEDRVT14_FDP_V2LP_2 VDD VSS VBP VBN Q QN CK D
Mxmn1 ckbb ckb VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn0 ckb CK VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn13 ibase#2fnet046 qf_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn12 mq_x ckbb ibase#2fnet048 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn11 ibase#2fnet048 mq VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn10 mq mq_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn9 qf ckb ibase#2fnet046 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn8 qf_x qf VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn6 mq_x ckb ibase#2fnet028 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn5 mq ckbb qf VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn0 ibase#2fnet028 D VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmi3#2fn0 QN qf VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmi2#2fn0 Q qf_x VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmp1 ckbb ckb VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp0 ckb CK VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp11 ibase#2fnet045 qf_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp10 mq_x ckb ibase#2fnet047 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp9 ibase#2fnet047 mq VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp8 mq mq_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp7 qf ckbb ibase#2fnet045 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp6 qf_x qf VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp4 mq_x ckbb ibase#2fnet027 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp3 qf ckb mq VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp1 ibase#2fnet027 D VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi3#2fp1 QN qf VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmi2#2fp1 Q qf_x VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_FDP_V2LP_2




.subckt SAEDRVT14_FILL16 VDD VSS VBP VBN
.ends SAEDRVT14_FILL16




.subckt SAEDRVT14_FILL2 VDD VSS VBP VBN
.ends SAEDRVT14_FILL2




.subckt SAEDRVT14_FILL32 VDD VSS VBP VBN
.ends SAEDRVT14_FILL32




.subckt SAEDRVT14_FILL3 VDD VSS VBP VBN
.ends SAEDRVT14_FILL3




.subckt SAEDRVT14_FILL4 VDD VSS VBP VBN
.ends SAEDRVT14_FILL4




.subckt SAEDRVT14_FILL5 VDD VSS VBP VBN
.ends SAEDRVT14_FILL5




.subckt SAEDRVT14_FILL64 VDD VSS VBP VBN
.ends SAEDRVT14_FILL64




.subckt SAEDRVT14_FILL8 VDD VSS VBP VBN
.ends SAEDRVT14_FILL8




.subckt SAEDRVT14_FILL_ECO_12 VDD VSS VBP VBN
Mxmmn1 net3 net3 net3 VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmmp1 net3 net3 net3 VBN n08 l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_FILL_ECO_12




.subckt SAEDRVT14_FILL_ECO_15 VDD VSS VBP VBN
Mxmmn1 net3 net3 net3 VBP p08 l=0.014u nf=5 m=1 nfin=4
Mxmmp1 net3 net3 net3 VBN n08 l=0.014u nf=5 m=1 nfin=4
.ends SAEDRVT14_FILL_ECO_15




.subckt SAEDRVT14_FILL_ECO_18 VDD VSS VBP VBN
Mxmmn1 net3 net3 net3 VBP p08 l=0.014u nf=6 m=1 nfin=4
Mxmmp1 net3 net3 net3 VBN n08 l=0.014u nf=6 m=1 nfin=4
.ends SAEDRVT14_FILL_ECO_18




.subckt SAEDRVT14_FILL_ECO_1 VDD VSS VBP VBN
.ends SAEDRVT14_FILL_ECO_1




.subckt SAEDRVT14_FILL_ECO_2 VDD VSS VBP VBN
.ends SAEDRVT14_FILL_ECO_2




.subckt SAEDRVT14_FILL_ECO_3 VDD VSS VBP VBN
Mxmmn1 net3 net3 net3 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp1 net3 net3 net3 VBN n08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FILL_ECO_3




.subckt SAEDRVT14_FILL_ECO_6 VDD VSS VBP VBN
Mxmmp1 net3 net3 net3 VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmmn1 net3 net3 net3 VBP p08 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_FILL_ECO_6




.subckt SAEDRVT14_FILL_ECO_9 VDD VSS VBP VBN
Mxmmp1 net3 net3 net3 VBN n08 l=0.014u nf=3 m=1 nfin=4
Mxmmn1 net3 net3 net3 VBP p08 l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_FILL_ECO_9




.subckt SAEDRVT14_FILL_NNWIV1Y2_2 VDD VSS VDDI
.ends SAEDRVT14_FILL_NNWIV1Y2_2




.subckt SAEDRVT14_FILL_NNWIV1Y2_3 VDD VSS VDDI
.ends SAEDRVT14_FILL_NNWIV1Y2_3




.subckt SAEDRVT14_FILL_NNWIY2_2 VDD VSS VDDI
.ends SAEDRVT14_FILL_NNWIY2_2




.subckt SAEDRVT14_FILL_NNWIY2_3 VDD VSS VDDI
.ends SAEDRVT14_FILL_NNWIY2_3




.subckt SAEDRVT14_FILL_NNWSPACERY2_7 VDD VSS VBP VBN
.ends SAEDRVT14_FILL_NNWSPACERY2_7




.subckt SAEDRVT14_FILL_NNWVDDBRKY2_3 VSS
.ends SAEDRVT14_FILL_NNWVDDBRKY2_3




.subckt SAEDRVT14_FILLP2 VDD VSS VDDR
.ends SAEDRVT14_FILLP2




.subckt SAEDRVT14_FILLP3 VDD VSS VDDR
.ends SAEDRVT14_FILLP3




.subckt SAEDRVT14_FILL_SPACER_7 VDD VSS
.ends SAEDRVT14_FILL_SPACER_7




.subckt SAEDRVT14_FILL_Y2_3 VDD VSS
.ends SAEDRVT14_FILL_Y2_3




.subckt SAEDRVT14_FSB2BDPRBQ_PV2_1 VDD VSS VDDR Q CK D SI SE RD B1 B2B
Mxn23 net035 mq net080 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn17 seb SE VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn10 net048 B2B net075 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn9 net079 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn8 mq ckbb qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn7 mq mq_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn6 net075 qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn4 net035 ckbb mq_x VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn3 net080 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn2 qf_x qf net079 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn1 ckbb ckb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn0 ckb CK VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn30 save_q B1 qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn29 save_qb save_q VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn28 save_q saveb net073 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn27 net073 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn26 net048 nrestoreb net077 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn25 net077 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn24 qf ckb net048 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn23 nrestoreb B2B VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn22 saveb B1 VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn5 mq_x ckb net025 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn4 net025 seb net029 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn3 net029 D VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn2 net025 SE net032 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn1 net032 SI VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn0 Q qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxp26 net035 ckb mq_x VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp25 net035 mq VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp24 net035 RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp15 seb SE VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp7 net048 nrestoreb net076 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp6 qf_x qf VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp5 net076 qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp4 qf ckb mq VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp2 mq_x ckbb net024 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp1 ckbb ckb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp0 ckb CK VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp30 save_q saveb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp29 save_qb save_q VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp28 net074 save_qb VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp27 save_q B1 net074 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp26 net078 save_qb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp25 net048 B2B net078 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp24 net048 ckbb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp23 nrestoreb B2B VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp22 saveb B1 VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp6 qf_x RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp5 mq mq_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp4 net024 SE net030 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp3 net030 D VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp2 net024 seb net031 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp1 net031 SI VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp0 Q qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FSB2BDPRBQ_PV2_1

.subckt SAEDRVT14_FSB2BDPRBQ4_PV2_1 VDD VSS VDDR Q0 Q1 Q2 Q3 CK D0 D1 D2 D3 SI SE RD B1 B2B
XI15 VDD VSS VDDR Q3 CK D3 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_1
XI14 VDD VSS VDDR Q2 CK D2 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_1
XI13 VDD VSS VDDR Q1 CK D1 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_1
XI12 VDD VSS VDDR Q0 CK D0 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_1
.ends SAEDRVT14_FSB2BDPRBQ4_PV2_1




.subckt SAEDRVT14_FSB2BDPRBQ_PV2_2 VDD VSS VDDR Q CK D SI SE RD B1 B2B
Mxn23 net035 mq net080 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn17 seb SE VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn10 net048 B2B net075 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn9 net079 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn8 mq ckbb qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn7 mq mq_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn6 net075 qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn4 net035 ckbb mq_x VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn3 net080 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn2 qf_x qf net079 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn1 ckbb ckb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn0 ckb CK VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn30 save_q B1 qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn29 save_qb save_q VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn28 save_q saveb net073 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn27 net073 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn26 net048 nrestoreb net077 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn25 net077 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn24 qf ckb net048 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn23 nrestoreb B2B VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn22 saveb B1 VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn5 mq_x ckb net025 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn4 net025 seb net029 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn3 net029 D VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn2 net025 SE net032 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn1 net032 SI VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn0 Q qf_x VSS VSS n08_hvt l=0.014u nf=2 m=1 nfin=4
Mxp26 net035 ckb mq_x VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp25 net035 mq VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp24 net035 RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp15 seb SE VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp7 net048 nrestoreb net076 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp6 qf_x qf VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp5 net076 qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp4 qf ckb mq VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp2 mq_x ckbb net024 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp1 ckbb ckb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp0 ckb CK VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp30 save_q saveb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp29 save_qb save_q VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp28 net074 save_qb VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp27 save_q B1 net074 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp26 net078 save_qb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp25 net048 B2B net078 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp24 net048 ckbb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp23 nrestoreb B2B VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp22 saveb B1 VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp6 qf_x RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp5 mq mq_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp4 net024 SE net030 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp3 net030 D VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp2 net024 seb net031 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp1 net031 SI VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp0 Q qf_x VDD VDDR p08_hvt l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_FSB2BDPRBQ_PV2_2

.subckt SAEDRVT14_FSB2BDPRBQ4_PV2_2 VDD VSS VDDR Q0 Q1 Q2 Q3 CK D0 D1 D2 D3 SI SE RD B1 B2B
XI11 VDD VSS VDDR Q3 CK D3 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_2
XI10 VDD VSS VDDR Q2 CK D2 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_2
XI9 VDD VSS VDDR Q1 CK D1 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_2
XI8 VDD VSS VDDR Q0 CK D0 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_2
.ends SAEDRVT14_FSB2BDPRBQ4_PV2_2




.subckt SAEDRVT14_FSB2BDPRBQ_PV2_4 VDD VSS VDDR Q CK D SI SE RD B1 B2B
Mxn23 net035 mq net080 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn17 seb SE VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn10 net048 B2B net075 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn9 net079 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn8 mq ckbb qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn7 mq mq_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn6 net075 qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn4 net035 ckbb mq_x VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn3 net080 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn2 qf_x qf net079 VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn1 ckbb ckb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn0 ckb CK VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn30 save_q B1 qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn29 save_qb save_q VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn28 save_q saveb net073 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn27 net073 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn26 net048 nrestoreb net077 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn25 net077 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn24 qf ckb net048 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn23 nrestoreb B2B VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn22 saveb B1 VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn5 mq_x ckb net025 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn4 net025 seb net029 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn3 net029 D VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn2 net025 SE net032 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn1 net032 SI VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn0 Q qf_x VSS VSS n08_hvt l=0.014u nf=4 m=1 nfin=4
Mxp26 net035 ckb mq_x VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp25 net035 mq VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp24 net035 RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp15 seb SE VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp7 net048 nrestoreb net076 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp6 qf_x qf VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=4
Mxp5 net076 qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp4 qf ckb mq VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp2 mq_x ckbb net024 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp1 ckbb ckb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp0 ckb CK VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp30 save_q saveb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp29 save_qb save_q VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp28 net074 save_qb VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp27 save_q B1 net074 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp26 net078 save_qb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp25 net048 B2B net078 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp24 net048 ckbb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp23 nrestoreb B2B VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp22 saveb B1 VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp6 qf_x RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=4
Mxmp5 mq mq_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp4 net024 SE net030 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp3 net030 D VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp2 net024 seb net031 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp1 net031 SI VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp0 Q qf_x VDD VDDR p08_hvt l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_FSB2BDPRBQ_PV2_4

.subckt SAEDRVT14_FSB2BDPRBQ4_PV2_4 VDD VSS VDDR Q0 Q1 Q2 Q3 CK D0 D1 D2 D3 SI SE RD B1 B2B
XI12 VDD VSS VDDR Q0 CK D0 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_4
XI11 VDD VSS VDDR Q3 CK D3 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_4
XI10 VDD VSS VDDR Q2 CK D2 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_4
XI9 VDD VSS VDDR Q1 CK D1 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_4
.ends SAEDRVT14_FSB2BDPRBQ4_PV2_4




.subckt SAEDRVT14_FSB2BDPRBQ_PV2_8 VDD VSS VDDR Q CK D SI SE RD B1 B2B
Mxn91 net0791 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn23 net035 mq net080 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn21 qf_x qf net0791 VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn17 seb SE VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn10 net048 B2B net075 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn9 net079 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn8 mq ckbb qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn7 mq mq_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn6 net075 qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn4 net035 ckbb mq_x VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn3 net080 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn2 qf_x qf net079 VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn1 ckbb ckb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn0 ckb CK VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn30 save_q B1 qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn29 save_qb save_q VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn28 save_q saveb net073 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn27 net073 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn26 net048 nrestoreb net077 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn25 net077 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn24 qf ckb net048 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn23 nrestoreb B2B VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn22 saveb B1 VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn5 mq_x ckb net025 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn4 net025 seb net029 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn3 net029 D VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn2 net025 SE net032 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn1 net032 SI VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn0 Q qf_x VSS VSS n08_hvt l=0.014u nf=8 m=1 nfin=4
Mxp26 net035 ckb mq_x VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp25 net035 mq VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp24 net035 RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp15 seb SE VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp7 net048 nrestoreb net076 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp6 qf_x qf VDD VDDR p08_hvt l=0.014u nf=2 m=1 nfin=4
Mxp5 net076 qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp4 qf ckb mq VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp2 mq_x ckbb net024 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp1 ckbb ckb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp0 ckb CK VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp30 save_q saveb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp29 save_qb save_q VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp28 net074 save_qb VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp27 save_q B1 net074 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp26 net078 save_qb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp25 net048 B2B net078 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp24 net048 ckbb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp23 nrestoreb B2B VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp22 saveb B1 VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp6 qf_x RD VDD VDDR p08_hvt l=0.014u nf=2 m=1 nfin=4
Mxmp5 mq mq_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp4 net024 SE net030 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp3 net030 D VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp2 net024 seb net031 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp1 net031 SI VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp0 Q qf_x VDD VDDR p08_hvt l=0.014u nf=8 m=1 nfin=4
.ends SAEDRVT14_FSB2BDPRBQ_PV2_8

.subckt SAEDRVT14_FSB2BDPRBQ4_PV2_8 VDD VSS VDDR Q0 Q1 Q2 Q3 CK D0 D1 D2 D3 SI SE RD B1 B2B
XI8 VDD VSS VDDR Q0 CK D0 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_8
XI9 VDD VSS VDDR Q1 CK D1 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_8
XI10 VDD VSS VDDR Q2 CK D2 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_8
XI11 VDD VSS VDDR Q3 CK D3 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_8
.ends SAEDRVT14_FSB2BDPRBQ4_PV2_8




.subckt SAEDRVT14_FSB2BDPRBQ_PV2_1 VDD VSS VDDR Q CK D SI SE RD B1 B2B
Mxn23 net035 mq net080 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn17 seb SE VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn10 net048 B2B net075 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn9 net079 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn8 mq ckbb qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn7 mq mq_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn6 net075 qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn4 net035 ckbb mq_x VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn3 net080 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn2 qf_x qf net079 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn1 ckbb ckb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn0 ckb CK VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn30 save_q B1 qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn29 save_qb save_q VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn28 save_q saveb net073 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn27 net073 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn26 net048 nrestoreb net077 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn25 net077 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn24 qf ckb net048 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn23 nrestoreb B2B VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn22 saveb B1 VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn5 mq_x ckb net025 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn4 net025 seb net029 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn3 net029 D VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn2 net025 SE net032 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn1 net032 SI VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn0 Q qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxp26 net035 ckb mq_x VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp25 net035 mq VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp24 net035 RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp15 seb SE VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp7 net048 nrestoreb net076 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp6 qf_x qf VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp5 net076 qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp4 qf ckb mq VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp2 mq_x ckbb net024 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp1 ckbb ckb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp0 ckb CK VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp30 save_q saveb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp29 save_qb save_q VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp28 net074 save_qb VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp27 save_q B1 net074 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp26 net078 save_qb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp25 net048 B2B net078 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp24 net048 ckbb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp23 nrestoreb B2B VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp22 saveb B1 VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp6 qf_x RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp5 mq mq_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp4 net024 SE net030 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp3 net030 D VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp2 net024 seb net031 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp1 net031 SI VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp0 Q qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FSB2BDPRBQ_PV2_1

.subckt SAEDRVT14_FSB2BDPRBQ8_PV2_1 VDD VSS VDDR Q0 Q1 Q2 Q3 CK D0 D1 D2 D3 SI SE RD B1 B2B D4 D5 D6 D7 Q4 Q5 Q6 Q7
XI31 VDD VSS VDDR Q3 CK D3 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_1
XI24 VDD VSS VDDR Q7 CK D7 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_1
XI25 VDD VSS VDDR Q5 CK D5 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_1
XI26 VDD VSS VDDR Q4 CK D4 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_1
XI29 VDD VSS VDDR Q1 CK D1 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_1
XI27 VDD VSS VDDR Q6 CK D6 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_1
XI28 VDD VSS VDDR Q0 CK D0 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_1
XI30 VDD VSS VDDR Q2 CK D2 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_1
.ends SAEDRVT14_FSB2BDPRBQ8_PV2_1




.subckt SAEDRVT14_FSB2BDPRBQ_PV2_2 VDD VSS VDDR Q CK D SI SE RD B1 B2B
Mxn23 net035 mq net080 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn17 seb SE VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn10 net048 B2B net075 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn9 net079 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn8 mq ckbb qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn7 mq mq_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn6 net075 qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn4 net035 ckbb mq_x VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn3 net080 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn2 qf_x qf net079 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn1 ckbb ckb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn0 ckb CK VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn30 save_q B1 qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn29 save_qb save_q VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn28 save_q saveb net073 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn27 net073 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn26 net048 nrestoreb net077 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn25 net077 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn24 qf ckb net048 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn23 nrestoreb B2B VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn22 saveb B1 VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn5 mq_x ckb net025 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn4 net025 seb net029 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn3 net029 D VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn2 net025 SE net032 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn1 net032 SI VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn0 Q qf_x VSS VSS n08_hvt l=0.014u nf=2 m=1 nfin=4
Mxp26 net035 ckb mq_x VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp25 net035 mq VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp24 net035 RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp15 seb SE VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp7 net048 nrestoreb net076 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp6 qf_x qf VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp5 net076 qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp4 qf ckb mq VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp2 mq_x ckbb net024 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp1 ckbb ckb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp0 ckb CK VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp30 save_q saveb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp29 save_qb save_q VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp28 net074 save_qb VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp27 save_q B1 net074 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp26 net078 save_qb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp25 net048 B2B net078 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp24 net048 ckbb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp23 nrestoreb B2B VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp22 saveb B1 VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp6 qf_x RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp5 mq mq_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp4 net024 SE net030 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp3 net030 D VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp2 net024 seb net031 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp1 net031 SI VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp0 Q qf_x VDD VDDR p08_hvt l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_FSB2BDPRBQ_PV2_2

.subckt SAEDRVT14_FSB2BDPRBQ8_PV2_2 VDD VSS VDDR Q0 Q1 Q2 Q3 CK D0 D1 D2 D3 SI SE RD B1 B2B D4 D5 D6 D7 Q4 Q5 Q6 Q7
XI19 VDD VSS VDDR Q3 CK D3 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_2
XI18 VDD VSS VDDR Q2 CK D2 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_2
XI17 VDD VSS VDDR Q1 CK D1 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_2
XI16 VDD VSS VDDR Q0 CK D0 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_2
XI13 VDD VSS VDDR Q5 CK D5 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_2
XI15 VDD VSS VDDR Q6 CK D6 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_2
XI14 VDD VSS VDDR Q4 CK D4 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_2
XI12 VDD VSS VDDR Q7 CK D7 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_2
.ends SAEDRVT14_FSB2BDPRBQ8_PV2_2




.subckt SAEDRVT14_FSB2BDPRBQ_PV2_4 VDD VSS VDDR Q CK D SI SE RD B1 B2B
Mxn23 net035 mq net080 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn17 seb SE VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn10 net048 B2B net075 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn9 net079 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn8 mq ckbb qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn7 mq mq_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn6 net075 qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn4 net035 ckbb mq_x VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn3 net080 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn2 qf_x qf net079 VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn1 ckbb ckb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn0 ckb CK VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn30 save_q B1 qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn29 save_qb save_q VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn28 save_q saveb net073 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn27 net073 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn26 net048 nrestoreb net077 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn25 net077 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn24 qf ckb net048 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn23 nrestoreb B2B VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn22 saveb B1 VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn5 mq_x ckb net025 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn4 net025 seb net029 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn3 net029 D VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn2 net025 SE net032 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn1 net032 SI VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn0 Q qf_x VSS VSS n08_hvt l=0.014u nf=4 m=1 nfin=4
Mxp26 net035 ckb mq_x VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp25 net035 mq VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp24 net035 RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp15 seb SE VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp7 net048 nrestoreb net076 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp6 qf_x qf VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=4
Mxp5 net076 qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp4 qf ckb mq VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp2 mq_x ckbb net024 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp1 ckbb ckb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp0 ckb CK VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp30 save_q saveb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp29 save_qb save_q VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp28 net074 save_qb VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp27 save_q B1 net074 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp26 net078 save_qb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp25 net048 B2B net078 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp24 net048 ckbb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp23 nrestoreb B2B VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp22 saveb B1 VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp6 qf_x RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=4
Mxmp5 mq mq_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp4 net024 SE net030 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp3 net030 D VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp2 net024 seb net031 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp1 net031 SI VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp0 Q qf_x VDD VDDR p08_hvt l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_FSB2BDPRBQ_PV2_4

.subckt SAEDRVT14_FSB2BDPRBQ8_PV2_4 VDD VSS VDDR Q0 Q1 Q2 Q3 CK D0 D1 D2 D3 SI SE RD B1 B2B D4 D5 D6 D7 Q4 Q5 Q6 Q7
XI19 VDD VSS VDDR Q3 CK D3 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_4
XI18 VDD VSS VDDR Q2 CK D2 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_4
XI17 VDD VSS VDDR Q1 CK D1 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_4
XI16 VDD VSS VDDR Q0 CK D0 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_4
XI13 VDD VSS VDDR Q5 CK D5 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_4
XI15 VDD VSS VDDR Q6 CK D6 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_4
XI14 VDD VSS VDDR Q4 CK D4 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_4
XI12 VDD VSS VDDR Q7 CK D7 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_4
.ends SAEDRVT14_FSB2BDPRBQ8_PV2_4




.subckt SAEDRVT14_FSB2BDPRBQ_PV2_8 VDD VSS VDDR Q CK D SI SE RD B1 B2B
Mxn91 net0791 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn23 net035 mq net080 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn21 qf_x qf net0791 VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn17 seb SE VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn10 net048 B2B net075 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn9 net079 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn8 mq ckbb qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn7 mq mq_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn6 net075 qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn4 net035 ckbb mq_x VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn3 net080 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn2 qf_x qf net079 VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn1 ckbb ckb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn0 ckb CK VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn30 save_q B1 qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn29 save_qb save_q VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn28 save_q saveb net073 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn27 net073 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn26 net048 nrestoreb net077 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn25 net077 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn24 qf ckb net048 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn23 nrestoreb B2B VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn22 saveb B1 VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn5 mq_x ckb net025 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn4 net025 seb net029 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn3 net029 D VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn2 net025 SE net032 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn1 net032 SI VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn0 Q qf_x VSS VSS n08_hvt l=0.014u nf=8 m=1 nfin=4
Mxp26 net035 ckb mq_x VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp25 net035 mq VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp24 net035 RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp15 seb SE VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp7 net048 nrestoreb net076 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp6 qf_x qf VDD VDDR p08_hvt l=0.014u nf=2 m=1 nfin=4
Mxp5 net076 qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp4 qf ckb mq VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp2 mq_x ckbb net024 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp1 ckbb ckb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp0 ckb CK VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp30 save_q saveb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp29 save_qb save_q VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp28 net074 save_qb VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp27 save_q B1 net074 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp26 net078 save_qb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp25 net048 B2B net078 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp24 net048 ckbb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp23 nrestoreb B2B VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp22 saveb B1 VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp6 qf_x RD VDD VDDR p08_hvt l=0.014u nf=2 m=1 nfin=4
Mxmp5 mq mq_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp4 net024 SE net030 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp3 net030 D VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp2 net024 seb net031 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp1 net031 SI VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp0 Q qf_x VDD VDDR p08_hvt l=0.014u nf=8 m=1 nfin=4
.ends SAEDRVT14_FSB2BDPRBQ_PV2_8

.subckt SAEDRVT14_FSB2BDPRBQ8_PV2_8 VDD VSS VDDR Q0 Q1 Q2 Q3 CK D0 D1 D2 D3 SI SE RD B1 B2B D4 D5 D6 D7 Q4 Q5 Q6 Q7
XI20 VDD VSS VDDR Q3 CK D3 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_8
XI19 VDD VSS VDDR Q2 CK D2 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_8
XI18 VDD VSS VDDR Q1 CK D1 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_8
XI17 VDD VSS VDDR Q0 CK D0 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_8
XI14 VDD VSS VDDR Q5 CK D5 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_8
XI16 VDD VSS VDDR Q6 CK D6 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_8
XI15 VDD VSS VDDR Q4 CK D4 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_8
XI13 VDD VSS VDDR Q7 CK D7 SI SE RD B1 B2B SAEDRVT14_FSB2BDPRBQ_PV2_8
.ends SAEDRVT14_FSB2BDPRBQ8_PV2_8




.subckt SAEDRVT14_FSB2BDPRBQ_PV2_1 VDD VSS VDDR Q CK D SI SE RD B1 B2B
Mxn23 net035 mq net080 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn17 seb SE VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn10 net048 B2B net075 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn9 net079 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn8 mq ckbb qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn7 mq mq_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn6 net075 qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn4 net035 ckbb mq_x VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn3 net080 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn2 qf_x qf net079 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn1 ckbb ckb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn0 ckb CK VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn30 save_q B1 qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn29 save_qb save_q VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn28 save_q saveb net073 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn27 net073 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn26 net048 nrestoreb net077 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn25 net077 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn24 qf ckb net048 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn23 nrestoreb B2B VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn22 saveb B1 VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn5 mq_x ckb net025 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn4 net025 seb net029 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn3 net029 D VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn2 net025 SE net032 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn1 net032 SI VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn0 Q qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxp26 net035 ckb mq_x VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp25 net035 mq VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp24 net035 RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp15 seb SE VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp7 net048 nrestoreb net076 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp6 qf_x qf VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp5 net076 qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp4 qf ckb mq VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp2 mq_x ckbb net024 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp1 ckbb ckb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp0 ckb CK VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp30 save_q saveb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp29 save_qb save_q VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp28 net074 save_qb VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp27 save_q B1 net074 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp26 net078 save_qb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp25 net048 B2B net078 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp24 net048 ckbb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp23 nrestoreb B2B VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp22 saveb B1 VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp6 qf_x RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp5 mq mq_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp4 net024 SE net030 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp3 net030 D VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp2 net024 seb net031 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp1 net031 SI VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp0 Q qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FSB2BDPRBQ_PV2_1




.subckt SAEDRVT14_FSB2BDPRBQ_PV2_2 VDD VSS VDDR Q CK D SI SE RD B1 B2B
Mxn23 net035 mq net080 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn17 seb SE VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn10 net048 B2B net075 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn9 net079 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn8 mq ckbb qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn7 mq mq_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn6 net075 qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn4 net035 ckbb mq_x VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn3 net080 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn2 qf_x qf net079 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn1 ckbb ckb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn0 ckb CK VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn30 save_q B1 qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn29 save_qb save_q VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn28 save_q saveb net073 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn27 net073 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn26 net048 nrestoreb net077 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn25 net077 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn24 qf ckb net048 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn23 nrestoreb B2B VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn22 saveb B1 VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn5 mq_x ckb net025 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn4 net025 seb net029 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn3 net029 D VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn2 net025 SE net032 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn1 net032 SI VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn0 Q qf_x VSS VSS n08_hvt l=0.014u nf=2 m=1 nfin=4
Mxp26 net035 ckb mq_x VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp25 net035 mq VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp24 net035 RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp15 seb SE VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp7 net048 nrestoreb net076 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp6 qf_x qf VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp5 net076 qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp4 qf ckb mq VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp2 mq_x ckbb net024 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp1 ckbb ckb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp0 ckb CK VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp30 save_q saveb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp29 save_qb save_q VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp28 net074 save_qb VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp27 save_q B1 net074 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp26 net078 save_qb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp25 net048 B2B net078 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp24 net048 ckbb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp23 nrestoreb B2B VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp22 saveb B1 VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp6 qf_x RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp5 mq mq_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp4 net024 SE net030 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp3 net030 D VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp2 net024 seb net031 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp1 net031 SI VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp0 Q qf_x VDD VDDR p08_hvt l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_FSB2BDPRBQ_PV2_2




.subckt SAEDRVT14_FSB2BDPRBQ_PV2_4 VDD VSS VDDR Q CK D SI SE RD B1 B2B
Mxn23 net035 mq net080 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn17 seb SE VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn10 net048 B2B net075 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn9 net079 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn8 mq ckbb qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn7 mq mq_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn6 net075 qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn4 net035 ckbb mq_x VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn3 net080 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn2 qf_x qf net079 VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn1 ckbb ckb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn0 ckb CK VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn30 save_q B1 qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn29 save_qb save_q VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn28 save_q saveb net073 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn27 net073 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn26 net048 nrestoreb net077 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn25 net077 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn24 qf ckb net048 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn23 nrestoreb B2B VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn22 saveb B1 VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn5 mq_x ckb net025 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn4 net025 seb net029 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn3 net029 D VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn2 net025 SE net032 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn1 net032 SI VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn0 Q qf_x VSS VSS n08_hvt l=0.014u nf=4 m=1 nfin=4
Mxp26 net035 ckb mq_x VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp25 net035 mq VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp24 net035 RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp15 seb SE VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp7 net048 nrestoreb net076 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp6 qf_x qf VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=4
Mxp5 net076 qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp4 qf ckb mq VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp2 mq_x ckbb net024 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp1 ckbb ckb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp0 ckb CK VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp30 save_q saveb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp29 save_qb save_q VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp28 net074 save_qb VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp27 save_q B1 net074 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp26 net078 save_qb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp25 net048 B2B net078 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp24 net048 ckbb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp23 nrestoreb B2B VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp22 saveb B1 VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp6 qf_x RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=4
Mxmp5 mq mq_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp4 net024 SE net030 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp3 net030 D VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp2 net024 seb net031 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp1 net031 SI VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp0 Q qf_x VDD VDDR p08_hvt l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_FSB2BDPRBQ_PV2_4




.subckt SAEDRVT14_FSB2BDPRBQ_PV2_8 VDD VSS VDDR Q CK D SI SE RD B1 B2B
Mxn91 net0791 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn23 net035 mq net080 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn21 qf_x qf net0791 VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn17 seb SE VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn10 net048 B2B net075 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn9 net079 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn8 mq ckbb qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn7 mq mq_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn6 net075 qf_x VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn4 net035 ckbb mq_x VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn3 net080 RD VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn2 qf_x qf net079 VSS n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxn1 ckbb ckb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxn0 ckb CK VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn30 save_q B1 qf VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn29 save_qb save_q VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn28 save_q saveb net073 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn27 net073 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn26 net048 nrestoreb net077 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn25 net077 save_qb VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn24 qf ckb net048 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn23 nrestoreb B2B VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn22 saveb B1 VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn5 mq_x ckb net025 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn4 net025 seb net029 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn3 net029 D VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn2 net025 SE net032 VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn1 net032 SI VSS VSS n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmn0 Q qf_x VSS VSS n08_hvt l=0.014u nf=8 m=1 nfin=4
Mxp26 net035 ckb mq_x VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp25 net035 mq VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp24 net035 RD VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp15 seb SE VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp7 net048 nrestoreb net076 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp6 qf_x qf VDD VDDR p08_hvt l=0.014u nf=2 m=1 nfin=4
Mxp5 net076 qf_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp4 qf ckb mq VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp2 mq_x ckbb net024 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp1 ckbb ckb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxp0 ckb CK VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp30 save_q saveb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp29 save_qb save_q VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp28 net074 save_qb VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp27 save_q B1 net074 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp26 net078 save_qb VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp25 net048 B2B net078 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp24 net048 ckbb qf VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp23 nrestoreb B2B VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp22 saveb B1 VDDR VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp6 qf_x RD VDD VDDR p08_hvt l=0.014u nf=2 m=1 nfin=4
Mxmp5 mq mq_x VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp4 net024 SE net030 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp3 net030 D VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp2 net024 seb net031 VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp1 net031 SI VDD VDDR p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmp0 Q qf_x VDD VDDR p08_hvt l=0.014u nf=8 m=1 nfin=4
.ends SAEDRVT14_FSB2BDPRBQ_PV2_8




.subckt SAEDRVT14_FSDN_V2_0P5 VDD VSS VBP VBN Q QN CK D SI SE
Mxmn1 ckbb ckb VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmn0 ckb CK VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn13 ibase#2fnet046 qf_x VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn12 mq_x ckb ibase#2fnet048 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn11 ibase#2fnet048 mq VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn10 mq mq_x VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn9 qf ckbb ibase#2fnet046 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn8 qf_x qf VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn6 mq_x ckbb net14 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn5 mq ckb qf VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi3#2fn0 Q qf_x VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmi2#2fn0 QN qf VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fn17 i0#2fseb SE VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn3 net14 D i0#2fnet22 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn2 i0#2fnet22 i0#2fseb VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn1 net14 SE i0#2fnet19 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn0 i0#2fnet19 SI VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmp1 ckbb ckb VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmp0 ckb CK VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp11 ibase#2fnet045 qf_x VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp10 mq_x ckbb ibase#2fnet047 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp9 ibase#2fnet047 mq VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp8 mq mq_x VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp7 qf ckb ibase#2fnet045 VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp6 qf_x qf VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp4 mq_x ckb net25 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp3 qf ckbb mq VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmi3#2fp1 Q qf_x VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmi2#2fp1 QN qf VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fp15 i0#2fseb SE VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp3 net25 D i0#2fnet21 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp2 i0#2fnet21 SE VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp1 net25 i0#2fseb i0#2fnet20 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp0 i0#2fnet20 SI VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_0P5

.subckt SAEDRVT14_FSDN2_V2_0P5 VDD VSS VBP VBN Q0 Q1 QN0 QN1 CK D0 D1 SI SE
XI9 VDD VSS VBP VBN Q0 QN0 CK D0 SI SE SAEDRVT14_FSDN_V2_0P5
XI10 VDD VSS VBP VBN Q1 QN1 CK D1 SI SE SAEDRVT14_FSDN_V2_0P5
.ends SAEDRVT14_FSDN2_V2_0P5




.subckt SAEDRVT14_FSDN_V2_1 VDD VSS VBP VBN Q QN CK D SI SE
Mxmn1 ckbb ckb VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmn0 ckb CK VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn13 ibase#2fnet046 qf_x VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn12 mq_x ckb ibase#2fnet048 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn11 ibase#2fnet048 mq VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn10 mq mq_x VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn9 qf ckbb ibase#2fnet046 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn8 qf_x qf VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn6 mq_x ckbb net14 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn5 mq ckb qf VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi3#2fn0 Q qf_x VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxmi2#2fn0 QN qf VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn17 i0#2fseb SE VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn3 net14 D i0#2fnet22 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn2 i0#2fnet22 i0#2fseb VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn1 net14 SE i0#2fnet19 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn0 i0#2fnet19 SI VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmp1 ckbb ckb VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmp0 ckb CK VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp11 ibase#2fnet045 qf_x VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp10 mq_x ckbb ibase#2fnet047 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp9 ibase#2fnet047 mq VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp8 mq mq_x VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp7 qf ckb ibase#2fnet045 VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp6 qf_x qf VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp4 mq_x ckb net25 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp3 qf ckbb mq VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmi3#2fp1 Q qf_x VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=4
Mxmi2#2fp1 QN qf VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp15 i0#2fseb SE VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp3 net25 D i0#2fnet21 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp2 i0#2fnet21 SE VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp1 net25 i0#2fseb i0#2fnet20 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp0 i0#2fnet20 SI VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_1

.subckt SAEDRVT14_FSDN2_V2_1 VDD VSS VBP VBN Q0 Q1 QN0 QN1 CK D0 D1 SI SE
XI2 VDD VSS VBP VBN Q0 QN0 CK D0 SI SE SAEDRVT14_FSDN_V2_1
XI3 VDD VSS VBP VBN Q1 QN1 CK D1 SI SE SAEDRVT14_FSDN_V2_1
.ends SAEDRVT14_FSDN2_V2_1




.subckt SAEDRVT14_FSDN_V2_2 VDD VSS VBP VBN Q QN CK D SI SE
Mxmn1 ckbb ckb VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmn0 ckb CK VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn13 ibase#2fnet046 qf_x VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn12 mq_x ckb ibase#2fnet048 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn11 ibase#2fnet048 mq VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn10 mq mq_x VSS VBN n08_hvt l=0.014u nf=2 m=1 nfin=3
Mxmibase#2fn9 qf ckbb ibase#2fnet046 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn8 qf_x qf VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn6 mq_x ckbb net017 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn5 mq ckb qf VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi3#2fn0 Q qf_x VSS VBN n08_hvt l=0.014u nf=2 m=1 nfin=4
Mxmi2#2fn0 QN qf VSS VBN n08_hvt l=0.014u nf=2 m=1 nfin=4
Mxmi0#2fn17 i0#2fseb SE VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn3 net017 D i0#2fnet22 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn2 i0#2fnet22 i0#2fseb VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn1 net017 SE i0#2fnet19 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn0 i0#2fnet19 SI VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmp1 ckbb ckb VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmp0 ckb CK VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp11 ibase#2fnet045 qf_x VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp10 mq_x ckbb ibase#2fnet047 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp9 ibase#2fnet047 mq VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp8 mq mq_x VDD VBP p08_hvt l=0.014u nf=2 m=1 nfin=3
Mxmibase#2fp7 qf ckb ibase#2fnet045 VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp6 qf_x qf VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp4 mq_x ckb net019 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp3 qf ckbb mq VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmi3#2fp1 Q qf_x VDD VBP p08_hvt l=0.014u nf=2 m=1 nfin=4
Mxmi2#2fp1 QN qf VDD VBP p08_hvt l=0.014u nf=2 m=1 nfin=4
Mxmi0#2fp15 i0#2fseb SE VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp3 net019 D i0#2fnet21 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp2 i0#2fnet21 SE VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp1 net019 i0#2fseb i0#2fnet20 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp0 i0#2fnet20 SI VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_2

.subckt SAEDRVT14_FSDN2_V2_2 VDD VSS VBP VBN Q0 Q1 QN0 QN1 CK D0 D1 SI SE
XI0 VDD VSS VBP VBN Q0 QN0 CK D0 SI SE SAEDRVT14_FSDN_V2_2
XI1 VDD VSS VBP VBN Q1 QN1 CK D1 SI SE SAEDRVT14_FSDN_V2_2
.ends SAEDRVT14_FSDN2_V2_2




.subckt SAEDRVT14_FSDN_V2_4 VDD VSS VBP VBN Q QN CK D SI SE
Mxmp1 ckbb ckb VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 ckb CK VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp11 ibase#2fnet045 qf_x VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp10 mq_x ckbb ibase#2fnet047 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp9 ibase#2fnet047 mq VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp8 mq mq_x VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmibase#2fp7 qf ckb ibase#2fnet045 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp6 qf_x qf VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp4 mq_x ckb net019 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp3 qf ckbb mq VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmi3#2fp1 Q qf_x VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmi2#2fp1 QN qf VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmi0#2fp15 i0#2fseb SE VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp3 net019 D i0#2fnet21 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp2 i0#2fnet21 SE VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp1 net019 i0#2fseb i0#2fnet20 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp0 i0#2fnet20 SI VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmn1 ckbb ckb VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 ckb CK VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn13 ibase#2fnet046 qf_x VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn12 mq_x ckb ibase#2fnet048 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn11 ibase#2fnet048 mq VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn10 mq mq_x VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmibase#2fn9 qf ckbb ibase#2fnet046 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn8 qf_x qf VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn6 mq_x ckbb net017 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn5 mq ckb qf VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi3#2fn0 Q qf_x VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmi2#2fn0 QN qf VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmi0#2fn17 i0#2fseb SE VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn3 net017 D i0#2fnet22 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn2 i0#2fnet22 i0#2fseb VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn1 net017 SE i0#2fnet19 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn0 i0#2fnet19 SI VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_4

.subckt SAEDRVT14_FSDN2_V2_4 VDD VSS VBP VBN Q0 Q1 QN0 QN1 CK D0 D1 SI SE
XI2 VDD VSS VBP VBN Q0 QN0 CK D0 SI SE SAEDRVT14_FSDN_V2_4
XI3 VDD VSS VBP VBN Q1 QN1 CK D1 SI SE SAEDRVT14_FSDN_V2_4
.ends SAEDRVT14_FSDN2_V2_4




.subckt SAEDRVT14_FSDN_V2_0P5 VDD VSS VBP VBN Q QN CK D SI SE
Mxmn1 ckbb ckb VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmn0 ckb CK VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn13 ibase#2fnet046 qf_x VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn12 mq_x ckb ibase#2fnet048 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn11 ibase#2fnet048 mq VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn10 mq mq_x VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn9 qf ckbb ibase#2fnet046 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn8 qf_x qf VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn6 mq_x ckbb net14 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn5 mq ckb qf VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi3#2fn0 Q qf_x VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmi2#2fn0 QN qf VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fn17 i0#2fseb SE VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn3 net14 D i0#2fnet22 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn2 i0#2fnet22 i0#2fseb VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn1 net14 SE i0#2fnet19 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn0 i0#2fnet19 SI VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmp1 ckbb ckb VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmp0 ckb CK VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp11 ibase#2fnet045 qf_x VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp10 mq_x ckbb ibase#2fnet047 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp9 ibase#2fnet047 mq VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp8 mq mq_x VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp7 qf ckb ibase#2fnet045 VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp6 qf_x qf VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp4 mq_x ckb net25 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp3 qf ckbb mq VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmi3#2fp1 Q qf_x VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmi2#2fp1 QN qf VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmi0#2fp15 i0#2fseb SE VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp3 net25 D i0#2fnet21 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp2 i0#2fnet21 SE VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp1 net25 i0#2fseb i0#2fnet20 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp0 i0#2fnet20 SI VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_0P5

.subckt SAEDRVT14_FSDN4_V2_0P5 VDD VSS VBP VBN Q0 Q1 Q2 Q3 QN0 QN1 QN2 QN3 CK D0 D1 D2 D3 SI SE
XI1 VDD VSS VBP VBN Q1 QN1 CK D1 SI SE SAEDRVT14_FSDN_V2_0P5
XI0 VDD VSS VBP VBN Q0 QN0 CK D0 SI SE SAEDRVT14_FSDN_V2_0P5
XI2 VDD VSS VBP VBN Q2 QN2 CK D2 SI SE SAEDRVT14_FSDN_V2_0P5
XI3 VDD VSS VBP VBN Q3 QN3 CK D3 SI SE SAEDRVT14_FSDN_V2_0P5
.ends SAEDRVT14_FSDN4_V2_0P5




.subckt SAEDRVT14_FSDN_V2_1 VDD VSS VBP VBN Q QN CK D SI SE
Mxmn1 ckbb ckb VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmn0 ckb CK VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn13 ibase#2fnet046 qf_x VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn12 mq_x ckb ibase#2fnet048 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn11 ibase#2fnet048 mq VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn10 mq mq_x VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn9 qf ckbb ibase#2fnet046 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn8 qf_x qf VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fn6 mq_x ckbb net14 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fn5 mq ckb qf VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi3#2fn0 Q qf_x VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxmi2#2fn0 QN qf VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fn17 i0#2fseb SE VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn3 net14 D i0#2fnet22 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn2 i0#2fnet22 i0#2fseb VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn1 net14 SE i0#2fnet19 VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmn0 i0#2fnet19 SI VSS VBN n08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmp1 ckbb ckb VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmp0 ckb CK VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp11 ibase#2fnet045 qf_x VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp10 mq_x ckbb ibase#2fnet047 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp9 ibase#2fnet047 mq VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp8 mq mq_x VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp7 qf ckb ibase#2fnet045 VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp6 qf_x qf VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmibase#2fp4 mq_x ckb net25 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmibase#2fp3 qf ckbb mq VBP p08_hvt l=0.014u nf=1 m=1 nfin=2
Mxmi3#2fp1 Q qf_x VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=4
Mxmi2#2fp1 QN qf VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=4
Mxmi0#2fp15 i0#2fseb SE VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp3 net25 D i0#2fnet21 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp2 i0#2fnet21 SE VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp1 net25 i0#2fseb i0#2fnet20 VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
Mxmi0#2fmp0 i0#2fnet20 SI VDD VBP p08_hvt l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_1

.subckt SAEDRVT14_FSDN4_V2_1 VDD VSS VBP VBN Q0 Q1 Q2 Q3 QN0 QN1 QN2 QN3 CK D0 D1 D2 D3 SI SE
XI3 VDD VSS VBP VBN Q3 QN3 CK D3 SI SE SAEDRVT14_FSDN_V2_1
XI2 VDD VSS VBP VBN Q2 QN2 CK D2 SI SE SAEDRVT14_FSDN_V2_1
XI1 VDD VSS VBP VBN Q1 QN1 CK D1 SI SE SAEDRVT14_FSDN_V2_1
XI0 VDD VSS VBP VBN Q0 QN0 CK D0 SI SE SAEDRVT14_FSDN_V2_1
.ends SAEDRVT14_FSDN4_V2_1




.subckt SAEDRVT14_FSDN_V2_2 vdd vss vbp vbn q qn ck d si se
xmn1 ckbb ckb vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_hvt l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb net017 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 q qf_x vss vbn n08_hvt l=0.014u nf=2 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_hvt l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net017 d i0#2fnet22 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net017 se i0#2fnet19 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_hvt l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb net019 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_hvt l=0.014u nf=2 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_hvt l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net019 d i0#2fnet21 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net019 i0#2fseb i0#2fnet20 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_2

.subckt SAEDRVT14_FSDN4_V2_2 vdd vss vbp vbn q0 q1 q2 q3 qn0 qn1 qn2 qn3 ck d0 d1 d2 d3 si se
xi3 vdd vss vbp vbn q3 qn3 ck d3 si se SAEDRVT14_FSDN_V2_2
xi2 vdd vss vbp vbn q2 qn2 ck d2 si se SAEDRVT14_FSDN_V2_2
xi1 vdd vss vbp vbn q1 qn1 ck d1 si se SAEDRVT14_FSDN_V2_2
xi0 vdd vss vbp vbn q0 qn0 ck d0 si se SAEDRVT14_FSDN_V2_2
.ends SAEDRVT14_FSDN4_V2_2




.subckt SAEDRVT14_FSDN_V2_4 vdd vss vbp vbn q qn ck d si se
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb net019 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net019 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net019 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb net017 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net017 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net017 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_4

.subckt SAEDRVT14_FSDN4_V2_4 vdd vss vbp vbn q0 q1 q2 q3 qn0 qn1 qn2 qn3 ck d0 d1 d2 d3 si se
xi3 vdd vss vbp vbn q3 qn3 ck d3 si se SAEDRVT14_FSDN_V2_4
xi2 vdd vss vbp vbn q2 qn2 ck d2 si se SAEDRVT14_FSDN_V2_4
xi1 vdd vss vbp vbn q1 qn1 ck d1 si se SAEDRVT14_FSDN_V2_4
xi0 vdd vss vbp vbn q0 qn0 ck d0 si se SAEDRVT14_FSDN_V2_4
.ends SAEDRVT14_FSDN4_V2_4




.subckt SAEDRVT14_FSDN_V2_0P5 vdd vss vbp vbn q qn ck d si se
xmn1 ckbb ckb vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb net14 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 q qf_x vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 qn qf vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net14 d i0#2fnet22 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net14 se i0#2fnet19 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb net25 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net25 d i0#2fnet21 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net25 i0#2fseb i0#2fnet20 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_0P5

.subckt SAEDRVT14_FSDN8_V2_0P5 vdd vss vbp vbn q0 q1 q2 q3 q4 q5 q6 q7 qn0 qn1 qn2 qn3 qn4 qn5 qn6 qn7 ck d0 d1 d2 d3 d4 d5 d6 d7 si se
xi7 vdd vss vbp vbn q7 qn7 ck d7 si se SAEDRVT14_FSDN_V2_0P5
xi6 vdd vss vbp vbn q6 qn6 ck d6 si se SAEDRVT14_FSDN_V2_0P5
xi5 vdd vss vbp vbn q5 qn5 ck d5 si se SAEDRVT14_FSDN_V2_0P5
xi4 vdd vss vbp vbn q4 qn4 ck d4 si se SAEDRVT14_FSDN_V2_0P5
xi3 vdd vss vbp vbn q3 qn3 ck d3 si se SAEDRVT14_FSDN_V2_0P5
xi2 vdd vss vbp vbn q2 qn2 ck d2 si se SAEDRVT14_FSDN_V2_0P5
xi1 vdd vss vbp vbn q1 qn1 ck d1 si se SAEDRVT14_FSDN_V2_0P5
xi0 vdd vss vbp vbn q0 qn0 ck d0 si se SAEDRVT14_FSDN_V2_0P5
.ends SAEDRVT14_FSDN8_V2_0P5




.subckt SAEDRVT14_FSDN_V2_1 vdd vss vbp vbn q qn ck d si se
xmn1 ckbb ckb vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb net14 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 q qf_x vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net14 d i0#2fnet22 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net14 se i0#2fnet19 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb net25 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net25 d i0#2fnet21 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net25 i0#2fseb i0#2fnet20 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_1

.subckt SAEDRVT14_FSDN8_V2_1 vdd vss vbp vbn q0 q1 q2 q3 q4 q5 q6 q7 qn0 qn1 qn2 qn3 qn4 qn5 qn6 qn7 ck d0 d1 d2 d3 d4 d5 d6 d7 si se
xi7 vdd vss vbp vbn q7 qn7 ck d7 si se SAEDRVT14_FSDN_V2_1
xi6 vdd vss vbp vbn q6 qn6 ck d6 si se SAEDRVT14_FSDN_V2_1
xi5 vdd vss vbp vbn q5 qn5 ck d5 si se SAEDRVT14_FSDN_V2_1
xi4 vdd vss vbp vbn q4 qn4 ck d4 si se SAEDRVT14_FSDN_V2_1
xi3 vdd vss vbp vbn q3 qn3 ck d3 si se SAEDRVT14_FSDN_V2_1
xi2 vdd vss vbp vbn q2 qn2 ck d2 si se SAEDRVT14_FSDN_V2_1
xi1 vdd vss vbp vbn q1 qn1 ck d1 si se SAEDRVT14_FSDN_V2_1
xi0 vdd vss vbp vbn q0 qn0 ck d0 si se SAEDRVT14_FSDN_V2_1
.ends SAEDRVT14_FSDN8_V2_1




.subckt SAEDRVT14_FSDN_V2_2 vdd vss vbp vbn q qn ck d si se
xmn1 ckbb ckb vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_hvt l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb net017 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 q qf_x vss vbn n08_hvt l=0.014u nf=2 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_hvt l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net017 d i0#2fnet22 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net017 se i0#2fnet19 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_hvt l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb net019 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_hvt l=0.014u nf=2 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_hvt l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net019 d i0#2fnet21 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net019 i0#2fseb i0#2fnet20 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_2

.subckt SAEDRVT14_FSDN8_V2_2 vdd vss vbp vbn q0 q1 q2 q3 q4 q5 q6 q7 qn0 qn1 qn2 qn3 qn4 qn5 qn6 qn7 ck d0 d1 d2 d3 d4 d5 d6 d7 si se
xi7 vdd vss vbp vbn q7 qn7 ck d7 si se SAEDRVT14_FSDN_V2_2
xi6 vdd vss vbp vbn q6 qn6 ck d6 si se SAEDRVT14_FSDN_V2_2
xi5 vdd vss vbp vbn q5 qn5 ck d5 si se SAEDRVT14_FSDN_V2_2
xi4 vdd vss vbp vbn q4 qn4 ck d4 si se SAEDRVT14_FSDN_V2_2
xi3 vdd vss vbp vbn q3 qn3 ck d3 si se SAEDRVT14_FSDN_V2_2
xi2 vdd vss vbp vbn q2 qn2 ck d2 si se SAEDRVT14_FSDN_V2_2
xi1 vdd vss vbp vbn q1 qn1 ck d1 si se SAEDRVT14_FSDN_V2_2
xi0 vdd vss vbp vbn q0 qn0 ck d0 si se SAEDRVT14_FSDN_V2_2
.ends SAEDRVT14_FSDN8_V2_2




.subckt SAEDRVT14_FSDN_V2_4 vdd vss vbp vbn q qn ck d si se
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb net019 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net019 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net019 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb net017 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net017 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net017 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_4

.subckt SAEDRVT14_FSDN8_V2_4 vdd vss vbp vbn q0 q1 q2 q3 q4 q5 q6 q7 qn0 qn1 qn2 qn3 qn4 qn5 qn6 qn7 ck d0 d1 d2 d3 d4 d5 d6 d7 si se
xi7 vdd vss vbp vbn q7 qn7 ck d7 si se SAEDRVT14_FSDN_V2_4
xi6 vdd vss vbp vbn q6 qn6 ck d6 si se SAEDRVT14_FSDN_V2_4
xi5 vdd vss vbp vbn q5 qn5 ck d5 si se SAEDRVT14_FSDN_V2_4
xi4 vdd vss vbp vbn q4 qn4 ck d4 si se SAEDRVT14_FSDN_V2_4
xi3 vdd vss vbp vbn q3 qn3 ck d3 si se SAEDRVT14_FSDN_V2_4
xi2 vdd vss vbp vbn q2 qn2 ck d2 si se SAEDRVT14_FSDN_V2_4
xi1 vdd vss vbp vbn q1 qn1 ck d1 si se SAEDRVT14_FSDN_V2_4
xi0 vdd vss vbp vbn q0 qn0 ck d0 si se SAEDRVT14_FSDN_V2_4
.ends SAEDRVT14_FSDN8_V2_4




.subckt SAEDRVT14_FSDNQ_V3_1 vdd vss vbp vbn q ck d si se
xmibase#2fsltn1 mq_x ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 qf_x ckbb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq ckb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn5 i0#2fnet016 i0#2fseb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn4 net049 d i0#2fnet016 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 net049 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltp1 qf_x ckbb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf_x ckb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp5 ibase#2fnet41 ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckbb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp5 i0#2fnet015 se vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp4 net049 d i0#2fnet015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDNQ_V3_1




.subckt SAEDRVT14_FSDNQ_V3_2 vdd vss vbp vbn q ck d si se
xmibase#2fsltn1 mq_x ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf_x ckbb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn20 mq ckb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn5 i0#2fnet016 i0#2fseb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn4 net049 d i0#2fnet016 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 net049 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltp1 qf_x ckbb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp14 qf_x ckb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet41 ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckbb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp5 i0#2fnet015 se vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp4 net049 d i0#2fnet015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDNQ_V3_2




.subckt SAEDRVT14_FSDNQ_V3_4 vdd vss vbp vbn q ck d si se
xmibase#2fsltn1 mq_x ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf_x ckbb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn20 mq ckb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckbb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn5 i0#2fnet016 i0#2fseb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn4 net049 d i0#2fnet016 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 net049 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltp1 qf_x ckbb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp14 qf_x ckb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet41 ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckbb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp5 i0#2fnet015 se vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp4 net049 d i0#2fnet015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDNQ_V3_4




.subckt SAEDRVT14_FSDN_V2_0P5 vdd vss vbp vbn q qn ck d si se
xmn1 ckbb ckb vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb net14 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 q qf_x vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 qn qf vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net14 d i0#2fnet22 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net14 se i0#2fnet19 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb net25 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net25 d i0#2fnet21 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net25 i0#2fseb i0#2fnet20 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_0P5




.subckt SAEDRVT14_FSDPRBQ_V2_4 vdd vss vbp vbn q ck d si se rd
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPRBQ_V2_4




.subckt SAEDRVT14_FSDN_V2_2 vdd vss vbp vbn q qn ck d si se
xmn1 ckbb ckb vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_hvt l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb net017 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 q qf_x vss vbn n08_hvt l=0.014u nf=2 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_hvt l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net017 d i0#2fnet22 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net017 se i0#2fnet19 vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_hvt l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_hvt l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb net019 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_hvt l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_hvt l=0.014u nf=2 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_hvt l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net019 d i0#2fnet21 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net019 i0#2fseb i0#2fnet20 vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_hvt l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_2




.subckt SAEDRVT14_FSDN_V2_4 vdd vss vbp vbn q qn ck d si se
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckbb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckb net019 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckbb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net019 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net019 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckbb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckbb net017 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net017 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net017 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDN_V2_4




.subckt SAEDRVT14_FSDPMQ_0P5 vdd vss vbp vbn q ck d0 d1 s si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn22 i0#2fnet17 s i0#2fnet39 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn21 i0#2fnet39 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn16 net050 i0#2fseb i0#2fnet17 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn15 i0#2fenb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet17 i0#2fenb i0#2fnet35 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet35 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet36 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet36 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp20 i0#2fnet18 i0#2fenb i0#2fnet38 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp19 i0#2fnet38 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp14 net050 se i0#2fnet18 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp13 i0#2fenb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnet34 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet18 s i0#2fnet34 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 i0#2fseb i0#2fnet37 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet37 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPMQ_0P5




.subckt SAEDRVT14_FSDPMQ_1 vdd vss vbp vbn q ck d0 d1 s si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn22 i0#2fnet17 s i0#2fnet39 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn21 i0#2fnet39 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn16 net050 i0#2fseb i0#2fnet17 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn15 i0#2fenb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet17 i0#2fenb i0#2fnet35 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet35 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet36 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet36 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp20 i0#2fnet18 i0#2fenb i0#2fnet38 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp19 i0#2fnet38 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp14 net050 se i0#2fnet18 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp13 i0#2fenb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnet34 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet18 s i0#2fnet34 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 i0#2fseb i0#2fnet37 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet37 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPMQ_1




.subckt SAEDRVT14_FSDPMQ_2 vdd vss vbp vbn q ck d0 d1 s si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet030 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn22 i0#2fnet17 s i0#2fnet39 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn21 i0#2fnet39 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn16 net050 i0#2fseb i0#2fnet17 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn15 i0#2fenb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet17 i0#2fenb i0#2fnet35 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet35 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet36 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet36 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp20 i0#2fnet18 i0#2fenb i0#2fnet38 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp19 i0#2fnet38 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp14 net050 se i0#2fnet18 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp13 i0#2fenb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnet34 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet18 s i0#2fnet34 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 i0#2fseb i0#2fnet37 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet37 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPMQ_2




.subckt SAEDRVT14_FSDPMQ_4 vdd vss vbp vbn q ck d0 d1 s si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet030 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fn22 i0#2fnet17 s i0#2fnet39 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn21 i0#2fnet39 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn16 net050 i0#2fseb i0#2fnet17 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn15 i0#2fenb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet17 i0#2fenb i0#2fnet35 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet35 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet36 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet36 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fp20 i0#2fnet18 i0#2fenb i0#2fnet38 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp19 i0#2fnet38 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp14 net050 se i0#2fnet18 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp13 i0#2fenb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnet34 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet18 s i0#2fnet34 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 i0#2fseb i0#2fnet37 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet37 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPMQ_4




.subckt SAEDRVT14_FSDPMQ_LP_0P5 vdd vss vbp vbn q ck d0 d1 s si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn22 i0#2fnet17 s i0#2fnet39 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn21 i0#2fnet39 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn16 net050 i0#2fseb i0#2fnet17 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn15 i0#2fenb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet17 i0#2fenb i0#2fnet35 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet35 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet36 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet36 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp20 i0#2fnet18 i0#2fenb i0#2fnet38 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp19 i0#2fnet38 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp14 net050 se i0#2fnet18 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp13 i0#2fenb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnet34 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet18 s i0#2fnet34 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 i0#2fseb i0#2fnet37 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet37 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPMQ_LP_0P5




.subckt SAEDRVT14_FSDPMQ_LP_1 vdd vss vbp vbn q ck d0 d1 s si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn22 i0#2fnet17 s i0#2fnet39 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn21 i0#2fnet39 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn16 net050 i0#2fseb i0#2fnet17 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn15 i0#2fenb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet17 i0#2fenb i0#2fnet35 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet35 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet36 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet36 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp20 i0#2fnet18 i0#2fenb i0#2fnet38 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp19 i0#2fnet38 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp14 net050 se i0#2fnet18 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp13 i0#2fenb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnet34 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet18 s i0#2fnet34 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 i0#2fseb i0#2fnet37 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet37 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPMQ_LP_1




.subckt SAEDRVT14_FSDPMQ_LP_ vdd vss vbp vbn q ck d0 d1 s si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn22 i0#2fnet17 s i0#2fnet39 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn21 i0#2fnet39 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn16 net050 i0#2fseb i0#2fnet17 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn15 i0#2fenb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet17 i0#2fenb i0#2fnet35 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet35 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet36 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet36 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp20 i0#2fnet18 i0#2fenb i0#2fnet38 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp19 i0#2fnet38 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp14 net050 se i0#2fnet18 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp13 i0#2fenb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnet34 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet18 s i0#2fnet34 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 i0#2fseb i0#2fnet37 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet37 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPMQ_LP_1




.subckt SAEDRVT14_FSDPQB_V2_0P5 vdd vss vbp vbn qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net015 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net015 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPQB_V2_0P5




.subckt SAEDRVT14_FSDPQB_V2_1 vdd vss vbp vbn qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net015 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net015 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPQB_V2_1




.subckt SAEDRVT14_FSDPQB_V2_2 vdd vss vbp vbn qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net015 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net015 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPQB_V2_2




.subckt SAEDRVT14_FSDPQB_V2_4 vdd vss vbp vbn qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net015 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net015 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPQB_V2_4




.subckt SAEDRVT14_FSDPQB_V2_8 vdd vss vbp vbn qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp3 net015 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1 net015 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_FSDPQB_V2_8




.subckt SAEDRVT14_FSDPQB_V2_0P5 vdd vss vbp vbn qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net015 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net015 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPQB_V2_0P5




.subckt SAEDRVT14_FSDPQB_V2LP_1 vdd vss vbp vbn qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net015 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net015 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQB_V2LP_1




.subckt SAEDRVT14_FSDPQB_V2LP_2 vdd vss vbp vbn qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net015 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net015 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQB_V2LP_2




.subckt SAEDRVT14_FSDPQB_V3_1 vdd vss vbp vbn qn ck d si se
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 qf_x ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn5 i0#2fnet016 i0#2fseb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn4 net049 d i0#2fnet016 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 net049 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf_x ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp5 i0#2fnet015 se vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp4 net049 d i0#2fnet015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQB_V3_1




.subckt SAEDRVT14_FSDPQB_V3_2 vdd vss vbp vbn qn ck d si se
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 qf_x ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn5 i0#2fnet016 i0#2fseb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn4 net049 d i0#2fnet016 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 net049 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf_x ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp5 i0#2fnet015 se vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp4 net049 d i0#2fnet015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQB_V3_2




.subckt SAEDRVT14_FSDPQB_V3_4 vdd vss vbp vbn qn ck d si se
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf_x ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn5 i0#2fnet016 i0#2fseb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn4 net049 d i0#2fnet016 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 net049 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf_x ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp5 i0#2fnet015 se vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp4 net049 d i0#2fnet015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQB_V3_4




.subckt SAEDRVT14_FSDPQB_V3_8 vdd vss vbp vbn qn ck d si se
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf_x ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn5 i0#2fnet016 i0#2fseb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn4 net049 d i0#2fnet016 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 net049 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf_x ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp5 i0#2fnet015 se vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp4 net049 d i0#2fnet015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQB_V3_8




.subckt SAEDRVT14_FSDPQM4_V2LPY2_1 vdd vss q0 q1 q2 q3 ck d0 d1 d2 d3 si se
xn0 ckb ck vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn0 ckbb ckb vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xibase#2fn13 ibase#2fnet046 qf0 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn12 mq0 ckbb ibase#2fnet048 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn11 ibase#2fnet048 mq_x0 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn10 mq_x0 mq0 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn9 sfbn ckb ibase#2fnet046 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn8 qf0 sfbn vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn6 mq0 ckb ibase#2fnet028 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn5 mq_x0 ckbb sfbn vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn0 ibase#2fnet028 net050 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi37#2fn0 q3 sfbn_3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi36#2fn13 i36#2fnet046 qf3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn12 mq3 ckbb i36#2fnet048 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn11 i36#2fnet048 mq_x3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn10 mq_x3 mq3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn9 sfbn_3 ckb i36#2fnet046 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn8 qf3 sfbn_3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn6 mq3 ckb i36#2fnet028 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn5 mq_x3 ckbb sfbn_3 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn0 i36#2fnet028 net027 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn17 i35#2fseb se vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmn3 net027 i35#2fseb i35#2fnet22 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmn2 i35#2fnet22 d3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmn1 net027 se i35#2fnet19 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmn0 i35#2fnet19 qf2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn17 i34#2fseb se vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmn3 net028 i34#2fseb i34#2fnet22 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmn2 i34#2fnet22 d2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmn1 net028 se i34#2fnet19 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmn0 i34#2fnet19 qf1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn13 i33#2fnet046 qf2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn12 mq2 ckbb i33#2fnet048 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn11 i33#2fnet048 mq_x2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn10 mq_x2 mq2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn9 sfbn_2 ckb i33#2fnet046 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn8 qf2 sfbn_2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn6 mq2 ckb i33#2fnet028 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn5 mq_x2 ckbb sfbn_2 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn0 i33#2fnet028 net028 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fn0 q2 sfbn_2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi31#2fn0 q1 sfbn_1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi30#2fn13 i30#2fnet046 qf1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn12 mq1 ckbb i30#2fnet048 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn11 i30#2fnet048 mq_x1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn10 mq_x1 mq1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn9 sfbn_1 ckb i30#2fnet046 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn8 qf1 sfbn_1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn6 mq1 ckb i30#2fnet028 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn5 mq_x1 ckbb sfbn_1 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn0 i30#2fnet028 net029 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn17 i29#2fseb se vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmn3 net029 i29#2fseb i29#2fnet22 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmn2 i29#2fnet22 d1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmn1 net029 se i29#2fnet19 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmn0 i29#2fnet19 qf0 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fn0 q0 sfbn vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn17 i0#2fseb se vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmn3 net050 i0#2fseb i0#2fnet22 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmn2 i0#2fnet22 d0 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmn1 net050 se i0#2fnet19 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmn0 i0#2fnet19 si vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xp0 ckb ck vdd vdd p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp0 ckbb ckb vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xibase#2fp11 ibase#2fnet045 qf0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp10 mq0 ckb ibase#2fnet047 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp9 ibase#2fnet047 mq_x0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp8 mq_x0 mq0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp7 sfbn ckbb ibase#2fnet045 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp6 qf0 sfbn vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp4 mq0 ckbb ibase#2fnet027 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp3 sfbn ckb mq_x0 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp1 ibase#2fnet027 net050 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi37#2fp1 q3 sfbn_3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi36#2fp11 i36#2fnet045 qf3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp10 mq3 ckb i36#2fnet047 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp9 i36#2fnet047 mq_x3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp8 mq_x3 mq3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp7 sfbn_3 ckbb i36#2fnet045 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp6 qf3 sfbn_3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp4 mq3 ckbb i36#2fnet027 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp3 sfbn_3 ckb mq_x3 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp1 i36#2fnet027 net027 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fp15 i35#2fseb se vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmp3 net027 se i35#2fnet21 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmp2 i35#2fnet21 d3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmp1 net027 i35#2fseb i35#2fnet20 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmp0 i35#2fnet20 qf2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fp15 i34#2fseb se vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmp3 net028 se i34#2fnet21 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmp2 i34#2fnet21 d2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmp1 net028 i34#2fseb i34#2fnet20 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmp0 i34#2fnet20 qf1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp11 i33#2fnet045 qf2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp10 mq2 ckb i33#2fnet047 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp9 i33#2fnet047 mq_x2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp8 mq_x2 mq2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp7 sfbn_2 ckbb i33#2fnet045 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp6 qf2 sfbn_2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp4 mq2 ckbb i33#2fnet027 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp3 sfbn_2 ckb mq_x2 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp1 i33#2fnet027 net028 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fp1 q2 sfbn_2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi31#2fp1 q1 sfbn_1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi30#2fp11 i30#2fnet045 qf1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp10 mq1 ckb i30#2fnet047 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp9 i30#2fnet047 mq_x1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp8 mq_x1 mq1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp7 sfbn_1 ckbb i30#2fnet045 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp6 qf1 sfbn_1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp4 mq1 ckbb i30#2fnet027 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp3 sfbn_1 ckb mq_x1 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp1 i30#2fnet027 net029 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fp15 i29#2fseb se vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmp3 net029 se i29#2fnet21 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmp2 i29#2fnet21 d1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmp1 net029 i29#2fseb i29#2fnet20 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmp0 i29#2fnet20 qf0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fp1 q0 sfbn vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp15 i0#2fseb se vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmp3 net050 se i0#2fnet21 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmp2 i0#2fnet21 d0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmp1 net050 i0#2fseb i0#2fnet20 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmp0 i0#2fnet20 si vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
.ends SAEDRVT14_FSDPQM4_V2LPY2_1




.subckt SAEDRVT14_FSDPQM4_V2Y2_1 vdd vss vbp vbn q0 q1 q2 q3 ck d0 d1 d2 d3 si se
xn0 ckb ck vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xmn0 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xibase#2fn13 ibase#2fnet046 qf0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn12 mq0 ckbb ibase#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn11 ibase#2fnet048 mq_x0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn10 mq_x0 mq0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn9 sfbn ckb ibase#2fnet046 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn8 qf0 sfbn vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn6 mq0 ckb ibase#2fnet028 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn5 mq_x0 ckbb sfbn vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi37#2fn0 q3 sfbn_3 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi36#2fn13 i36#2fnet046 qf3 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn12 mq3 ckbb i36#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn11 i36#2fnet048 mq_x3 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn10 mq_x3 mq3 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn9 sfbn_3 ckb i36#2fnet046 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn8 qf3 sfbn_3 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn6 mq3 ckb i36#2fnet028 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn5 mq_x3 ckbb sfbn_3 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn0 i36#2fnet028 net027 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn17 i35#2fseb se vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmn3 net027 i35#2fseb i35#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmn2 i35#2fnet22 d3 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmn1 net027 se i35#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmn0 i35#2fnet19 qf2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn17 i34#2fseb se vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmn3 net028 i34#2fseb i34#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmn2 i34#2fnet22 d2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmn1 net028 se i34#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmn0 i34#2fnet19 qf1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn13 i33#2fnet046 qf2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn12 mq2 ckbb i33#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn11 i33#2fnet048 mq_x2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn10 mq_x2 mq2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn9 sfbn_2 ckb i33#2fnet046 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn8 qf2 sfbn_2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn6 mq2 ckb i33#2fnet028 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn5 mq_x2 ckbb sfbn_2 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn0 i33#2fnet028 net028 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fn0 q2 sfbn_2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi31#2fn0 q1 sfbn_1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi30#2fn13 i30#2fnet046 qf1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn12 mq1 ckbb i30#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn11 i30#2fnet048 mq_x1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn10 mq_x1 mq1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn9 sfbn_1 ckb i30#2fnet046 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn8 qf1 sfbn_1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn6 mq1 ckb i30#2fnet028 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn5 mq_x1 ckbb sfbn_1 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn0 i30#2fnet028 net029 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn17 i29#2fseb se vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmn3 net029 i29#2fseb i29#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmn2 i29#2fnet22 d1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmn1 net029 se i29#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmn0 i29#2fnet19 qf0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fn0 q0 sfbn vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn17 i0#2fseb se vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmn3 net050 i0#2fseb i0#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmn2 i0#2fnet22 d0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmn0 i0#2fnet19 si vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xp0 ckb ck vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xmp0 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xibase#2fp11 ibase#2fnet045 qf0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp10 mq0 ckb ibase#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp9 ibase#2fnet047 mq_x0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp8 mq_x0 mq0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp7 sfbn ckbb ibase#2fnet045 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp6 qf0 sfbn vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp4 mq0 ckbb ibase#2fnet027 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp3 sfbn ckb mq_x0 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi37#2fp1 q3 sfbn_3 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi36#2fp11 i36#2fnet045 qf3 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp10 mq3 ckb i36#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp9 i36#2fnet047 mq_x3 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp8 mq_x3 mq3 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp7 sfbn_3 ckbb i36#2fnet045 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp6 qf3 sfbn_3 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp4 mq3 ckbb i36#2fnet027 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp3 sfbn_3 ckb mq_x3 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp1 i36#2fnet027 net027 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fp15 i35#2fseb se vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmp3 net027 se i35#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmp2 i35#2fnet21 d3 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmp1 net027 i35#2fseb i35#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fmp0 i35#2fnet20 qf2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fp15 i34#2fseb se vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmp3 net028 se i34#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmp2 i34#2fnet21 d2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmp1 net028 i34#2fseb i34#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fmp0 i34#2fnet20 qf1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp11 i33#2fnet045 qf2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp10 mq2 ckb i33#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp9 i33#2fnet047 mq_x2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp8 mq_x2 mq2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp7 sfbn_2 ckbb i33#2fnet045 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp6 qf2 sfbn_2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp4 mq2 ckbb i33#2fnet027 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp3 sfbn_2 ckb mq_x2 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp1 i33#2fnet027 net028 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fp1 q2 sfbn_2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi31#2fp1 q1 sfbn_1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi30#2fp11 i30#2fnet045 qf1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp10 mq1 ckb i30#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp9 i30#2fnet047 mq_x1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp8 mq_x1 mq1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp7 sfbn_1 ckbb i30#2fnet045 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp6 qf1 sfbn_1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp4 mq1 ckbb i30#2fnet027 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp3 sfbn_1 ckb mq_x1 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp1 i30#2fnet027 net029 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fp15 i29#2fseb se vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmp3 net029 se i29#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmp2 i29#2fnet21 d1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmp1 net029 i29#2fseb i29#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fmp0 i29#2fnet20 qf0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fp1 q0 sfbn vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp15 i0#2fseb se vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmp3 net050 se i0#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmp2 i0#2fnet21 d0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmp1 net050 i0#2fseb i0#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
.ends SAEDRVT14_FSDPQM4_V2Y2_1




.subckt SAEDRVT14_FSDPQ_V2_0P5 vdd vss vbp vbn q ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 i0#2fseb i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net050 se i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net050 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQ_V2_0P5




.subckt SAEDRVT14_FSDPQ_V2_1 vdd vss vbp vbn q ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 i0#2fseb i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net050 se i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net050 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQ_V2_1



.subckt SAEDRVT14_FSDPQ_V2_2 vdd vss vbp vbn q ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 i0#2fseb i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net050 se i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net050 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQ_V2_2




.subckt SAEDRVT14_FSDPQ_V2_4 vdd vss vbp vbn q ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet030 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 i0#2fseb i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net050 se i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net050 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQ_V2_4




.subckt SAEDRVT14_FSDPQ_V2LP_0P5 vdd vss vbp vbn q ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 i0#2fseb i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net050 se i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net050 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQ_V2LP_0P5




.subckt SAEDRVT14_FSDPQ_V2LP_1 vdd vss vbp vbn q ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 i0#2fseb i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net050 se i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net050 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQ_V2LP_1




.subckt SAEDRVT14_FSDPQ_V2LP_2 vdd vss vbp vbn q ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 i0#2fseb i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net050 se i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net050 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQ_V2LP_2




.subckt SAEDRVT14_FSDPQ_V3_1 vdd vss vbp vbn q ck d si se
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 qf_x ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn5 i0#2fnet016 i0#2fseb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn4 net049 d i0#2fnet016 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 net049 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf_x ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp5 i0#2fnet015 se vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp4 net049 d i0#2fnet015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQ_V3_1




.subckt SAEDRVT14_FSDPQ_V3_2 vdd vss vbp vbn q ck d si se
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf_x ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn5 i0#2fnet016 i0#2fseb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn4 net049 d i0#2fnet016 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 net049 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp14 qf_x ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp5 i0#2fnet015 se vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp4 net049 d i0#2fnet015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQ_V3_2




.subckt SAEDRVT14_FSDPQ_V3_4 vdd vss vbp vbn q ck d si se
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf_x ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn5 i0#2fnet016 i0#2fseb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn4 net049 d i0#2fnet016 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 net049 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp14 qf_x ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp5 i0#2fnet015 se vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp4 net049 d i0#2fnet015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPQ_V3_4




.subckt SAEDRVT14_FSDPRBQ_V2_0P5 vdd vss vbp vbn q ck d si se rd
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPRBQ_V2_0P5




.subckt SAEDRVT14_FSDPRBQ_V2_1 vdd vss vbp vbn q ck d si se rd
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPRBQ_V2_1




.subckt SAEDRVT14_FSDPRBQ_V2_2 vdd vss vbp vbn q ck d si se rd
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPRBQ_V2_2




.subckt SAEDRVT14_FSDPRBQ_V2_4 vdd vss vbp vbn q ck d si se rd
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPRBQ_V2_4




.subckt SAEDRVT14_FSDPRBQ_V2LP_0P5 vdd vss vbp vbn q ck d si se rd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPRBQ_V2LP_0P5




.subckt SAEDRVT14_FSDPRBQ_V2LP_1 vdd vss vbp vbn q ck d si se rd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPRBQ_V2LP_1




.subckt SAEDRVT14_FSDPRBQ_V2LP_2 vdd vss vbp vbn q ck d si se rd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet14 mq ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 qf ckb ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet31 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn4 ibase#2fnet14 ckbb mq_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 qf_x qf ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet015 ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet015 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet015 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet42 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet42 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 qf_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPRBQ_V2LP_2




.subckt SAEDRVT14_FSDPRBQ_V3_1 vdd vss vbp vbn q ck d si se rd
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn32 ibase#2fnet025 ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn31 ibase#2fnet025 qf ibase#2fnet031 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn30 ibase#2fnet031 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn21 ibase#2fnet032 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq ibase#2fnet032 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn5 i0#2fnet016 i0#2fseb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn4 net049 d i0#2fnet016 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 net049 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp31 qf_x ckbb ibase#2fnet025 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp30 ibase#2fnet025 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp29 ibase#2fnet025 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp21 mq_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp5 i0#2fnet015 se vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp4 net049 d i0#2fnet015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPRBQ_V3_1




.subckt SAEDRVT14_FSDPRBQ_V3_2 vdd vss vbp vbn q ck d si se rd
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn32 ibase#2fnet025 ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn31 ibase#2fnet025 qf ibase#2fnet031 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn30 ibase#2fnet031 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet038 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn21 ibase#2fnet032 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq ibase#2fnet032 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet038 ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn5 i0#2fnet016 i0#2fseb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn4 net049 d i0#2fnet016 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 net049 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp31 qf_x ckbb ibase#2fnet025 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp30 ibase#2fnet025 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp29 ibase#2fnet025 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet037 ckbb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp21 mq_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmp17 mq net049 ibase#2fnet037 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp5 i0#2fnet015 se vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp4 net049 d i0#2fnet015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPRBQ_V3_2




.subckt SAEDRVT14_FSDPRBQ_V3_4 vdd vss vbp vbn q ck d si se rd
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn32 ibase#2fnet025 ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn31 ibase#2fnet025 qf ibase#2fnet031 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn30 ibase#2fnet031 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet038 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn21_2 ibase#2fnet032_2 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn18_2 mq_x mq ibase#2fnet032_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn21 ibase#2fnet032 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq ibase#2fnet032 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet038 ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn5 i0#2fnet016 i0#2fseb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmn4 net049 d i0#2fnet016 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 net049 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp31 qf_x ckbb ibase#2fnet025 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp30 ibase#2fnet025 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp29 ibase#2fnet025 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet037 ckbb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp21 mq_x rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp17 mq net049 ibase#2fnet037 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp5 i0#2fnet015 se vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fmp4 net049 d i0#2fnet015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPRBQ_V3_4




.subckt SAEDRVT14_FSDPRBSBQ_V2_0P5 vdd vss vbp vbn q ck d si se rd sd
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 i2 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet038 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet038 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 i1 ckb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net10 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net10 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp26 ibase#2fnet016 ckb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckbb ibase#2fnet026 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 ibase#2fnet026 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 i98 ckb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 ibase#2fnet026 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 i1 ckbb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net11 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net11 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPRBSBQ_V2_0P5




.subckt SAEDRVT14_FSDPRBSBQ_V2_1 vdd vss vbp vbn q ck d si se rd sd
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn8 i2 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet038 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet038 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn1 i1 ckb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net10 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net10 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp26 ibase#2fnet016 ckb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckbb ibase#2fnet026 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 ibase#2fnet026 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 i98 ckb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 ibase#2fnet026 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 i1 ckbb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net11 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net11 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPRBSBQ_V2_1




.subckt SAEDRVT14_FSDPRBSBQ_V2_2 vdd vss vbp vbn q ck d si se rd sd
xmibase#2fn9_1 ibase#2fnet43_1 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn2_1 i99 i98 ibase#2fnet43_1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn8 i2 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet027 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet027 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn1 i1 ckb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net10 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net10 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp26 ibase#2fnet016 ckb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckbb ibase#2fnet026 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 ibase#2fnet026 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 i98 ckb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 ibase#2fnet026 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 i1 ckbb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net11 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net11 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPRBSBQ_V2_2




.subckt SAEDRVT14_FSDPRBSBQ_V2_4 vdd vss vbp vbn q ck d si se rd sd
xmibase#2fn9_1 ibase#2fnet43_1 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn2_1 i99 i98 ibase#2fnet43_1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn8 i2 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet027 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet027 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn4 ibase#2fnet14 ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn1 i1 ckb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net10 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net10 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp26 ibase#2fnet016 ckb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckbb ibase#2fnet026 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 ibase#2fnet026 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 i98 ckb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 ibase#2fnet026 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 i1 ckbb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net11 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net11 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPRBSBQ_V2_4




.subckt SAEDRVT14_FSDPRBSBQ_V2LP_0P5 vdd vss vbp vbn q ck d si se rd sd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 i2 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet027 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet027 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn4 ibase#2fnet14 ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 i1 ckb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net10 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net10 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet016 ckb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckbb ibase#2fnet039 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 ibase#2fnet039 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 i98 ckb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 ibase#2fnet039 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 i1 ckbb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net11 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net11 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPRBSBQ_V2LP_0P5




.subckt SAEDRVT14_FSDPRBSBQ_V2LP_1 vdd vss vbp vbn q ck d si se rd sd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 i2 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet027 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet027 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn4 ibase#2fnet14 ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 i1 ckb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net10 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net10 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet016 ckb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckbb ibase#2fnet039 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 ibase#2fnet039 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 i98 ckb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 ibase#2fnet039 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 i1 ckbb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net11 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net11 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPRBSBQ_V2LP_1




.subckt SAEDRVT14_FSDPRBSBQ_V2LP_2 vdd vss vbp vbn q ck d si se rd sd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet14 i2 ibase#2fnet44 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 ibase#2fnet035 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 ibase#2fnet43 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 i2 ckbb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 ibase#2fnet027 ckb i98 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 ibase#2fnet027 i99 ibase#2fnet035 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 i2 i1 ibase#2fnet034 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn4 ibase#2fnet14 ckbb i1 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn3 ibase#2fnet44 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn2 i99 i98 ibase#2fnet43 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 i1 ckb net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet034 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q i99 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net10 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net10 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp26 ibase#2fnet016 ckb i1 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp25 ibase#2fnet016 i2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp24 ibase#2fnet016 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 i98 ckbb ibase#2fnet039 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 ibase#2fnet039 i99 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 i99 i98 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 i2 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 i98 ckb i2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 ibase#2fnet039 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 i1 ckbb net11 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 i99 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp0 i2 i1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q i99 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net11 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net11 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPRBSBQ_V2LP_2




.subckt SAEDRVT14_FSDPSBQ_V2_0P5 vdd vss vbp vbn q ck d si se sd
xmibase#2fp23 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp22 ibase#2fnet025 ckbb qf vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp20 mq sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp19 ibase#2fnet025 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet025 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp10 mq_x ckb ibase#2fnet31 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet31 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn25 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn24 ibase#2fnet24 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet33 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn22 mq mq_x ibase#2fnet33 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 ibase#2fnet30 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet24 qf_x ibase#2fnet30 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet32 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPSBQ_V2_0P5




.subckt SAEDRVT14_FSDPSBQ_V2_1 vdd vss vbp vbn q ck d si se sd
xmibase#2fp23 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp22 ibase#2fnet025 ckbb qf vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp20 mq sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp19 ibase#2fnet025 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet025 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp10 mq_x ckb ibase#2fnet31 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet31 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn25 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn24 ibase#2fnet24 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet33 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn22 mq mq_x ibase#2fnet33 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 ibase#2fnet30 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet24 qf_x ibase#2fnet30 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet32 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPSBQ_V2_1




.subckt SAEDRVT14_FSDPSBQ_V2_2 vdd vss vbp vbn q ck d si se sd
xmibase#2fp23 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp22 ibase#2fnet025 ckbb qf vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp20 mq sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp19 ibase#2fnet025 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp11 ibase#2fnet025 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp10 mq_x ckb ibase#2fnet31 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet31 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn25 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn24 ibase#2fnet24 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet33 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn22 mq mq_x ibase#2fnet33 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 ibase#2fnet30 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn13 ibase#2fnet24 qf_x ibase#2fnet30 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn12 mq_x ckbb ibase#2fnet32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet32 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPSBQ_V2_2




.subckt SAEDRVT14_FSDPSBQ_V2_4 vdd vss vbp vbn q ck d si se sd
xmibase#2fp23 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp22 ibase#2fnet025 ckbb qf vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp20 mq sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp19 ibase#2fnet025 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp11 ibase#2fnet025 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp10 mq_x ckb ibase#2fnet31 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet31 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn25 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn24 ibase#2fnet24 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet33 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn22 mq mq_x ibase#2fnet33 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 ibase#2fnet30 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn13 ibase#2fnet24 qf_x ibase#2fnet30 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn12 mq_x ckbb ibase#2fnet32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet32 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDPSBQ_V2_4




.subckt SAEDRVT14_FSDPSBQ_V2LP_0P5 vdd vss vbp vbn q ck d si se sd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn25 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn24 ibase#2fnet24 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet33 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn22 mq mq_x ibase#2fnet33 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn17 ibase#2fnet30 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet24 qf_x ibase#2fnet30 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet32 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp23 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp22 ibase#2fnet025 ckbb qf vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp20 mq sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp19 ibase#2fnet025 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet025 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet31 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet31 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSBQ_V2LP_0P5




.subckt SAEDRVT14_FSDPSBQ_V2LP_1 vdd vss vbp vbn q ck d si se sd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn25 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn24 ibase#2fnet24 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet33 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn22 mq mq_x ibase#2fnet33 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn17 ibase#2fnet30 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet24 qf_x ibase#2fnet30 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet32 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp23 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp22 ibase#2fnet025 ckbb qf vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp20 mq sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp19 ibase#2fnet025 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet025 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet31 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet31 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSBQ_V2LP_1




.subckt SAEDRVT14_FSDPSBQ_V2LP_2 vdd vss vbp vbn q ck d si se sd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn25 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn24 ibase#2fnet24 ckb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn23 ibase#2fnet33 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn22 mq mq_x ibase#2fnet33 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn17 ibase#2fnet30 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet24 qf_x ibase#2fnet30 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet32 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn1 mq_x ckb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net050 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net050 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp23 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp22 ibase#2fnet025 ckbb qf vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp20 mq sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp19 ibase#2fnet025 sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet025 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet31 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet31 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp2 mq_x ckbb net049 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net049 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net049 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSBQ_V2LP_2




.subckt SAEDRVT14_FSDPSYNRBQM4_V2LPY2_1 vdd vss q0 q1 q2 q3 ck d0 d1 d2 d3 si se rd
xn0 ckb ck vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=2
xmn0 ckbb ckb vss vss n08_rev l=0.014u nf=2 m=1 nfin=2
xibase#2fn13 ibase#2fnet046 qf0 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn12 mq0 ckbb ibase#2fnet048 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn11 ibase#2fnet048 mq_x0 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn10 mq_x0 mq0 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn9 sfbn ckb ibase#2fnet046 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn8 qf0 sfbn vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn6 mq0 ckb ibase#2fnet028 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn5 mq_x0 ckbb sfbn vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn0 ibase#2fnet028 net050 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi37#2fn0 q3 sfbn_3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi36#2fn13 i36#2fnet046 qf3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn12 mq3 ckbb i36#2fnet048 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn11 i36#2fnet048 mq_x3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn10 mq_x3 mq3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn9 sfbn_3 ckb i36#2fnet046 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn8 qf3 sfbn_3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn6 mq3 ckb i36#2fnet028 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn5 mq_x3 ckbb sfbn_3 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn0 i36#2fnet028 net021 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn17 i35#2fseb se vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn14 i35#2fnet23 rd vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn4 i35#2fnd_out d3 i35#2fnet23 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn3 i35#2fnd_out i35#2fseb net021 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn2 i35#2fnet21 qf2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn0 net021 se i35#2fnet21 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn17 i34#2fseb se vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn14 i34#2fnet23 rd vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn4 i34#2fnd_out d2 i34#2fnet23 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn3 i34#2fnd_out i34#2fseb net020 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn2 i34#2fnet21 qf1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn0 net020 se i34#2fnet21 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn13 i33#2fnet046 qf2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn12 mq2 ckbb i33#2fnet048 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn11 i33#2fnet048 mq_x2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn10 mq_x2 mq2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn9 sfbn_2 ckb i33#2fnet046 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn8 qf2 sfbn_2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn6 mq2 ckb i33#2fnet028 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn5 mq_x2 ckbb sfbn_2 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn0 i33#2fnet028 net020 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fn0 q2 sfbn_2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi31#2fn0 q1 sfbn_1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi30#2fn13 i30#2fnet046 qf1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn12 mq1 ckbb i30#2fnet048 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn11 i30#2fnet048 mq_x1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn10 mq_x1 mq1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn9 sfbn_1 ckb i30#2fnet046 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn8 qf1 sfbn_1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn6 mq1 ckb i30#2fnet028 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn5 mq_x1 ckbb sfbn_1 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn0 i30#2fnet028 net019 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn17 i29#2fseb se vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn14 i29#2fnet23 rd vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn4 i29#2fnd_out d1 i29#2fnet23 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn3 i29#2fnd_out i29#2fseb net019 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn2 i29#2fnet21 qf0 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn0 net019 se i29#2fnet21 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fn0 q0 sfbn vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn17 i0#2fseb se vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn14 i0#2fnet23 rd vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn4 i0#2fnd_out d0 i0#2fnet23 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn3 i0#2fnd_out i0#2fseb net050 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn2 i0#2fnet21 si vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn0 net050 se i0#2fnet21 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xp0 ckb ck vdd vdd p08_rev2 l=0.014u nf=2 m=1 nfin=2
xmp0 ckbb ckb vdd vdd p08_rev l=0.014u nf=2 m=1 nfin=2
xibase#2fp11 ibase#2fnet045 qf0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp10 mq0 ckb ibase#2fnet047 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp9 ibase#2fnet047 mq_x0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp8 mq_x0 mq0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp7 sfbn ckbb ibase#2fnet045 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp6 qf0 sfbn vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp4 mq0 ckbb ibase#2fnet027 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp3 sfbn ckb mq_x0 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp1 ibase#2fnet027 net050 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi37#2fp1 q3 sfbn_3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi36#2fp11 i36#2fnet045 qf3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp10 mq3 ckb i36#2fnet047 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp9 i36#2fnet047 mq_x3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp8 mq_x3 mq3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp7 sfbn_3 ckbb i36#2fnet045 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp6 qf3 sfbn_3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp4 mq3 ckbb i36#2fnet027 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp3 sfbn_3 ckb mq_x3 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp1 i36#2fnet027 net021 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fp15 i35#2fseb se vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fp12 i35#2fnd_out d3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fp3 net021 i35#2fseb i35#2fnet22 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fp2 i35#2fnd_out rd vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fp1 net021 se i35#2fnd_out vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fp0 i35#2fnet22 qf2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fp15 i34#2fseb se vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fp12 i34#2fnd_out d2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fp3 net020 i34#2fseb i34#2fnet22 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fp2 i34#2fnd_out rd vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fp1 net020 se i34#2fnd_out vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fp0 i34#2fnet22 qf1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp11 i33#2fnet045 qf2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp10 mq2 ckb i33#2fnet047 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp9 i33#2fnet047 mq_x2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp8 mq_x2 mq2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp7 sfbn_2 ckbb i33#2fnet045 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp6 qf2 sfbn_2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp4 mq2 ckbb i33#2fnet027 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp3 sfbn_2 ckb mq_x2 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp1 i33#2fnet027 net020 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fp1 q2 sfbn_2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi31#2fp1 q1 sfbn_1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi30#2fp11 i30#2fnet045 qf1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp10 mq1 ckb i30#2fnet047 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp9 i30#2fnet047 mq_x1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp8 mq_x1 mq1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp7 sfbn_1 ckbb i30#2fnet045 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp6 qf1 sfbn_1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp4 mq1 ckbb i30#2fnet027 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp3 sfbn_1 ckb mq_x1 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp1 i30#2fnet027 net019 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fp15 i29#2fseb se vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fp12 i29#2fnd_out d1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fp3 net019 i29#2fseb i29#2fnet22 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fp2 i29#2fnd_out rd vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fp1 net019 se i29#2fnd_out vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fp0 i29#2fnet22 qf0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fp1 q0 sfbn vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp15 i0#2fseb se vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp12 i0#2fnd_out d0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp3 net050 i0#2fseb i0#2fnet22 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp2 i0#2fnd_out rd vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp1 net050 se i0#2fnd_out vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp0 i0#2fnet22 si vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
.ends SAEDRVT14_FSDPSYNRBQM4_V2LPY2_1




.subckt SAEDRVT14_FSDPSYNRBQM4_V2Y2_1 vdd vss q0 q1 q2 q3 ck d0 d1 d2 d3 si se rd
xn0 ckb ck vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xmn0 ckbb ckb vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xibase#2fn13 ibase#2fnet046 qf0 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn12 mq0 ckbb ibase#2fnet048 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn11 ibase#2fnet048 mq_x0 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn10 mq_x0 mq0 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn9 sfbn ckb ibase#2fnet046 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn8 qf0 sfbn vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn6 mq0 ckb ibase#2fnet028 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn5 mq_x0 ckbb sfbn vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fn0 ibase#2fnet028 net050 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi37#2fn0 q3 sfbn_3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi36#2fn13 i36#2fnet046 qf3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn12 mq3 ckbb i36#2fnet048 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn11 i36#2fnet048 mq_x3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn10 mq_x3 mq3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn9 sfbn_3 ckb i36#2fnet046 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn8 qf3 sfbn_3 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn6 mq3 ckb i36#2fnet028 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn5 mq_x3 ckbb sfbn_3 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fn0 i36#2fnet028 net021 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn17 i35#2fseb se vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn14 i35#2fnet23 rd vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn4 i35#2fnd_out d3 i35#2fnet23 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn3 i35#2fnd_out i35#2fseb net021 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn2 i35#2fnet21 qf2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn0 net021 se i35#2fnet21 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn17 i34#2fseb se vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn14 i34#2fnet23 rd vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn4 i34#2fnd_out d2 i34#2fnet23 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn3 i34#2fnd_out i34#2fseb net020 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn2 i34#2fnet21 qf1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn0 net020 se i34#2fnet21 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn13 i33#2fnet046 qf2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn12 mq2 ckbb i33#2fnet048 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn11 i33#2fnet048 mq_x2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn10 mq_x2 mq2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn9 sfbn_2 ckb i33#2fnet046 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn8 qf2 sfbn_2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn6 mq2 ckb i33#2fnet028 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn5 mq_x2 ckbb sfbn_2 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fn0 i33#2fnet028 net020 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fn0 q2 sfbn_2 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi31#2fn0 q1 sfbn_1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi30#2fn13 i30#2fnet046 qf1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn12 mq1 ckbb i30#2fnet048 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn11 i30#2fnet048 mq_x1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn10 mq_x1 mq1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn9 sfbn_1 ckb i30#2fnet046 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn8 qf1 sfbn_1 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn6 mq1 ckb i30#2fnet028 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn5 mq_x1 ckbb sfbn_1 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fn0 i30#2fnet028 net019 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn17 i29#2fseb se vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn14 i29#2fnet23 rd vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn4 i29#2fnd_out d1 i29#2fnet23 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn3 i29#2fnd_out i29#2fseb net019 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn2 i29#2fnet21 qf0 vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn0 net019 se i29#2fnet21 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fn0 q0 sfbn vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn17 i0#2fseb se vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn14 i0#2fnet23 rd vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn4 i0#2fnd_out d0 i0#2fnet23 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn3 i0#2fnd_out i0#2fseb net050 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn2 i0#2fnet21 si vss vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn0 net050 se i0#2fnet21 vss n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xp0 ckb ck vdd vdd p08_rev2 l=0.014u nf=2 m=1 nfin=4
xmp0 ckbb ckb vdd vdd p08_rev l=0.014u nf=2 m=1 nfin=4
xibase#2fp11 ibase#2fnet045 qf0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp10 mq0 ckb ibase#2fnet047 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp9 ibase#2fnet047 mq_x0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp8 mq_x0 mq0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp7 sfbn ckbb ibase#2fnet045 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp6 qf0 sfbn vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp4 mq0 ckbb ibase#2fnet027 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp3 sfbn ckb mq_x0 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xibase#2fp1 ibase#2fnet027 net050 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi37#2fp1 q3 sfbn_3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi36#2fp11 i36#2fnet045 qf3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp10 mq3 ckb i36#2fnet047 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp9 i36#2fnet047 mq_x3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp8 mq_x3 mq3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp7 sfbn_3 ckbb i36#2fnet045 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp6 qf3 sfbn_3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp4 mq3 ckbb i36#2fnet027 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp3 sfbn_3 ckb mq_x3 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi36#2fp1 i36#2fnet027 net021 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fp15 i35#2fseb se vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fp12 i35#2fnd_out d3 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fp2 i35#2fnd_out rd vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fp1 net021 se i35#2fnd_out vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fp0 i35#2fnet22 qf2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi35#2fn1 net021 i35#2fseb i35#2fnet22 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fp15 i34#2fseb se vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fp12 i34#2fnd_out d2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fp2 i34#2fnd_out rd vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fp1 net020 se i34#2fnd_out vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fp0 i34#2fnet22 qf1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi34#2fn1 net020 i34#2fseb i34#2fnet22 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp11 i33#2fnet045 qf2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp10 mq2 ckb i33#2fnet047 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp9 i33#2fnet047 mq_x2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp8 mq_x2 mq2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp7 sfbn_2 ckbb i33#2fnet045 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp6 qf2 sfbn_2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp4 mq2 ckbb i33#2fnet027 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp3 sfbn_2 ckb mq_x2 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi33#2fp1 i33#2fnet027 net020 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fp1 q2 sfbn_2 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi31#2fp1 q1 sfbn_1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi30#2fp11 i30#2fnet045 qf1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp10 mq1 ckb i30#2fnet047 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp9 i30#2fnet047 mq_x1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp8 mq_x1 mq1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp7 sfbn_1 ckbb i30#2fnet045 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp6 qf1 sfbn_1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp4 mq1 ckbb i30#2fnet027 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp3 sfbn_1 ckb mq_x1 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi30#2fp1 i30#2fnet027 net019 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fp15 i29#2fseb se vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fp12 i29#2fnd_out d1 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fp2 i29#2fnd_out rd vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fp1 net019 se i29#2fnd_out vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fp0 i29#2fnet22 qf0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi29#2fn1 net019 i29#2fseb i29#2fnet22 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fp1 q0 sfbn vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp15 i0#2fseb se vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp12 i0#2fnd_out d0 vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp2 i0#2fnd_out rd vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp1 net050 se i0#2fnd_out vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp0 i0#2fnet22 si vdd vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn1 net050 i0#2fseb i0#2fnet22 vdd p08_rev3 l=0.014u nf=1 m=1 nfin=2   
.ends SAEDRVT14_FSDPSYNRBQM4_V2Y2_1




.subckt SAEDRVT14_FSDPSYNRBQ_V2_0P5 vdd vss vbp vbn q ck d si se rd
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnd_out rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 net050 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet23 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnd_out d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnd_out i0#2fseb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V2_0P5




.subckt SAEDRVT14_FSDPSYNRBQ_V2_1 vdd vss vbp vbn q ck d si se rd
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnd_out rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 net050 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet23 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnd_out d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnd_out i0#2fseb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V2_1




.subckt SAEDRVT14_FSDPSYNRBQ_V2_2 vdd vss vbp vbn q ck d si se rd
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnd_out rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 net050 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet23 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnd_out d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnd_out i0#2fseb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V2_2




.subckt SAEDRVT14_FSDPSYNRBQ_V2_4 vdd vss vbp vbn q ck d si se rd
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnd_out rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 net050 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet030 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet23 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnd_out d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnd_out i0#2fseb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V2_4




.subckt SAEDRVT14_FSDPSYNRBQ_V2LP_0P5 vdd vss vbp vbn q ck d si se rd
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 net050 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnd_out rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet23 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnd_out d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnd_out i0#2fseb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V2LP_0P5




.subckt SAEDRVT14_FSDPSYNRBQ_V2LP_1 vdd vss vbp vbn q ck d si se rd
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 net050 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnd_out rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet23 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnd_out d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnd_out i0#2fseb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V2LP_1




.subckt SAEDRVT14_FSDPSYNRBQ_V2LP_2 vdd vss vbp vbn q ck d si se rd
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 net050 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnd_out rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet23 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnd_out d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnd_out i0#2fseb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V2LP_2




.subckt SAEDRVT14_FSDPSYNRBQ_V3_1 vdd vss vbp vbn q ck d si se rd
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp14 qf_x ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnd_out rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net049 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 net049 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn17 qf_x ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet23 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn4 i0#2fnd_out d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn3 i0#2fnd_out i0#2fseb net049 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net049 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V3_1




.subckt SAEDRVT14_FSDPSYNRBQ_V3_2 vdd vss vbp vbn q ck d si se rd
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp14 qf_x ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnd_out rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net049 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 net049 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf_x ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet23 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn4 i0#2fnd_out d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn3 i0#2fnd_out i0#2fseb net049 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net049 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V3_2




.subckt SAEDRVT14_FSDPSYNRBQ_V3_4 ck d q rd se si vbn vbp vdd vss
xmibase#2fsltp1 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp15 ibase#2fnet27 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp14 qf_x ckbb ibase#2fnet27 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp12 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp5 ibase#2fnet41 ckbb vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmibase#2fmp20 ibase#2fnet30 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp19 mq ckb ibase#2fnet30 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmp18 mq_x mq vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fmp17 mq net049 ibase#2fnet41 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fp0 ckb ck vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnd_out rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net049 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 net049 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fsltn1 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fn17 qf_x ckb ibase#2fnet28 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn16 ibase#2fnet28 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn14 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn7 mq net049 ibase#2fnet31 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fmn20 mq ckbb ibase#2fnet29 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn19 ibase#2fnet29 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fmn18 mq_x mq vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmibase#2fmn17 ibase#2fnet31 ckb vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn1 ckbb ckb vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi1#2fn0 ckb ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnet23 rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn4 i0#2fnd_out d i0#2fnet23 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn3 i0#2fnd_out i0#2fseb net049 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net049 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V3_4




.subckt SAEDRVT14_FSDPSYNRBQ_V2_0P5 vdd vss vbp vbn q ck d si se sd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn15 i0#2fsnb sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnd_out i0#2fsnb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnd_out d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnd_out i0#2fseb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp13 i0#2fsnb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d i0#2fnet024 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet024 i0#2fsnb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 net050 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V2_0P5




.subckt SAEDRVT14_FSDPSYNRBQ_V2_1 vdd vss vbp vbn q ck d si se sd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn15 i0#2fsnb sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnd_out i0#2fsnb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnd_out d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnd_out i0#2fseb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp13 i0#2fsnb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d i0#2fnet024 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet024 i0#2fsnb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 net050 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V2_1




.subckt SAEDRVT14_FSDPSYNRBQ_V2_2 vdd vss vbp vbn q ck d si se sd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn15 i0#2fsnb sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnd_out i0#2fsnb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnd_out d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnd_out i0#2fseb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp13 i0#2fsnb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d i0#2fnet024 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet024 i0#2fsnb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 net050 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V2_2




.subckt SAEDRVT14_FSDPSYNRBQ_V2_4 vdd vss vbp vbn q ck d si se sd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet030 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn0 ibase#2fnet030 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn15 i0#2fsnb sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnd_out i0#2fsnb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnd_out d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnd_out i0#2fseb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet029 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmibase#2fp1 ibase#2fnet029 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp13 i0#2fsnb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d i0#2fnet024 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet024 i0#2fsnb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 net050 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V2_4




.subckt SAEDRVT14_FSDPSYNRBQ_V2LP_0P5 vdd vss vbp vbn q ck d si se sd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn15 i0#2fsnb sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnd_out i0#2fsnb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnd_out d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnd_out i0#2fseb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp13 i0#2fsnb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d i0#2fnet024 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 net050 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet024 i0#2fsnb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V2LP_0P5




.subckt SAEDRVT14_FSDPSYNRBQ_V2LP_1 vdd vss vbp vbn q ck d si se sd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn15 i0#2fsnb sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnd_out i0#2fsnb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnd_out d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnd_out i0#2fseb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp13 i0#2fsnb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d i0#2fnet024 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 net050 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet024 i0#2fsnb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V2LP_1




.subckt SAEDRVT14_FSDPSYNRBQ_V2LP_2 vdd vss vbp vbn q ck d si se sd
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq_x mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf_x ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq ckb ibase#2fnet028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq_x ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn0 ibase#2fnet028 net050 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn15 i0#2fsnb sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn14 i0#2fnd_out i0#2fsnb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnd_out d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnd_out i0#2fseb net050 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet21 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 net050 se i0#2fnet21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq_x mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf_x ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq ckbb ibase#2fnet027 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf_x ckb mq_x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp1 ibase#2fnet027 net050 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp13 i0#2fsnb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fnd_out d i0#2fnet024 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 net050 i0#2fseb i0#2fnet22 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet024 i0#2fsnb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 net050 se i0#2fnd_out vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet22 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDPSYNRBQ_V2LP_2




.subckt SAEDRVT14_FSDP_V2_0P5 vdd vss vbp vbn q qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net14 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net14 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net14 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net25 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net25 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net25 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDP_V2_0P5




.subckt SAEDRVT14_FSDP_V2_1 vdd vss vbp vbn q qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net14 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net14 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net14 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net25 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net25 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net25 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDP_V2_1




.subckt SAEDRVT14_FSDP_V2_2 vdd vss vbp vbn q qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net017 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net017 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net017 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net019 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net019 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net019 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDP_V2_2




.subckt SAEDRVT14_FSDP_V2_4 vdd vss vbp vbn q qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fn6 mq_x ckb net017 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn3 net017 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 net017 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net019 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp3 net019 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 net019 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_FSDP_V2_4




.subckt SAEDRVT14_FSDP_V2LP_0P5 vdd vss vbp vbn q qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net14 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net14 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net14 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net25 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net25 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net25 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDP_V2LP_0P5




.subckt SAEDRVT14_FSDP_V2LP_1 vdd vss vbp vbn q qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net14 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net14 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net14 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net25 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net25 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net25 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDP_V2LP_1




.subckt SAEDRVT14_FSDP_V2LP_2 vdd vss vbp vbn q qn ck d si se
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn13 ibase#2fnet046 qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn12 mq_x ckbb ibase#2fnet048 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn11 ibase#2fnet048 mq vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn10 mq mq_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn9 qf ckb ibase#2fnet046 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn8 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fn6 mq_x ckb net017 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fn5 mq ckbb qf vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi3#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fn0 qn qf vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn17 i0#2fseb se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn3 net017 d i0#2fnet22 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn2 i0#2fnet22 i0#2fseb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn1 net017 se i0#2fnet19 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmn0 i0#2fnet19 si vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb ck vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp11 ibase#2fnet045 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp10 mq_x ckb ibase#2fnet047 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp9 ibase#2fnet047 mq vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp8 mq mq_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp7 qf ckbb ibase#2fnet045 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp6 qf_x qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmibase#2fp4 mq_x ckbb net019 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmibase#2fp3 qf ckb mq vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi3#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fp1 qn qf vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp15 i0#2fseb se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp3 net019 d i0#2fnet21 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp2 i0#2fnet21 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 net019 i0#2fseb i0#2fnet20 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0 i0#2fnet20 si vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_FSDP_V2LP_2




.subckt SAEDRVT14_INV_0P5 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 x a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_INV_0P5




.subckt SAEDRVT14_INV_0P75 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_INV_0P75




.subckt SAEDRVT14_INV_10 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=10 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=10 m=1 nfin=4
.ends SAEDRVT14_INV_10




.subckt SAEDRVT14_INV_12 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=12 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=12 m=1 nfin=4
.ends SAEDRVT14_INV_12




.subckt SAEDRVT14_INV_16 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=16 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=16 m=1 nfin=4
.ends SAEDRVT14_INV_16




.subckt SAEDRVT14_INV_1P5 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_INV_1P5




.subckt SAEDRVT14_INV_1 vdd vss vbp vbn x a
xmmn0 x a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 x a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_INV_1




.subckt SAEDRVT14_INV_20 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=20 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=20 m=1 nfin=4
.ends SAEDRVT14_INV_20




.subckt SAEDRVT14_INV_2 vdd vss vbp vbn x a
xmmn0 x a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmp0 x a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_INV_2




.subckt SAEDRVT14_INV_3 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmp1 x a vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
.ends SAEDRVT14_INV_3




.subckt SAEDRVT14_INV_4 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_INV_4




.subckt SAEDRVT14_INV_6 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
.ends SAEDRVT14_INV_6




.subckt SAEDRVT14_INV_8 vdd vss vbp vbn x a
xmmn0 x a vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmmp0 x a vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
.ends SAEDRVT14_INV_8




.subckt SAEDRVT14_INV_ECO_1 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_INV_ECO_1




.subckt SAEDRVT14_INV_ECO_2 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_INV_ECO_2




.subckt SAEDRVT14_INV_ECO_3 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_INV_ECO_3




.subckt SAEDRVT14_INV_ECO_4 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_INV_ECO_4




.subckt SAEDRVT14_INV_ECO_6 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
.ends SAEDRVT14_INV_ECO_6




.subckt SAEDRVT14_INV_ECO_8 vdd vss vbp vbn x a
xmn0 x a vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
.ends SAEDRVT14_INV_ECO_8




.subckt SAEDRVT14_INV_OR2_AN2_1 a a1 a2 vbn vbp vdd vss x
xmp1 x a vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=4
xm20 x int_zn vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=2
xm19 int_zn a1 i0#2fmidp_a_b vbp p08_lvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fp0 i0#2fint_zn a2 vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fp1 i0#2fint_zn a1 vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fp2 x i0#2fint_zn vdd vbp p08_lvt l=0.014u nf=1 m=1 nfin=4
xmn0 x a vss vbn n08_lvt l=0.014u nf=1 m=1 nfin=4
xm17 int_zn a1 vss vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xm18 x int_zn vss vbn n08_lvt l=0.014u nf=1 m=1 nfin=4
xmi0#2fn3 int_zn a2 vss vbn n08_lvt l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fint_zn a1 i0#2fmidn_a_b vbn n08_lvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fn1 i0#2fmidn_a_b a2 vss vbn n08_lvt l=0.014u nf=1 m=1 nfin=3
xmi0#2fn2 x i0#2fint_zn vss vbn n08_lvt l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_INV_OR2_AN2_1




.subckt SAEDRVT14_INV_OR2_AN2_2 a a1 a2 vbn vbp vdd vss x
xm6 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi0#2fn1 i0#2fmidn_a_b a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xm5 i0#2fint_zn a1 i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn3 int_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn0 int_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn0 x a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xm8 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xm7 i0#2fint_zn a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0 i0#2fint_zn a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp2 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp1 int_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmmp0 x a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_INV_OR2_AN2_2




.subckt SAEDRVT14_INV_PECO_12 vdd vss vddr vbp vbn x a
xn1 x a vss vbn n08_rev2 l=0.014u nf=12 m=1 nfin=4
xp1 x a vddr vbp p08_rev2 l=0.014u nf=12 m=1 nfin=4
.ends SAEDRVT14_INV_PECO_12




.subckt SAEDRVT14_INV_PECO_1 vdd vss vddr vbp vbn x a
xn1 x a vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn1 net10 net10 net10 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xp1 x a vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp1 net10 net10 net10 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_INV_PECO_1




.subckt SAEDRVT14_INV_PECO_2 vdd vss vddr vbp vbn x a
xn1 x a vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xp1 x a vddr vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_INV_PECO_2




.subckt SAEDRVT14_INV_PECO_4 vdd vss vddr vbp vbn x a
xn1 x a vss vbn n08_rev2 l=0.014u nf=4 m=1 nfin=4
xp1 x a vddr vbp p08_rev2 l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_INV_PECO_4




.subckt SAEDRVT14_INV_PECO_8 vdd vss vddr vbp vbn x a
xn1 x a vss vbn n08_rev2 l=0.014u nf=8 m=1 nfin=4
xp1 x a vddr vbp p08_rev2 l=0.014u nf=8 m=1 nfin=4
.ends SAEDRVT14_INV_PECO_8




.subckt SAEDRVT14_INV_PS_1 vdd vss vddr x a
xn1 x a vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 x a vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_INV_PS_1




.subckt SAEDRVT14_INV_PS_2 vdd vss vddr x a
xn1 x a vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xp1 x a vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_INV_PS_2




.subckt SAEDRVT14_INV_PS_3 vdd vss vddr x a
xn1 x a vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xp1 x a vddr vddr p08_rev2 l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_INV_PS_3




.subckt SAEDRVT14_INV_PS_6 vdd vss vddr x a
xn1 x a vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xp1 x a vddr vddr p08_rev2 l=0.014u nf=6 m=1 nfin=4
.ends SAEDRVT14_INV_PS_6




.subckt SAEDRVT14_INV_S_0P5 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 x a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_INV_S_0P5




.subckt SAEDRVT14_INV_S_0P75 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_INV_S_0P75




.subckt SAEDRVT14_LDNQOR2_2 vdd vss vbp vbn q g ten en
xmn22 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn18 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi35#2fn23 i35#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn20 nmosdb ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi35#2fn12 qf_x ckbb i35#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi35#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn1 nmosdb en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn0 nmosdb ten vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp16 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi35#2fp21 qf_x ckb i35#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp18 qf_x ckbb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp9 i35#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp1 pmosdb ten i34#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp0 i34#2fmidp_a_b en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDNQOR2_2




.subckt SAEDRVT14_INV_S_12 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=12 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=12 m=1 nfin=4
.ends SAEDRVT14_INV_S_12




.subckt SAEDRVT14_INV_S_16 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=16 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=16 m=1 nfin=4
.ends SAEDRVT14_INV_S_16




.subckt SAEDRVT14_INV_S_1P5 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmp1 x a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_INV_S_1P5




.subckt SAEDRVT14_INV_S_1 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_INV_S_1




.subckt SAEDRVT14_INV_S_20 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=20 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=20 m=1 nfin=4
.ends SAEDRVT14_INV_S_20




.subckt SAEDRVT14_INV_S_2 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_INV_S_2




.subckt SAEDRVT14_INV_S_3 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_INV_S_3



.subckt SAEDRVT14_INV_S_4 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_INV_S_4




.subckt SAEDRVT14_INV_S_5 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=4
.ends SAEDRVT14_INV_S_5




.subckt SAEDRVT14_INV_S_6 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
.ends SAEDRVT14_INV_S_6




.subckt SAEDRVT14_INV_S_7 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=7 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=7 m=1 nfin=4
.ends SAEDRVT14_INV_S_7




.subckt SAEDRVT14_INV_S_8 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
.ends SAEDRVT14_INV_S_8




.subckt SAEDRVT14_INV_S_9 vdd vss vbp vbn x a
xmn1 x a vss vbn n08_rev l=0.014u nf=9 m=1 nfin=4
xmp1 x a vdd vbp p08_rev l=0.014u nf=9 m=1 nfin=4
.ends SAEDRVT14_INV_S_9




.subckt SAEDRVT14_ISOFSDPQ_PECO_4 vdd vss vddr q ck d si se ison
xn13 net80 qf vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn12 mq ckbb net82 vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn11 net82 mq_x vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn10 mq_x mq vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn9 qf_x ckb net80 vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn8 qf qf_x vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn6 mq ckb net83 vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn5 mq_x ckbb qf_x vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net44 net39 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn1 midn_en_ck ison vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 net39 si midn_en_ck vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn17_merged net85 sen_iso net85 vss n08_rev l=0.0140u nf=2 m=1 nfin=4
xmn21 vss net87 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn20 mq_x ckbb mq_x vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn16 net_052 net_052 net_052 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn15 mq mq mq vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn14 net55 net55 net55 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn13 net_068 net_068 net_068 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn10 sen_iso seb vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn9 seb se net054 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn8 net054 ison vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn7 ckbb ckb vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn6 ckb ck vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 q qf_x vss vss n08_rev l=0.014u nf=4 m=1 nfin=4
xmn4 net83 net55 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 net55 seb net85 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 net85 d vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 net55 sen_iso net88 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 net88 net44 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp11 net79 qf vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp10 mq ckb net81 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp9 net81 mq_x vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp8 mq_x mq vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp7 qf_x ckbb net79 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp6 qf qf_x vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 mq ckbb net84 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 qf_x ckb mq_x vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net44 net39 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 net39 si vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp0 net39 ison vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp17_merged net86 sen_iso net86 vddr p08_rev l=0.0140u nf=2 m=1 nfin=4
xmp21 net87 net87 net87 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp20 qf_x ckbb qf_x vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp16 net_052 net_052 net_052 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp15 mq mq mq vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp14 net55 net55 net55 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp13 net_068 net_068 net_068 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp10 sen_iso seb vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp9 seb ison vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp8 seb se vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp7 ckbb ckb vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp6 ckb ck vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp5 q qf_x vddr vddr p08_rev l=0.014u nf=4 m=1 nfin=4
xmp4 net84 net55 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 net55 sen_iso net86 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 net86 d vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 net55 seb net87 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 net87 net44 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ISOFSDPQ_PECO_4




.subckt SAEDRVT14_ISOFSDPQ_PECO_8 vdd vss vddr q ck d si se ison
xn13 net80 qf vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn12 mq ckbb net82 vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn11 net82 mq_x vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn10 mq_x mq vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn9 qf_x ckb net80 vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn8 qf qf_x vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn6 mq ckb net83 vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn5 mq_x ckbb qf_x vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net44 net39 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn1 midn_en_ck ison vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 net39 si midn_en_ck vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn17_merged net85 sen_iso net85 vss n08_rev l=0.0140u nf=2 m=1 nfin=4
xmn21 vss net87 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn20 mq_x ckbb mq_x vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn16 net_057 net_057 net_057 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn15 mq mq mq vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn14 net55 net55 net55 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn13 net_068 net_068 net_068 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn10 sen_iso seb vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn9 seb se net054 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn8 net054 ison vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn7 ckbb ckb vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn6 ckb ck vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 q qf_x vss vss n08_rev l=0.014u nf=8 m=1 nfin=4
xmn4 net83 net55 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 net55 seb net85 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 net85 d vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 net55 sen_iso net88 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 net88 net44 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp11 net79 qf vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp10 mq ckb net81 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp9 net81 mq_x vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp8 mq_x mq vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp7 qf_x ckbb net79 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp6 qf qf_x vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 mq ckbb net84 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 qf_x ckb mq_x vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net44 net39 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 net39 si vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp0 net39 ison vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp17_merged net86 sen_iso net86 vddr p08_rev l=0.0140u nf=2 m=1 nfin=4
xmp21 net87 net87 net87 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp20 qf_x ckbb qf_x vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp16 net_057 net_057 net_057 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp15 mq mq mq vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp14 net55 net55 net55 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp13 net_068 net_068 net_068 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp10 sen_iso seb vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp9 seb ison vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp8 seb se vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp7 ckbb ckb vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp6 ckb ck vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp5 q qf_x vddr vddr p08_rev l=0.014u nf=8 m=1 nfin=4
xmp4 net84 net55 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 net55 sen_iso net86 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 net86 d vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 net55 seb net87 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 net87 net44 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ISOFSDPQ_PECO_8




.subckt SAEDRVT14_ISOS0CL1_P_2 a en0 vbn vbp vdd vddr vss x
xn3 int_zn en0 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=2
xn0 int_zn a vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xp3 midp_a_b en0 vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp2 x int_zn vddr vbp p08_rev2 l=0.014u nf=2 m=1 nfin=2
xp1 int_zn a midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ISOS0CL1_P_2




.subckt SAEDRVT14_ISOS0CL1_P_8 a en0 vbn vbp vdd vddr vss x
xn3 int_zn en0 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn0 int_zn a vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 midp_a_b en0 vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x int_zn vddr vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp1 int_zn a midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ISOS0CL1_P_8




.subckt SAEDRVT14_ISOS0CL1_PECO_1 a en0 vbn vbp vdd vddr vss x
xn3 int_zn en0 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 int_zn a vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xmn4 vss int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xp3 midp_a_b en0 vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x int_zn vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 int_zn a midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xmp4 vddr int_zn vddr vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ISOS0CL1_PECO_1




.subckt SAEDRVT14_ISOS0CL1_PECO_2 a en0 vbn vbp vdd vddr vss x
xn3 int_zn en0 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=2
xn0 int_zn a vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 midp_a_b en0 vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x int_zn vddr vbp p08_rev2 l=0.014u nf=2 m=1 nfin=2
xp1 int_zn a midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ISOS0CL1_PECO_2




.subckt SAEDRVT14_ISOS0CL1_PECO4_1 vdd vss vddr x1 x2 x3 x4 a1 a2 a3 a4 en0
xn3 int_zn_1 en0 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net4 int_zn_1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 int_zn_1 a1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 vss int_zn_1 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x2 int_zn_2_2 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 int_zn_2_2 net5 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm3_1 net5 int_zn_2 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm2_1 int_zn_2 a2 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm11_1 net3 int_zn_3 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm10_1 int_zn_3 a3 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm20 int_zn_4 en0 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm19 net6 int_zn_4 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm18 int_zn_4 a4 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm16 vss int_zn_4 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm12 int_zn_3 en0 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm11 x4 int_zn_4_4 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm10 int_zn_4_4 net6 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm8 vss int_zn_3 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm7 x3 int_zn_3_3 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm6 int_zn_3_3 net3 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm4 int_zn_2 en0 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm3 x1 int_zn_1_1 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm2 int_zn_1_1 net4 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 vss int_zn_2 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp3 midp_a_b_1 en0 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net4 int_zn_1 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 int_zn_1 a1 midp_a_b_1 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 vddr int_zn_1 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x2 int_zn_2_2 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 int_zn_2_2 net5 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm9_1 vddr int_zn_3 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm8_1 int_zn_3_3 net3 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm7_1 midp_a_b_2 en0 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm6_1 net5 int_zn_2 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm5_1 int_zn_2 a2 midp_a_b_2 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm4_1 int_zn_1_1 net4 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm13_1 int_zn_3 a3 midp_a_b_3 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm12_1 int_zn_4_4 net6 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm23 midp_a_b_4 en0 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm22 net6 int_zn_4 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm21 int_zn_4 a4 midp_a_b_4 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm17 vddr int_zn_4 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm15 midp_a_b_3 en0 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm14 net3 int_zn_3 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm13 x4 int_zn_4_4 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm9 x3 int_zn_3_3 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 x1 int_zn_1_1 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm1 vddr int_zn_2 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ISOS0CL1_PECO4_1




.subckt SAEDRVT14_ISOS0CL1_PECO4_2 vdd vss vddr en0 a1 a2 a3 a4 x1 x2 x3 x4
xm18 int_zn_4 en0 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm17 net23 int_zn_4 vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm16 int_zn_4 a4 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm31 x2 int_zn_2_2 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm26 x3 int_zn_3_3 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm36 x1 int_zn_1_1 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm10 int_zn_3 en0 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm9 net20 int_zn_3 vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm8 int_zn_3 a3 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x4 int_zn_4_4 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm25 int_zn_3_3 net20 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm2 int_zn_2 en0 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm1 net21 int_zn_2 vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm0 int_zn_2 a2 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm29 int_zn_2_2 net21 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 int_zn_4_4 net23 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xm34 int_zn_1_1 net22 vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xn3 int_zn_1 en0 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net22 int_zn_1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn0 int_zn_1 a1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xm21 midp_a_b_4 en0 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm20 net23 int_zn_4 vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xm19 int_zn_4 a4 midp_a_b_4 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 int_zn_4_4 net23 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm27 int_zn_3_3 net20 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm13 midp_a_b_3 en0 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm12 net20 int_zn_3 vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xm11 int_zn_3 a3 midp_a_b_3 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm28 x3 int_zn_3_3 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm32 int_zn_2_2 net21 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm35 int_zn_1_1 net22 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm5 midp_a_b_2 en0 vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm4 net21 int_zn_2 vddr vddr p08_rev l=0.014u nf=2 m=1 nfin=4
xm3 int_zn_2 a2 midp_a_b_2 vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xm30 x2 int_zn_2_2 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xm33 x1 int_zn_1_1 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 x4 int_zn_4_4 vdd vddr p08_rev l=0.014u nf=1 m=1 nfin=2
xp3 midp_a_b_1 en0 vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net22 int_zn_1 vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp1 int_zn_1 a1 midp_a_b_1 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ISOS0CL1_PECO4_2




.subckt SAEDRVT14_ISOS0CL1_PECO_4 a en0 vbn vbp vdd vddr vss x
xn3 int_zn en0 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=3
xn0 int_zn a vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 midp_a_b en0 vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x int_zn vddr vbp p08_rev2 l=0.014u nf=2 m=1 nfin=3
xp1 int_zn a midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ISOS0CL1_PECO_4




.subckt SAEDRVT14_ISOS0CL1_PECO_8 a en0 vbn vbp vdd vddr vss x
xn3 int_zn en0 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn0 int_zn a vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 midp_a_b en0 vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x int_zn vddr vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp1 int_zn a midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ISOS0CL1_PECO_8




.subckt SAEDRVT14_ISOS1CL0_P_2 a en vbn vbp vdd vddr vss x
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=3
xn1 midn_en_ck en vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 int_zn a midn_en_ck vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xp2 x int_zn vddr vbp p08_rev2 l=0.014u nf=2 m=1 nfin=3
xp1 int_zn a vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 int_zn en vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ISOS1CL0_P_2




.subckt SAEDRVT14_ISOS1CL0_P_8 a en vbn vbp vdd vddr vss x
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn1 midn_en_ck en vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 int_zn a midn_en_ck vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp2 x int_zn vddr vbp p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp1 int_zn a vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 int_zn en vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ISOS1CL0_P_2




.subckt SAEDRVT14_ISOS1CL0_PECO_1 a en vbn vbp vdd vddr vss x
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn1 midn_en_ck en vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 int_zn a midn_en_ck vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xmn4 vss int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xp2 x int_zn vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp1 int_zn a vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 int_zn en vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xmp4 vddr int_zn vddr vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ISOS1CL0_PECO_1




.subckt SAEDRVT14_ISOS1CL0_PECO_2 a en vbn vbp vdd vddr vss x
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=2
xn1 midn_en_ck en vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 int_zn a midn_en_ck vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp2 x int_zn vddr vbp p08_rev2 l=0.014u nf=2 m=1 nfin=2
xp1 int_zn a vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 int_zn en vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ISOS1CL0_PECO_2




.subckt SAEDRVT14_ISOS1CL0_PECO_4 a en vbn vbp vdd vddr vss x
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=3
xn1 midn_en_ck en vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 int_zn a midn_en_ck vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xp2 x int_zn vddr vbp p08_rev2 l=0.014u nf=2 m=1 nfin=3
xp1 int_zn a vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 int_zn en vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ISOS1CL0_PECO_4




.subckt SAEDRVT14_ISOS1CL0_PECO_8 a en vbn vbp vdd vddr vss x
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn1 midn_en_ck en vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 int_zn a midn_en_ck vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x int_zn vddr vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp1 int_zn a vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 int_zn en vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ISOS1CL0_PECO_8




.subckt SAEDRVT14_LDCKNR2PQ_5 vdd vss vbp vbn q g1 g2 d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 ckb g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn7 ckb g1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 qf_x ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp01 ckb g1 net131 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 ckb g1 net13 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp71 net131 g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp7 net13 g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp21 qf_x ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_LDCKNR2PQ_5




.subckt SAEDRVT14_LDND2NQ_1 vdd vss vbp vbn q g en se
xmn22 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn23 i35#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn20 net17 ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn12 qf_x ckbb i35#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn1 i34#2fmidn_a_b en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi34#2fn0 net17 se i34#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp20 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp16 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp21 qf_x ckb i35#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp18 qf_x ckbb net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp9 i35#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp1 net16 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi34#2fp0 net16 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_LDND2NQ_1




.subckt SAEDRVT14_LDND2NQ_2 vdd vss vbp vbn q g en se
xmn22 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn23 i35#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn20 net17 ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn12 qf_x ckbb i35#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn1 i34#2fmidn_a_b en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi34#2fn0 net17 se i34#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp20 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp16 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp21 qf_x ckb i35#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp18 qf_x ckbb net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp9 i35#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp1 net16 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi34#2fp0 net16 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_LDND2NQ_2




.subckt SAEDRVT14_LDND2NQ_4 vdd vss vbp vbn q g en se
xmn22 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn23 i35#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn20 net17 ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi35#2fn12 qf_x ckbb i35#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi34#2fn1 i34#2fmidn_a_b en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi34#2fn0 net17 se i34#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp20 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp16 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp21 qf_x ckb i35#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp18 qf_x ckbb net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi35#2fp9 i35#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi34#2fp1 net16 se vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi34#2fp0 net16 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_LDND2NQ_1




.subckt SAEDRVT14_LDNQ_1 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn12 qf_x ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp21 qf_x ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckbb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDNQ_1




.subckt SAEDRVT14_LDNQ_2 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn12 qf_x ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp21 qf_x ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckbb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDNQ_2




.subckt SAEDRVT14_LDNQ_3 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 qf_x ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmi1#2fp21 qf_x ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckbb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LDNQ_3




.subckt SAEDRVT14_LDNQ_4 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 qf_x ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp21 qf_x ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_LDNQ_4




.subckt SAEDRVT14_LDNQ_5 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 qf_x ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=4
xmi1#2fp21 qf_x ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckbb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LDNQ_5




.subckt SAEDRVT14_LDNQ_6 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 qf_x ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmi1#2fp21 qf_x ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckbb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LDNQ_6




.subckt SAEDRVT14_LDNQ_8 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 qf_x ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmi1#2fp21 qf_x ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckbb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_LDNQ_8




.subckt SAEDRVT14_LDNQOR2_1 vdd vss vbp vbn q g ten en
xmn22 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn18 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi35#2fn23 i35#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn20 nmosdb ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi35#2fn12 qf_x ckbb i35#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi35#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn1 nmosdb en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn0 nmosdb ten vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp16 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi35#2fp21 qf_x ckb i35#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp18 qf_x ckbb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp9 i35#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp1 pmosdb ten i34#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp0 i34#2fmidp_a_b en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDNQOR2_1




.subckt SAEDRVT14_LDNQOR2_2 vdd vss vbp vbn q g ten en
xmn22 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn18 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi35#2fn23 i35#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn20 nmosdb ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi35#2fn12 qf_x ckbb i35#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi35#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn1 nmosdb en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn0 nmosdb ten vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp16 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi35#2fp21 qf_x ckb i35#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp18 qf_x ckbb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp9 i35#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp1 pmosdb ten i34#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp0 i34#2fmidp_a_b en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDNQOR2_2




.subckt SAEDRVT14_LDNQOR2_4 vdd vss vbp vbn q g ten en
xmn22 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn18 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi35#2fn23 i35#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn20 nmosdb ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi35#2fn12 qf_x ckbb i35#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi34#2fn1 nmosdb en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi34#2fn0 nmosdb ten vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp20 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp16 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi35#2fp21 qf_x ckb i35#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp18 qf_x ckbb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi35#2fp9 i35#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi34#2fp1 pmosdb ten i34#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi34#2fp0 i34#2fmidp_a_b en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LDNQOR2_4




.subckt SAEDRVT14_LDNQ_U_0P5 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn12 qf_x ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp21 qf_x ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckbb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDNQ_U_0P5




.subckt SAEDRVT14_LDNQ_V1_1 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 qf_x ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp21 qf_x ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckbb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDNQ_V1_1




.subckt SAEDRVT14_LDNQ_V1_2 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 qf_x ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp21 qf_x ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckbb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDNQ_V1_2




.subckt SAEDRVT14_LDNQ_V1_4 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 qf_x ckbb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp21 qf_x ckb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckbb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LDNQ_V1_4




.subckt SAEDRVT14_LDNR2PQ_1 en g q se vbn vbp vdd vss
xmp20 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp16 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp21 qf_x ckb i35#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp18 qf_x ckbb net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp9 i35#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp1 net16 se i34#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp0 i34#2fmidp_a_b en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn22 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn23 i35#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn20 net17 ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn12 qf_x ckbb i35#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn1 net17 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn0 net17 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDNR2PQ_1




.subckt SAEDRVT14_LDNR2PQ_2 en g q se vbn vbp vdd vss
xmn22 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn23 i35#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn20 net17 ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn12 qf_x ckbb i35#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn1 net17 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn0 net17 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp16 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp21 qf_x ckb i35#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp18 qf_x ckbb net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp9 i35#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp1 net16 se i34#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp0 i34#2fmidp_a_b en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDNR2PQ_2




.subckt SAEDRVT14_LDNR2PQ_4 en g q se vbn vbp vdd vss
xmn22 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn23 i35#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn20 net17 ckb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi35#2fn12 qf_x ckbb i35#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi34#2fn1 net17 en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi34#2fn0 net17 se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp20 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp16 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp21 qf_x ckb i35#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp18 qf_x ckbb net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi35#2fp9 i35#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi34#2fp1 net16 se i34#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi34#2fp0 i34#2fmidp_a_b en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LDNR2PQ_4




.subckt SAEDRVT14_LDNRBQ_V2_0P5 vdd vss vbp vbn q g d rd
xmn29 net35 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn24 qf_x ckb net35 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn23 net32 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn14 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn12 qf_x ckbb net32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 qf rb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 rb rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn9 ckb rb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn8 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp27 net36 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 qf_x ckbb net36 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp21 qf_x ckb net33 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp14 net34 rb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp11 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp10 net33 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 rb rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 qf qf_x net34 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp9 net026 rb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp8 ckb g net026 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDNRBQ_V2_0P5




.subckt SAEDRVT14_LDNRBQ_V2_1 vdd vss vbp vbn q g d rd
xmn29 net35 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn24 qf_x ckb net35 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn23 net32 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn14 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 qf_x ckbb net32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 qf rb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 rb rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn9 ckb rb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn8 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp27 net36 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 qf_x ckbb net36 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp21 qf_x ckb net33 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp14 net34 rb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp11 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp10 net33 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 rb rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 qf qf_x net34 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp9 net026 rb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp8 ckb g net026 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDNRBQ_V2_1




.subckt SAEDRVT14_LDNRBQ_V2_2 vdd vss vbp vbn q g d rd
xmn29 net35 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn24 qf_x ckb net35 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn23 net32 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn14 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn12 qf_x ckbb net32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 qf rb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 rb rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn9 ckb rb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn8 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp27 net36 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp23 qf_x ckbb net36 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp21 qf_x ckb net33 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp14 net34 rb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp11 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp10 net33 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 rb rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 qf qf_x net34 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp9 net026 rb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp8 ckb g net026 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDNRBQ_V2_2




.subckt SAEDRVT14_LDNRBQ_V2_4 vdd vss vbp vbn q g d rd
xmn29 net35 d vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn24 qf_x ckb net35 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn23 net32 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn14 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn12 qf_x ckbb net32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 qf rb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 rb rd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn9 ckb rb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn8 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp27 net36 d vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp23 qf_x ckbb net36 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp21 qf_x ckb net33 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp14 net34 rb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp11 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp10 net33 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 rb rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 qf qf_x net34 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp9 net026 rb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp8 ckb g net026 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDNRBQ_V2_4




.subckt SAEDRVT14_LDOR2PQ_1 vdd vss vbp vbn q g en se
xmn22 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn23 i35#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn20 nmose_nr_te ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn12 qf_x ckb i35#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn1 nmose_nr_te en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn0 nmose_nr_te se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp16 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp21 qf_x ckbb i35#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp18 qf_x ckb pmose_nr_te vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp9 i35#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp1 pmose_nr_te se i34#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp0 i34#2fmidp_a_b en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDOR2PQ_1




.subckt SAEDRVT14_LDOR2PQ_2 vdd vss vbp vbn q g en se
xmn22 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn23 i35#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn20 nmose_nr_te ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn12 qf_x ckb i35#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn1 nmose_nr_te en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fn0 nmose_nr_te se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp20 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp16 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp21 qf_x ckbb i35#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp18 qf_x ckb pmose_nr_te vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp9 i35#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp1 pmose_nr_te se i34#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi34#2fp0 i34#2fmidp_a_b en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDOR2PQ_2




.subckt SAEDRVT14_LDOR2PQ_4 vdd vss vbp vbn q g en se
xmn22 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn23 i35#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn20 nmose_nr_te ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi35#2fn12 qf_x ckb i35#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi34#2fn1 nmose_nr_te en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi34#2fn0 nmose_nr_te se vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp20 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp16 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp21 qf_x ckbb i35#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp18 qf_x ckb pmose_nr_te vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi35#2fp9 i35#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi35#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi34#2fp1 pmose_nr_te se i34#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi34#2fp0 i34#2fmidp_a_b en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LDOR2PQ_4




.subckt SAEDRVT14_LDPQ_1 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn12 qf_x ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp21 qf_x ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDPQ_1




.subckt SAEDRVT14_LDPQ_2 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn12 qf_x ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp21 qf_x ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDPQ_2




.subckt SAEDRVT14_LDPQ_3 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 qf_x ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmi1#2fp21 qf_x ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LDPQ_3




.subckt SAEDRVT14_LDPQ_4 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 qf_x ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp21 qf_x ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_LDPQ_4




.subckt SAEDRVT14_LDPQ_5 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 qf_x ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=4
xmi1#2fp21 qf_x ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LDPQ_5




.subckt SAEDRVT14_LDPQ_6 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 qf_x ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmi1#2fp21 qf_x ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LDPQ_6




.subckt SAEDRVT14_LDPQ_8 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 qf_x ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmi1#2fp21 qf_x ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_LDPQ_8




.subckt SAEDRVT14_LDPQ_ECO_1 vdd vss vbp vbn q g d
xmn23 net27 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 qf_x ckb net27 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn9 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn8 net26 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn7 qf_x ckbb net26 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp21 qf_x ckbb net28 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp9 net28 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp9 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp8 qf_x ckb net25 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp7 net25 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LDPQ_ECO_1




.subckt SAEDRVT14_LDPQ_U_0P5 vdd vss vbp vbn q g d
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn12 qf_x ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp21 qf_x ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDPQ_U_0P5




.subckt SAEDRVT14_LDPQ_V1_1 d g q vbn vbp vdd vss
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 qf_x ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp21 qf_x ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDPQ_V1_1




.subckt SAEDRVT14_LDPQ_V1_2 d g q vbn vbp vdd vss
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn12 qf_x ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi1#2fp21 qf_x ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDPQ_V1_2




.subckt SAEDRVT14_LDPQ_V1_4 d g q vbn vbp vdd vss
xmp23 pmosdb d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp1 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fp21 qf_x ckbb i1#2fnet98 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp18 qf_x ckb pmosdb vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp9 i1#2fnet98 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp8 qf qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmn24 nmosdb d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi1#2fn23 i1#2fnet61 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn20 nmosdb ckbb qf_x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn12 qf_x ckb i1#2fnet61 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn10 qf qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_LDPQ_V1_4




.subckt SAEDRVT14_LDPRSQB_1 d g qn rd sd vbn vbp vdd vss
xmn29 net35 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn24 qf_x ckbb net35 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn23 net32 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn14 qn qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn13 net23 sethb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn12 qf_x ckb net32 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn10 qf rd net23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 qf qf_x net23 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 sethb sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 ckb g vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp27 net36 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 qf_x ckb net36 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp21 qf_x ckbb net33 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp15 qf sethb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp14 net34 rd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp11 qn qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp10 net33 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 sethb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 qf qf_x net34 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDPRSQB_1




.subckt SAEDRVT14_LDPSBQ_V2_0P5 d g q sd vbn vbp vdd vss
xmn29 net024 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn28 qf qf_x net56 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn27 net56 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn26 net76 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn24 qf_x ckbb net024 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn23 net60 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 ckb g net76 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn14 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn12 qf_x ckb net60 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp27 net025 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp26 qf sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp25 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp24 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 qf_x ckb net025 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp21 qf_x ckbb net105 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp16 ckb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp11 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp9 net105 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDPSBQ_V2_0P5




.subckt SAEDRVT14_LDPSBQ_V2_1 d g q sd vbn vbp vdd vss
xmn29 net024 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn28 qf qf_x net56 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn27 net56 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn26 net76 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn24 qf_x ckbb net024 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn23 net60 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 ckb g net76 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn14 q qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 qf_x ckb net60 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp27 net025 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp26 qf sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp25 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp24 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 qf_x ckb net025 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp21 qf_x ckbb net105 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp16 ckb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp11 q qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp9 net105 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDPSBQ_V2_1




.subckt SAEDRVT14_LDPSBQ_V2_2 d g q sd vbn vbp vdd vss
xmn29 net024 d vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn28 qf qf_x net56 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn27 net56 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn26 net76 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn24 qf_x ckbb net024 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn23 net60 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 ckb g net76 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn14 q qf_x vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn12 qf_x ckb net60 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp27 net025 d vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp26 qf sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp25 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp24 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 qf_x ckb net025 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp21 qf_x ckbb net105 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp16 ckb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp11 q qf_x vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp9 net105 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDPSBQ_V2_2




.subckt SAEDRVT14_LDPSBQ_V2_4 d g q sd vbn vbp vdd vss
xmn29 net024 d vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn28 qf qf_x net56 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn27 net56 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn26 net76 sd vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn24 qf_x ckbb net024 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn23 net60 qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn19 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn18 ckb g net76 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn14 q qf_x vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn12 qf_x ckb net60 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp27 net025 d vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp26 qf sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp25 qf qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp24 ckb g vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp23 qf_x ckb net025 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp21 qf_x ckbb net105 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp17 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp16 ckb sd vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp11 q qf_x vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp9 net105 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LDPSBQ_V2_4




.subckt SAEDRVT14_LSRDPQ_1 d q qn vdd vddr vss ck
xm15 net29 net31 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm17 net30 net29 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm19 net30 ckn net31 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm13 d ckp net31 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm21 net29 ckn net28 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm8 ckn ck vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm9 ckp ckn vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm23 q net28 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm25 qn q vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm27 qn ckp net28 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm16 net29 net31 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm18 net30 net29 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm20 net30 ckp net31 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm14 d ckn net31 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm22 net29 ckp net28 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm7 ckn ck vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm24 q net28 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm10 ckp ckn vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm26 qn q vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm28 qn ckn net28 vss n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LSRDPQ_1




.subckt SAEDRVT14_LSRDPQ_2 d q qn vdd vddr vss ck
xm15 net29 net31 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm17 net30 net29 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm19 net30 ckn net31 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm13 d ckp net31 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm21 net29 ckn net28 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm8 ckn ck vdd vdd p08_rev l=0.014u nf=2 m=1 nfin=4
xm9 ckp ckn vdd vdd p08_rev l=0.014u nf=2 m=1 nfin=4
xm23 q net28 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm25 qn q vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm27 qn ckp net28 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm16 net29 net31 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm18 net30 net29 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm20 net30 ckp net31 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm14 d ckn net31 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm22 net29 ckp net28 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm7 ckn ck vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm24 q net28 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm10 ckp ckn vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm26 qn q vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm28 qn ckn net28 vss n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LSRDPQ_2




.subckt SAEDRVT14_LSRDPQ4_1 d1 d2 d3 d4 q1 q2 q3 q4 qn1 qn2 qn3 qn4 vdd vddr vss ck
xm88 net123 net125 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm86 net124 net123 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm84 net124 ckn net125 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm82 d4 ckp net125 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm81 net123 ckn net122 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm77 q4 net122 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm76 qn4 q4 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm70 ckn ck vdd vdd p08_rev l=0.014u nf=4 m=1 nfin=4
xm69 ckp ckn vdd vdd p08_rev l=0.014u nf=4 m=1 nfin=4
xm67 q3 net118 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm66 qn3 q3 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm62 qn3 ckp net118 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm61 net120 ckn net121 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm59 d3 ckp net121 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm56 net120 net119 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm55 net119 net121 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm53 net119 ckn net118 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm51 q2 net114 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm50 qn2 q2 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm46 qn2 ckp net114 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm45 net116 ckn net117 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm43 d2 ckp net117 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm23 q1 net110 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm25 qn1 q1 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm27 qn1 ckp net110 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm19 net112 ckn net113 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm13 d1 ckp net113 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm21 net111 ckn net110 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm37 net116 net115 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm38 net115 net117 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm15 net111 net113 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm17 net112 net111 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm40 net115 ckn net114 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm74 qn4 ckp net122 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm87 net123 net125 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm85 net124 net123 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm83 net124 ckp net125 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm80 d4 ckn net125 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm79 net123 ckp net122 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm78 q4 net122 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm75 qn4 q4 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm72 ckn ck vss vss n08_rev l=0.014u nf=4 m=1 nfin=4
xm71 ckp ckn vss vss n08_rev l=0.014u nf=4 m=1 nfin=4
xm68 q3 net118 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm65 net120 net119 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm64 qn3 q3 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm63 net119 ckp net118 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm60 qn3 ckn net118 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm58 d3 ckn net121 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm57 net120 ckp net121 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm54 net119 net121 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm52 q2 net114 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm49 net116 net115 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm48 qn2 q2 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm47 net115 ckp net114 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm44 qn2 ckn net114 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm42 d2 ckn net117 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm41 net116 ckp net117 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm24 q1 net110 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm18 net112 net111 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm26 qn1 q1 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm22 net111 ckp net110 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm28 qn1 ckn net110 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm14 d1 ckn net113 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm20 net112 ckp net113 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm16 net111 net113 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm39 net115 net117 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm73 qn4 ckn net122 vss n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LSRDPQ4_1




.subckt SAEDRVT14_LSRDPQ4_2 d1 d2 d3 d4 q1 q2 q3 q4 qn1 qn2 qn3 qn4 vdd vddr vss ck
xm76 net114 net116 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm74 net115 net114 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm72 net115 ckn net116 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm70 d4 ckp net116 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm69 net114 ckn net113 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm65 q4 net113 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm64 qn4 q4 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm62 qn4 ckp net113 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm60 net110 net112 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm58 net111 net110 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm56 net111 ckn net112 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm54 d3 ckp net112 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm53 net110 ckn net109 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm49 qn3 q3 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm48 q3 net109 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm46 qn3 ckp net109 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm44 net106 net108 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm42 net107 net106 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm40 net107 ckn net108 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm38 d2 ckp net108 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm37 net106 ckn net105 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm15 net102 net104 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm32 qn2 q2 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm33 q2 net105 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm25 qn1 q1 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm23 q1 net101 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm27 qn1 ckp net101 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm30 qn2 ckp net105 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm19 net103 ckn net104 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm8 ckn ck vdd vdd p08_rev l=0.014u nf=8 m=1 nfin=4
xm17 net103 net102 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm21 net102 ckn net101 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm13 d1 ckp net104 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm9 ckp ckn vdd vdd p08_rev l=0.014u nf=8 m=1 nfin=4
xm75 net114 net116 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm73 net115 net114 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm71 net115 ckp net116 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm68 d4 ckn net116 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm67 net114 ckp net113 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm66 q4 net113 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm63 qn4 q4 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm61 qn4 ckn net113 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm59 net110 net112 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm57 net111 net110 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm55 net111 ckp net112 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm52 d3 ckn net112 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm51 net110 ckp net109 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm50 q3 net109 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm47 qn3 ckn net109 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm45 qn3 q3 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm43 net106 net108 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm41 net107 net106 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm39 net107 ckp net108 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm36 d2 ckn net108 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm35 net106 ckp net105 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm34 q2 net105 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm26 qn1 q1 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm28 qn1 ckn net101 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm29 qn2 ckn net105 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm7 ckn ck vss vss n08_rev l=0.014u nf=8 m=1 nfin=4
xm10 ckp ckn vss vss n08_rev l=0.014u nf=8 m=1 nfin=4
xm18 net103 net102 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm22 net102 ckp net101 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm14 d1 ckn net104 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm24 q1 net101 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm16 net102 net104 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm20 net103 ckp net104 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm31 qn2 q2 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LSRDPQ4_2




.subckt SAEDRVT14_LVLDBUFE0_IY2_10 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=2
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2_10




.subckt SAEDRVT14_LVLDBUFE0_IY2_12 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=2
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2_12




.subckt SAEDRVT14_LVLDBUFE0_IY2_1 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2_1




.subckt SAEDRVT14_LVLDBUFE0_IY2_2 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2_2




.subckt SAEDRVT14_LVLDBUFE0_IY2_3 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2_3




.subckt SAEDRVT14_LVLDBUFE0_IY2_4 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2_4




.subckt SAEDRVT14_LVLDBUFE0_IY2_6 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=2 m=1 nfin=2
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLDBUFE0_IY2_6




.subckt SAEDRVT14_LVLDBUFE0_IY2_8 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=2 m=1 nfin=2
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2_8




.subckt SAEDRVT14_LVLDBUFE0_IY2V1_10 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=3
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=3
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2V1_10




.subckt SAEDRVT14_LVLDBUFE0_IY2V1_12 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=3
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=3
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2V1_12




.subckt SAEDRVT14_LVLDBUFE0_IY2V1_1 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2V1_1




.subckt SAEDRVT14_LVLDBUFE0_IY2V1_2 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2V1_2




.subckt SAEDRVT14_LVLDBUFE0_IY2V1_3 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2V1_3




.subckt SAEDRVT14_LVLDBUFE0_IY2V1_4 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2V1_4




.subckt SAEDRVT14_LVLDBUFE0_IY2V1_6 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=3
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2V1_6




.subckt SAEDRVT14_LVLDBUFE0_IY2V1_8 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=3
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 vddl vddl p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY2V1_3




.subckt SAEDRVT14_LVLDBUFE1_IY2_10 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLDBUFE1_IY2_10




.subckt SAEDRVT14_LVLDBUFE1_IY2_12 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLDBUFE1_IY2_12




.subckt SAEDRVT14_LVLDBUFE1_IY2_1 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE1_IY2_1




.subckt SAEDRVT14_LVLDBUFE1_IY2_2 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=3
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE1_IY2_2




.subckt SAEDRVT14_LVLDBUFE1_IY2_3 vddi vss vdd x a en
xn5 x net16 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddi vddi p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp4 net16 net1 net_025 vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddi vddi p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddi p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddi p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vdd vdd p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddi vddi p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE1_IY2_3




.subckt SAEDRVT14_LVLDBUFE1_IY2_4 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE1_IY2_4




.subckt SAEDRVT14_LVLDBUFE1_IY2_6 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE1_IY2_6




.subckt SAEDRVT14_LVLDBUFE1_IY2_8 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_LVLDBUFE1_IY2_8




.subckt SAEDRVT14_LVLDBUFE1_IY2V1_10 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLDBUFE1_IY2V1_10




.subckt SAEDRVT14_LVLDBUFE1_IY2V1_12 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLDBUFE1_IY2V1_12




.subckt SAEDRVT14_LVLDBUFE1_IY2V1_1 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE1_IY2V1_1




.subckt SAEDRVT14_LVLDBUFE1_IY2V1_2 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=3
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE1_IY2V1_2




.subckt SAEDRVT14_LVLDBUFE1_IY2V1_3 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE1_IY2V1_3




.subckt SAEDRVT14_LVLDBUFE1_IY2V1_4 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE1_IY2V1_4




.subckt SAEDRVT14_LVLDBUFE1_IY2V1_6 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE1_IY2V1_6




.subckt SAEDRVT14_LVLDBUFE1_IY2V1_8 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddl vddl p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 net_025 vddl p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddl vddl p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_LVLDBUFE1_IY2V1_10




.subckt SAEDRVT14_LVLDBUF_IY2V1_10 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=7 m=1 nfin=4
xp4 x net14 vddl vddl p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp3 net14 net1 vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUF_IY2V1_10




.subckt SAEDRVT14_LVLDBUF_IY2V1_12 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=7 m=1 nfin=4
xp4 x net14 vddl vddl p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp3 net14 net1 vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUF_IY2V1_12




.subckt SAEDRVT14_LVLDBUF_IY2V1_1 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=5 m=1 nfin=4
xp4 x net14 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net14 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net1 net2 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUF_IY2V1_1




.subckt SAEDRVT14_LVLDBUF_IY2V1_2 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=5 m=1 nfin=4
xp4 x net14 vddl vddl p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net14 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net1 net2 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUF_IY2V1_2




.subckt SAEDRVT14_LVLDBUF_IY2V1_3 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=5 m=1 nfin=4
xp4 x net14 vddl vddl p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net14 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net1 net2 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUF_IY2V1_3




.subckt SAEDRVT14_LVLDBUF_IY2V1_4 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=5 m=1 nfin=4
xp4 x net14 vddl vddl p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp3 net14 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net1 net2 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUF_IY2V1_4




.subckt SAEDRVT14_LVLDBUF_IY2V1_6 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=7 m=1 nfin=4
xp4 x net14 vddl vddl p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp3 net14 net1 vddl vddl p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp2 net1 net2 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUF_IY2V1_6




.subckt SAEDRVT14_LVLDBUF_IY2V1_8 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=7 m=1 nfin=4
xp4 x net14 vddl vddl p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp3 net14 net1 vddl vddl p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp2 net1 net2 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUF_IY2V1_8




.subckt SAEDRVT14_LVLDBUFE0_IY_2 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLDBUFE0_IY_2



.subckt SAEDRVT14_LVLUBUF4E0_IY2_2 vss en a1 a2 a3 a4 vddh vddl x1 x2 x3 x4
xi6 vss x4 a4 en vddh vddl SAEDRVT14_LVLUBUFE0_IY2_2
xi5 vss x3 a3 en vddh vddl SAEDRVT14_LVLUBUFE0_IY2_2
xi4 vss x2 a2 en vddh vddl SAEDRVT14_LVLUBUFE0_IY2_2
xi0 vss x1 a1 en vddh vddl SAEDRVT14_LVLUBUFE0_IY2_2
.ends SAEDRVT14_LVLUBUF4E0_IY2_2




.subckt SAEDRVT14_LVLUBUFE0_IY2_4 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE0_IY2_4



.subckt SAEDRVT14_LVLUBUF4E0_IY2_4 vss en a1 a2 a3 a4 vddh vddl x1 x2 x3 x4
xi0 vss x1 a1 en vddh vddl SAEDRVT14_LVLUBUFE0_IY2_4
xi6 vss x4 a4 en vddh vddl SAEDRVT14_LVLUBUFE0_IY2_4
xi5 vss x3 a3 en vddh vddl SAEDRVT14_LVLUBUFE0_IY2_4
xi4 vss x2 a2 en vddh vddl SAEDRVT14_LVLUBUFE0_IY2_4
.ends SAEDRVT14_LVLUBUF4E0_IY2_4




.subckt SAEDRVT14_LVLUBUFE0_IY2_8 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE0_IY2_8

.subckt SAEDRVT14_LVLUBUF4E0_IY2_8 vss en a1 a2 a3 a4 vddh vddl x1 x2 x3 x4
xi0 vss x1 a1 en vddh vddl SAEDRVT14_LVLUBUFE0_IY2_8
xi6 vss x4 a4 en vddh vddl SAEDRVT14_LVLUBUFE0_IY2_8
xi5 vss x3 a3 en vddh vddl SAEDRVT14_LVLUBUFE0_IY2_8
xi4 vss x2 a2 en vddh vddl SAEDRVT14_LVLUBUFE0_IY2_8
.ends SAEDRVT14_LVLUBUF4E0_IY2_8




.subckt SAEDRVT14_LVLUBUFE0_IY2_10 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE0_IY2_10




.subckt SAEDRVT14_LVLUBUFE0_IY2_12 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp4 net16 net1 vddh vddh p08 l=0.014u nf=1
!Error: Error: Error while looking for the value of parameter "m" for the instance xp4 in the design rvt/SAEDRVT14_LVLUBUFE0_IY2_12/schematic: parse failed: "NFIN=4" char(5) (NETLISTING-017)
 nfin=1
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE0_IY2_12



.subckt SAEDRVT14_LVLUBUFE0_IY2_1 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE0_IY2_1




.subckt SAEDRVT14_LVLUBUFE0_IY2_2 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE0_IY2_2




.subckt SAEDRVT14_LVLUBUFE0_IY2_3 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE0_IY2_3




.subckt SAEDRVT14_LVLUBUFE0_IY2_4 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE0_IY2_4




.subckt SAEDRVT14_LVLUBUFE0_IY2_6 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE0_IY2_6




.subckt SAEDRVT14_LVLUBUFE0_IY2_8 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE0_IY2_8




.subckt SAEDRVT14_LVLUBUFE0_IY2V1_10 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE0_IY2V1_10




.subckt SAEDRVT14_LVLUBUFE0_IY2V1_12 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE0_IY2V1_12




.subckt SAEDRVT14_LVLUBUFE0_IY2V1_1 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE0_IY2V1_1




.subckt SAEDRVT14_LVLUBUFE0_IY2V1_2 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE0_IY2V1_2




.subckt SAEDRVT14_LVLUBUFE0_IY2V1_3 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE0_IY2V1_3




.subckt SAEDRVT14_LVLUBUFE0_IY2V1_4 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE0_IY2V1_4




.subckt SAEDRVT14_LVLUBUFE0_IY2V1_6 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE0_IY2V1_6




.subckt SAEDRVT14_LVLUBUFE0_IY2V1_8 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net1 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_fet vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=2
xn0 net8 net_fet vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_fet a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=2
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 vddh vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_fet vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp6 net_fet a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE0_IY2V1_3




.subckt SAEDRVT14_LVLUBUFE1_IY2_10 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE1_IY2_10




.subckt SAEDRVT14_LVLUBUFE1_IY2_12 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE1_IY2_12




.subckt SAEDRVT14_LVLUBUFE1_IY2_1 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE1_IY2_1




.subckt SAEDRVT14_LVLUBUFE1_IY2_2 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE1_IY2_2




.subckt SAEDRVT14_LVLUBUFE1_IY2_3 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE1_IY2_3




.subckt SAEDRVT14_LVLUBUFE1_IY2_4 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE1_IY2_4




.subckt SAEDRVT14_LVLUBUFE1_IY2_6 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE1_IY2_6




.subckt SAEDRVT14_LVLUBUFE1_IY2_8 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_LVLUBUFE1_IY2_8




.subckt SAEDRVT14_LVLUBUFE1_IY2V1_10 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE1_IY2V1_10




.subckt SAEDRVT14_LVLUBUFE1_IY2V1_12 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUFE1_IY2V1_12




.subckt SAEDRVT14_LVLUBUFE1_IY2V1_1 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_09 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_09 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_09 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_09 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_09 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE1_IY2V1_1




.subckt SAEDRVT14_LVLUBUFE1_IY2V1_2 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE1_IY2V1_2




.subckt SAEDRVT14_LVLUBUFE1_IY2V1_3 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE1_IY2V1_3




.subckt SAEDRVT14_LVLUBUFE1_IY2V1_4 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=3
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE1_IY2V1_4




.subckt SAEDRVT14_LVLUBUFE1_IY2V1_6 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUFE1_IY2V1_6




.subckt SAEDRVT14_LVLUBUFE1_IY2V1_8 vss x a en vddh vddl
xn5 x net16 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn4 net16 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net16 iso vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn6 net_08 a vss vss n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 iso en vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp5 x net16 vddh vddh p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp4 net16 net1 net_025 vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net_012 iso vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 net_012 vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp7 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 net_025 iso vddh vddh p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 iso en vddh vddh p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_LVLUBUFE1_IY2V1_8




.subckt SAEDRVT14_LVLUBUF_IY2_10 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=3
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=10 m=1 nfin=3
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUF_IY2_10




.subckt SAEDRVT14_LVLUBUF_IY2_12 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=3
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=12 m=1 nfin=3
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUF_IY2_12




.subckt SAEDRVT14_LVLUBUF_IY2_1 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUF_IY2_1




.subckt SAEDRVT14_LVLUBUF_IY2_2 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUF_IY2_2




.subckt SAEDRVT14_LVLUBUF_IY2_3 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUF_IY2_3




.subckt SAEDRVT14_LVLUBUF_IY2_4 vdd vss vddi x a
xn4 x net14 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp4 x net14 vdd vdd p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp3 net14 net1 vdd vdd p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp2 net1 net2 vdd vdd p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vdd vdd p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddi vddi p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddi vddi p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUF_IY2_4




.subckt SAEDRVT14_LVLUBUF_IY2_6 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=7 m=1 nfin=4
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUF_IY2_6




.subckt SAEDRVT14_LVLUBUF_IY2_8 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_LVLUBUF_IY2_8




.subckt SAEDRVT14_LVLUBUF_IY2V1_10 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=10 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=7 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=10 m=1 nfin=4
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUF_IY2V1_10




.subckt SAEDRVT14_LVLUBUF_IY2V1_12 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=12 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=7 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=12 m=1 nfin=4
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUF_IY2V1_12




.subckt SAEDRVT14_LVLUBUF_IY2V1_1 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=5 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUF_IY2V1_1




.subckt SAEDRVT14_LVLUBUF_IY2V1_2 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=5 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUF_IY2V1_2




.subckt SAEDRVT14_LVLUBUF_IY2V1_3 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=5 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUF_IY2V1_3




.subckt SAEDRVT14_LVLUBUF_IY2V1_4 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=5 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUF_IY2V1_4




.subckt SAEDRVT14_LVLUBUF_IY2V1_6 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=7 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUF_IY2V1_6




.subckt SAEDRVT14_LVLUBUF_IY2V1_8 vss x a vddh vddl
xn4 x net14 vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn3 net14 net1 vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 net1 net_08 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn1 net2 net8 vss vss n08_rev2 l=0.014u nf=7 m=1 nfin=4
xn0 net8 net_08 vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn4 net_08 a vss vss n08_rev l=0.014u nf=7 m=1 nfin=4
xp4 x net14 vddh vddh p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp3 net14 net1 vddh vddh p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp2 net1 net2 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net2 net1 vddh vddh p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net8 net_08 vddl vddl p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp4 net_08 a vddl vddl p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_LVLUBUF_IY2V1_8





.subckt SAEDRVT14_MUX2_1P5 d0 d1 s vbn vbp vdd vss x
xmn4 x net77 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmmn5 net09 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn4 i0#2fnet20 net09 net77 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn3 i0#2fnet18 s net77 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x net77 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmmp5 net09 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp4 i0#2fnet21 s net77 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fnet19 net09 net77 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_MUX2_1P5




.subckt SAEDRVT14_MUX2_1 d0 d1 s vbn vbp vdd vss x
xmn4 x net77 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn5 net09 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net09 net77 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnet18 s net77 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 x net77 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp5 net09 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s net77 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fnet19 net09 net77 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_MUX2_1




.subckt SAEDRVT14_MUX2_2 d0 d1 s vbn vbp vdd vss x
xmn4 x net77 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn5 net09 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net09 net77 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn3 i0#2fnet18 s net77 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x net77 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp5 net09 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s net77 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fnet19 net09 net77 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_MUX2_2




.subckt SAEDRVT14_MUX2_4 vdd vss vbp vbn x d0 d1 s
xmp4 x net77 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmmp5 net09 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp41 i0#2fnet211 s net77 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp31 i0#2fnet191 net09 net77 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp21 i0#2fnet211 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp01 i0#2fnet191 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp4 i0#2fnet21 s net77 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fnet19 net09 net77 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 x net77 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmmn5 net09 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn41 i0#2fnet201 net09 net77 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn31 i0#2fnet181 s net77 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn21 i0#2fnet201 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn01 i0#2fnet181 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn4 i0#2fnet20 net09 net77 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn3 i0#2fnet18 s net77 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_MUX2_4




.subckt SAEDRVT14_MUX2_ECO_1 vdd vss vbp vbn x d0 d1 s
xmp4 x net77 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp9 net77 sb net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp8 net015 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp7 net013 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp6 net77 s net013 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp5 sb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 x net77 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn9 net77 s net014 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn8 net014 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn7 net012 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn6 net77 sb net012 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn5 sb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_MUX2_ECO_1




.subckt SAEDRVT14_MUX2_ECO_2 vdd vss vbp vbn x d0 d1 s
xmmp11 x net9 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp10 net9 sb net19 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp9 net19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp8 sb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp7 net20 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp6 net9 s net20 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmn11 x net9 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn10 net18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn9 net9 s net18 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn8 net9 sb net21 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn7 net21 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn6 sb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_MUX2_ECO_2




.subckt SAEDRVT14_MUX2_MM_0P5 vdd vss vbp vbn x d0 d1 s
xmp4 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp5 net9 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fnet19 net9 int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn5 net9 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net9 int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnet18 s int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_MUX2_MM_0P5




.subckt SAEDRVT14_MUX2_MM_1 vdd vss vbp vbn x d0 d1 s
xmp4 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp5 net9 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fnet19 net9 int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn5 net9 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net9 int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnet18 s int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_MUX2_MM_1




.subckt SAEDRVT14_MUX2_MM_2 vdd vss vbp vbn x d0 d1 s
xmp4 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp5 net9 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp4 i0#2fnet21 s int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fnet19 net9 int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn5 net9 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn4 i0#2fnet20 net9 int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn3 i0#2fnet18 s int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_MUX2_MM_2




.subckt SAEDRVT14_MUX2_MM_4 vdd vss vbp vbn x d0 d1 s
xmp4 x int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmmp5 net9 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp41 i0#2fnet211 s int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp31 i0#2fnet191 net9 int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp21 i0#2fnet211 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp01 i0#2fnet191 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp4 i0#2fnet21 s int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fnet19 net9 int_zn vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 x int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmmn5 net9 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn41 i0#2fnet201 net9 int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn31 i0#2fnet181 s int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn21 i0#2fnet201 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn01 i0#2fnet181 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn4 i0#2fnet20 net9 int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn3 i0#2fnet18 s int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_MUX2_MM_4




.subckt SAEDRVT14_MUX2_U_0P5 vdd vss vbp vbn x d0 d1 s
xmp4 x net77 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp5 net08 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s net77 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fnet19 net08 net77 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 x net77 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn5 net08 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net08 net77 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnet18 s net77 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_MUX2_U_0P5




.subckt SAEDRVT14_MUX3_V1M_0P5 vdd vss vbp vbn x d0 d1 d2 s0 s1
xmn3 x net015 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 net017 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 net125 d2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 net016 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xi1#2fn4 net018 net017 net015 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn3 net125 s1 net015 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn4 i0#2fnet20 net016 net018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn3 i0#2fnet18 s0 net018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xmp3 x net015 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 net017 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 net125 d2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 net016 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xi1#2fp4 net018 s1 net015 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp3 net125 net017 net015 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp4 i0#2fnet21 s0 net018 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp3 i0#2fnet19 net016 net018 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
.ends SAEDRVT14_MUX3_V1M_0P5




.subckt SAEDRVT14_MUX3_V1M_1 vdd vss vbp vbn x d0 d1 d2 s0 s1
xmn3 x net015 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 net017 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 net125 d2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 net016 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xi1#2fn4 net018 net017 net015 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn3 net125 s1 net015 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn4 i0#2fnet20 net016 net018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn3 i0#2fnet18 s0 net018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xmp3 x net015 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 net017 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 net125 d2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 net016 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xi1#2fp4 net018 s1 net015 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp3 net125 net017 net015 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp4 i0#2fnet21 s0 net018 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp3 i0#2fnet19 net016 net018 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
.ends SAEDRVT14_MUX3_V1M_1




.subckt SAEDRVT14_MUX3_V1M_2 vdd vss vbp vbn x d0 d1 d2 s0 s1
xmn3 x net015 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn2 net017 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 net125 d2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 net016 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xi1#2fn4 net018 net017 net015 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn3 net125 s1 net015 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn4 i0#2fnet20 net016 net018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn3 i0#2fnet18 s0 net018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xmp3 x net015 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp2 net017 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 net125 d2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 net016 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xi1#2fp4 net018 s1 net015 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp3 net125 net017 net015 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp4 i0#2fnet21 s0 net018 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp3 i0#2fnet19 net016 net018 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
.ends SAEDRVT14_MUX3_V1M_2




.subckt SAEDRVT14_MUX3_V1M_4 vdd vss vbp vbn x d0 d1 d2 s0 s1
xmn3 x net015 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn2 net017 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 net125 d2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 net016 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xi1#2fn4 net018 net017 net015 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn3 net125 s1 net015 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn41 i0#2fnet201 net016 net018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn31 i0#2fnet181 s0 net018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn21 i0#2fnet201 d0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn01 i0#2fnet181 d1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn4 i0#2fnet20 net016 net018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn3 i0#2fnet18 s0 net018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xmp3 x net015 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp2 net017 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 net125 d2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 net016 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xi1#2fp4 net018 s1 net015 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp3 net125 net017 net015 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp41 i0#2fnet211 s0 net018 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp31 i0#2fnet191 net016 net018 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp21 i0#2fnet211 d0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp01 i0#2fnet191 d1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp4 i0#2fnet21 s0 net018 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp3 i0#2fnet19 net016 net018 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
.ends SAEDRVT14_MUX3_V1M_4




.subckt SAEDRVT14_MUX4_V1M_1 vdd vss vbp vbn x d0 d1 d2 d3 s0 s1
xmn13 net18 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn12 x net15 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn5 net12 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xi2#2fn4 net17 net18 net15 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn3 net16 s1 net15 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn4 i1#2fnet20 net12 net17 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn3 i1#2fnet18 s0 net17 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn2 i1#2fnet20 d0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn0 i1#2fnet18 d1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn4 i0#2fnet20 net12 net16 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn3 i0#2fnet18 s0 net16 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn2 i0#2fnet20 d2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn0 i0#2fnet18 d3 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xmp13 net18 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp12 x net15 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 net12 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xi2#2fp4 net17 s1 net15 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp3 net16 net18 net15 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp4 i1#2fnet21 s0 net17 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp3 i1#2fnet19 net12 net17 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp2 i1#2fnet21 d0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp0 i1#2fnet19 d1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp4 i0#2fnet21 s0 net16 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp3 i0#2fnet19 net12 net16 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp2 i0#2fnet21 d2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp0 i0#2fnet19 d3 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
.ends SAEDRVT14_MUX4_V1M_1




.subckt SAEDRVT14_MUX4_V1M_2 vdd vss vbp vbn x d0 d1 d2 d3 s0 s1
xmn13 net18 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 x net15 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 net12 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xi2#2fn4 net17 net18 net15 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn3 net16 s1 net15 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn4 i1#2fnet20 net12 net17 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn3 i1#2fnet18 s0 net17 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn2 i1#2fnet20 d0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn0 i1#2fnet18 d1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn4 i0#2fnet20 net12 net16 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn3 i0#2fnet18 s0 net16 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn2 i0#2fnet20 d2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn0 i0#2fnet18 d3 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xmp13 net18 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp12 x net15 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp5 net12 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xi2#2fp4 net17 s1 net15 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp3 net16 net18 net15 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp4 i1#2fnet21 s0 net17 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp3 i1#2fnet19 net12 net17 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp2 i1#2fnet21 d0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp0 i1#2fnet19 d1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp4 i0#2fnet21 s0 net16 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp3 i0#2fnet19 net12 net16 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp2 i0#2fnet21 d2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp0 i0#2fnet19 d3 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
.ends SAEDRVT14_MUX4_V1M_2




.subckt SAEDRVT14_MUX4_V1M_4 vdd vss vbp vbn x d0 d1 d2 d3 s0 s1
xmn13 net18 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 x net15 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn5 net12 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xi2#2fn4 net17 net18 net15 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn3 net16 s1 net15 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn41 i1#2fnet201 net12 net17 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn31 i1#2fnet181 s0 net17 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn21 i1#2fnet201 d0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn01 i1#2fnet181 d1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn4 i1#2fnet20 net12 net17 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn3 i1#2fnet18 s0 net17 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn2 i1#2fnet20 d0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn0 i1#2fnet18 d1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn41 i0#2fnet201 net12 net16 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn31 i0#2fnet181 s0 net16 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn21 i0#2fnet201 d2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn01 i0#2fnet181 d3 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn4 i0#2fnet20 net12 net16 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn3 i0#2fnet18 s0 net16 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn2 i0#2fnet20 d2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn0 i0#2fnet18 d3 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xmp13 net18 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp12 x net15 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp5 net12 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xi2#2fp4 net17 s1 net15 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp3 net16 net18 net15 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp41 i1#2fnet211 s0 net17 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp31 i1#2fnet191 net12 net17 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp21 i1#2fnet211 d0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp01 i1#2fnet191 d1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp4 i1#2fnet21 s0 net17 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp3 i1#2fnet19 net12 net17 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp2 i1#2fnet21 d0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp0 i1#2fnet19 d1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp41 i0#2fnet211 s0 net16 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp31 i0#2fnet191 net12 net16 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp21 i0#2fnet211 d2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp01 i0#2fnet191 d3 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp4 i0#2fnet21 s0 net16 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp3 i0#2fnet19 net12 net16 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp2 i0#2fnet21 d2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp0 i0#2fnet19 d3 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
.ends SAEDRVT14_MUX4_V1M_4




.subckt SAEDRVT14_MUX4_V1U_0P5 vdd vss vbp vbn x d0 d1 d2 d3 s0 s1
xmn13 net18 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn12 x net15 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn5 net12 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xi2#2fn4 net17 net18 net15 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn3 net16 s1 net15 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn4 i1#2fnet20 net12 net17 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn3 i1#2fnet18 s0 net17 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn2 i1#2fnet20 d0 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn0 i1#2fnet18 d1 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn4 i0#2fnet20 net12 net16 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn3 i0#2fnet18 s0 net16 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn2 i0#2fnet20 d2 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn0 i0#2fnet18 d3 vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xmp13 net18 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp12 x net15 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 net12 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xi2#2fp4 net17 s1 net15 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp3 net16 net18 net15 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp4 i1#2fnet21 s0 net17 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp3 i1#2fnet19 net12 net17 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp2 i1#2fnet21 d0 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp0 i1#2fnet19 d1 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp4 i0#2fnet21 s0 net16 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp3 i0#2fnet19 net12 net16 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp2 i0#2fnet21 d2 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp0 i0#2fnet19 d3 vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
.ends SAEDRVT14_MUX4_V1U_0P5




.subckt SAEDRVT14_MUXI2_0P5 vdd vss vbp vbn x d0 d1 s
xmmp7 x net029 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp6 net029 net028 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp5 net036 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s net028 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fnet19 net036 net028 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmn7 x net029 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn6 net029 net028 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn5 net036 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net036 net028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnet18 s net028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_MUXI2_0P5




.subckt SAEDRVT14_MUXI2_1 vdd vss vbp vbn x d0 d1 s
xmmp7 x net029 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp6 net029 net028 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp5 net036 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s net028 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fnet19 net036 net028 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmn7 x net029 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn6 net029 net028 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn5 net036 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net036 net028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnet18 s net028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_MUXI2_1




.subckt SAEDRVT14_MUXI2_2 vdd vss vbp vbn x d0 d1 s
xmmp7 x net029 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp6 net029 net028 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmmp5 net036 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s net028 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fnet19 net036 net028 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmn7 x net029 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn6 net029 net028 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmmn5 net036 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net036 net028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnet18 s net028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_MUXI2_2




.subckt SAEDRVT14_MUXI2_4 vdd vss vbp vbn x d0 d1 s
xmmp7 x net029 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmmp6 net029 net028 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp5 net036 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s net028 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fnet19 net036 net028 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmn7 x net029 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmmn6 net029 net028 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn5 net036 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net036 net028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnet18 s net028 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_MUXI2_4




.subckt SAEDRVT14_MUXI2_B_1 vdd vss vbp vbn x d0 d1 s
xmmp5 net036 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp4 i0#2fnet21 s x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fnet19 net036 x vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmn5 net036 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn4 i0#2fnet20 net036 x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn3 i0#2fnet18 s x vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_MUXI2_B_1




.subckt SAEDRVT14_MUXI2_ECO_1 vdd vss vbp vbn x d0 d1 s
xmmp11 net028 sb net014 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp10 net014 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp9 net028 s net013 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp8 net013 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp7 x net029 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp6 net029 net028 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp5 sb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmn11 net015 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn10 net028 s net015 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn9 net028 sb net016 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn8 net016 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn7 x net029 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn6 net029 net028 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn5 sb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_MUXI2_ECO_1




.subckt SAEDRVT14_MUXI2_ECO_2 vdd vss vbp vbn x d0 d1 s
xmmp11 net9 sb net20 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp10 net20 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp9 net9 s net19 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp8 net19 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp7 x net17 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp6 net17 net9 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp5 sb s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmn11 net22 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn10 net9 s net22 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn9 net9 sb net21 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn8 net21 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn7 x net17 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn6 net17 net9 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn5 sb s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_MUXI2_ECO_2




.subckt SAEDRVT14_MUXI2_U_0P5 vdd vss vbp vbn x d0 d1 s
xmmp5 net036 s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fnet19 net036 x vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmn5 net036 s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net036 x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnet18 s x vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_MUXI2_U_0P5




.subckt SAEDRVT14_MUXI3_0P5 vdd vss vbp vbn x d0 d1 d2 s0 s1
xmmn4 x net021 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn3 net021 net015 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn2 net017 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn1 net125 d2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn0 net016 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn4 net018 net017 net015 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn3 net125 s1 net015 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net016 net018 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnet18 s0 net018 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmp4 x net021 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp3 net021 net015 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp2 net017 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp1 net125 d2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp0 net016 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp4 net018 s1 net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp3 net125 net017 net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s0 net018 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fnet19 net016 net018 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_MUXI3_0P5




.subckt SAEDRVT14_MUXI3_1 vdd vss vbp vbn x d0 d1 d2 s0 s1
xmmn4 x net021 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn3 net021 net015 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn2 net017 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn1 net125 d2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn0 net016 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn4 net018 net017 net015 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn3 net125 s1 net015 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net016 net018 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnet18 s0 net018 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmp4 x net021 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp3 net021 net015 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp2 net017 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp1 net125 d2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp0 net016 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp4 net018 s1 net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp3 net125 net017 net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s0 net018 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fnet19 net016 net018 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_MUXI3_1




.subckt SAEDRVT14_MUXI3_2 vdd vss vbp vbn x d0 d1 d2 s0 s1
xmmn4 x net021 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn3 net021 net015 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn2 net017 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn1 net125 d2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn0 net016 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn4 net018 net017 net015 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn3 net125 s1 net015 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn4 i0#2fnet20 net016 net018 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn3 i0#2fnet18 s0 net018 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmp4 x net021 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp3 net021 net015 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp2 net017 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 net125 d2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 net016 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp4 net018 s1 net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp3 net125 net017 net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp4 i0#2fnet21 s0 net018 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fnet19 net016 net018 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_MUXI3_2




.subckt SAEDRVT14_MUXI3_4 vdd vss vbp vbn x d0 d1 d2 s0 s1
xmmn4 x net021 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmmn3 net021 net015 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn2 net017 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn1 net125 d2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn0 net016 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn4 net018 net017 net015 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn3 net125 s1 net015 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn4 i0#2fnet20 net016 net018 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn3 i0#2fnet18 s0 net018 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn2 i0#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 i0#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmp4 x net021 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmmp3 net021 net015 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp2 net017 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 net125 d2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 net016 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp4 net018 s1 net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp3 net125 net017 net015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp4 i0#2fnet21 s0 net018 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fnet19 net016 net018 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 i0#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0 i0#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_MUXI3_4




.subckt SAEDRVT14_MUXI4_2 vdd vss vbp vbn x d0 d1 d2 d3 s0 s1
xmmn13 net18 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn12 x net15 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn5 net12 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn4 i2#2fnet20 net18 net15 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn3 i2#2fnet18 s1 net15 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn2 i2#2fnet20 net17 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 i2#2fnet18 net16 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn4 i1#2fnet20 net12 net17 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn3 i1#2fnet18 s0 net17 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn2 i1#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn0 i1#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net12 net16 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnet18 s0 net16 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet20 d2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fnet18 d3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmp13 net18 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp12 x net15 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp5 net12 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp4 i2#2fnet21 s1 net15 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp3 i2#2fnet19 net18 net15 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp2 i2#2fnet21 net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp0 i2#2fnet19 net16 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp4 i1#2fnet21 s0 net17 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp3 i1#2fnet19 net12 net17 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp2 i1#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 i1#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s0 net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fnet19 net12 net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet21 d2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet19 d3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_MUXI4_2




.subckt SAEDRVT14_MUXI4_4 vdd vss vbp vbn x d0 d1 d2 d3 s0 s1
xmmn13 net18 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn12 x net15 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn5 net12 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn4 i2#2fnet20 net18 net15 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn3 i2#2fnet18 s1 net15 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn2 i2#2fnet20 net17 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fn0 i2#2fnet18 net16 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fn4 i1#2fnet20 net12 net17 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn3 i1#2fnet18 s0 net17 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn2 i1#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn0 i1#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net12 net16 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnet18 s0 net16 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet20 d2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fnet18 d3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmp13 net18 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp12 x net15 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp5 net12 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp4 i2#2fnet21 s1 net15 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp3 i2#2fnet19 net18 net15 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp2 i2#2fnet21 net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi2#2fp0 i2#2fnet19 net16 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi1#2fp4 i1#2fnet21 s0 net17 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp3 i1#2fnet19 net12 net17 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp2 i1#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 i1#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s0 net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fnet19 net12 net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet21 d2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet19 d3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_MUXI4_4




.subckt SAEDRVT14_MUXI4_U_0P5 vdd vss vbp vbn x d0 d1 d2 d3 s0 s1
xmmn13 net18 s1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn12 x net15 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn5 net12 s0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn4 i2#2fnet20 net18 net15 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn3 i2#2fnet18 s1 net15 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn2 i2#2fnet20 net17 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fn0 i2#2fnet18 net16 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn4 i1#2fnet20 net12 net17 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn3 i1#2fnet18 s0 net17 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn2 i1#2fnet20 d0 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fn0 i1#2fnet18 d1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn4 i0#2fnet20 net12 net16 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn3 i0#2fnet18 s0 net16 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 i0#2fnet20 d2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fnet18 d3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmp13 net18 s1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp12 x net15 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp5 net12 s0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp4 i2#2fnet21 s1 net15 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp3 i2#2fnet19 net18 net15 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp2 i2#2fnet21 net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi2#2fp0 i2#2fnet19 net16 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp4 i1#2fnet21 s0 net17 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp3 i1#2fnet19 net12 net17 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp2 i1#2fnet21 d0 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi1#2fp0 i1#2fnet19 d1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp4 i0#2fnet21 s0 net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fnet19 net12 net16 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 i0#2fnet21 d2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp0 i0#2fnet19 d3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_MUXI4_U_0P5




.subckt SAEDRVT14_ND2_0P5 vdd vss vbp vbn x a1 a2
xmi0#2fmn1_2 x a1 i0#2fmidn_a_b_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn0_2 i0#2fmidn_a_b_2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn1 x a1 i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fmidn_a_b a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1_2 x a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp0_2 x a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 x a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 x a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ND2_0P5




.subckt SAEDRVT14_ND2_16 vdd vss vbp vbn x a1 a2
xmi0#2fn1_16 i0#2fmidn_a_b_16 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_15 i0#2fmidn_a_b_15 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_14 i0#2fmidn_a_b_14 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_13 i0#2fmidn_a_b_13 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_12 i0#2fmidn_a_b_12 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_11 i0#2fmidn_a_b_11 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_10 i0#2fmidn_a_b_10 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_9 i0#2fmidn_a_b_9 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_8 i0#2fmidn_a_b_8 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_7 i0#2fmidn_a_b_7 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_6 i0#2fmidn_a_b_6 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_5 i0#2fmidn_a_b_5 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_4 i0#2fmidn_a_b_4 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_3 i0#2fmidn_a_b_3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_2 i0#2fmidn_a_b_2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_16 x a1 i0#2fmidn_a_b_16 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_15 x a1 i0#2fmidn_a_b_15 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_14 x a1 i0#2fmidn_a_b_14 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_13 x a1 i0#2fmidn_a_b_13 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_12 x a1 i0#2fmidn_a_b_12 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_11 x a1 i0#2fmidn_a_b_11 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_10 x a1 i0#2fmidn_a_b_10 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_9 x a1 i0#2fmidn_a_b_9 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_8 x a1 i0#2fmidn_a_b_8 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_7 x a1 i0#2fmidn_a_b_7 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_6 x a1 i0#2fmidn_a_b_6 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_5 x a1 i0#2fmidn_a_b_5 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_4 x a1 i0#2fmidn_a_b_4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_3 x a1 i0#2fmidn_a_b_3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_2 x a1 i0#2fmidn_a_b_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1 i0#2fmidn_a_b a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 x a1 i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1_2 x a1 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=3
xmi0#2fp0_2 x a2 vdd vbp p08_rev l=0.014u nf=14 m=1 nfin=3
xmi0#2fp1 x a1 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=2
xmi0#2fp0 x a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_ND2_16




.subckt SAEDRVT14_ND2_1P5 vdd vss vbp vbn x a1 a2
xmi0#2fmn1_3 x a1 i0#2fmidn_a_b_3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1_2 x a1 i0#2fmidn_a_b_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn0_3 i0#2fmidn_a_b_3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn0_2 i0#2fmidn_a_b_2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 x a1 i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmn0 i0#2fmidn_a_b a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0_3 x a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 x a2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmi0#2fmp0 x a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_ND2_1P5




.subckt SAEDRVT14_ND2_1 vdd vss vbp vbn x a1 a2
xmi0#2fmn1_2 x a1 i0#2fmidn_a_b_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn0_2 i0#2fmidn_a_b_2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 x a1 i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn0 i0#2fmidn_a_b a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp1_2 x a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp0_2 x a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 x a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 x a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ND2_1




.subckt SAEDRVT14_ND2_2 vdd vss vbp vbn x a1 a2
xmi0#2fmn1_3 x a1 i0#2fmidn_a_b_3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1_2 x a1 i0#2fmidn_a_b_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn0_3 i0#2fmidn_a_b_3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn0_2 i0#2fmidn_a_b_2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn1 x a1 i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn0 i0#2fmidn_a_b a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0_3 x a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 x a2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmi0#2fmp0 x a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_ND2_2




.subckt SAEDRVT14_ND2_3 vdd vss vbp vbn x a1 a2
xmi0#2fn1_4 i0#2fmidn_a_b_4 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_3 i0#2fmidn_a_b_3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_2 i0#2fmidn_a_b_2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_4 x a1 i0#2fmidn_a_b_4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_3 x a1 i0#2fmidn_a_b_3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_2 x a1 i0#2fmidn_a_b_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1 i0#2fmidn_a_b a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 x a1 i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1_2 x a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi0#2fp0_2 x a2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmi0#2fp1 x a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp0 x a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ND2_3




.subckt SAEDRVT14_ND2_4 vdd vss vbp vbn x a1 a2
xmi0#2fn1_5 i0#2fmidn_a_b_5 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_4 i0#2fmidn_a_b_4 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_3 i0#2fmidn_a_b_3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_2 i0#2fmidn_a_b_2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_5 x a1 i0#2fmidn_a_b_5 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_4 x a1 i0#2fmidn_a_b_4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_3 x a1 i0#2fmidn_a_b_3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_2 x a1 i0#2fmidn_a_b_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1 i0#2fmidn_a_b a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 x a1 i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1_2 x a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi0#2fp1 x a1 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=2
xmi0#2fp0 x a2 vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=3
.ends SAEDRVT14_ND2_4




.subckt SAEDRVT14_ND2_5 vdd vss vbp vbn x a1 a2
xmi0#2fn1_6 i0#2fmidn_a_b_6 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_5 i0#2fmidn_a_b_5 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_4 i0#2fmidn_a_b_4 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_3 i0#2fmidn_a_b_3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_2 i0#2fmidn_a_b_2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_6 x a1 i0#2fmidn_a_b_6 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_5 x a1 i0#2fmidn_a_b_5 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_4 x a1 i0#2fmidn_a_b_4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_3 x a1 i0#2fmidn_a_b_3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_2 x a1 i0#2fmidn_a_b_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1 i0#2fmidn_a_b a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 x a1 i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1_2 x a1 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmi0#2fp1 x a1 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=2
xmi0#2fp0 x a2 vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=3
.ends SAEDRVT14_ND2_5




.subckt SAEDRVT14_ND2_6 vdd vss vbp vbn x a1 a2
xmi0#2fn1_7 i0#2fmidn_a_b_7 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_6 i0#2fmidn_a_b_6 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_5 i0#2fmidn_a_b_5 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_4 i0#2fmidn_a_b_4 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_3 i0#2fmidn_a_b_3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_2 i0#2fmidn_a_b_2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_7 x a1 i0#2fmidn_a_b_7 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_6 x a1 i0#2fmidn_a_b_6 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_5 x a1 i0#2fmidn_a_b_5 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_4 x a1 i0#2fmidn_a_b_4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_3 x a1 i0#2fmidn_a_b_3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_2 x a1 i0#2fmidn_a_b_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1 i0#2fmidn_a_b a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 x a1 i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1_2 x a1 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmi0#2fp1 x a1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmi0#2fp0 x a2 vdd vbp p08_rev l=0.014u nf=7 m=1 nfin=3
.ends SAEDRVT14_ND2_6




.subckt SAEDRVT14_ND2_8 vdd vss vbp vbn x a1 a2
xmi0#2fn1_9 i0#2fmidn_a_b_9 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_8 i0#2fmidn_a_b_8 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_7 i0#2fmidn_a_b_7 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_6 i0#2fmidn_a_b_6 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_5 i0#2fmidn_a_b_5 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_4 i0#2fmidn_a_b_4 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_3 i0#2fmidn_a_b_3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1_2 i0#2fmidn_a_b_2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_9 x a1 i0#2fmidn_a_b_9 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_8 x a1 i0#2fmidn_a_b_8 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_7 x a1 i0#2fmidn_a_b_7 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_6 x a1 i0#2fmidn_a_b_6 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_5 x a1 i0#2fmidn_a_b_5 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_4 x a1 i0#2fmidn_a_b_4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_3 x a1 i0#2fmidn_a_b_3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0_2 x a1 i0#2fmidn_a_b_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1 i0#2fmidn_a_b a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 x a1 i0#2fmidn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1_2 x a1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmi0#2fp1 x a1 vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=2
xmi0#2fp0 x a2 vdd vbp p08_rev l=0.014u nf=9 m=1 nfin=3
.ends SAEDRVT14_ND2_8




.subckt SAEDRVT14_ND2B_0P75 vdd vss vbp vbn x a b
xmn5 x int_zn yn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn4 yn int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn3 int_zn x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn2 midn_ab_b b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn1 x1 ab midn_ab_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn0 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 x int_zn yp vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 yp int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 int_zn x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmmp2 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmmp1 x1 b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmmp0 x1 ab vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ND2B_0P75




.subckt SAEDRVT14_ND2B_1P5 vdd vss vbp vbn x a b
xmn5 x int_zn yn vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn4 yn int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn3 int_zn x1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmmn2 midn_ab_b b vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmmn1 x1 ab midn_ab_b vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn0 ab a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmp5 x int_zn yp vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp4 yp int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp3 int_zn x1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmmp2 ab a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmmp1 x1 b vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmmp0 x1 ab vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_ND2B_1P5




.subckt SAEDRVT14_ND2B_1 vdd vss vbp vbn x a b
xmn5 x int_zn yn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn4 yn int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn3 int_zn x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn2 midn_ab_b b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn1 x1 ab midn_ab_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn0 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 x int_zn yp vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 yp int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 int_zn x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmmp2 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmmp1 x1 b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmmp0 x1 ab vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ND2B_1




.subckt SAEDRVT14_ND2B_2 vdd vss vbp vbn x a b
xmn5 x int_zn yn vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn4 yn int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn3 int_zn x1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmmn2 midn_ab_b b vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmmn1 x1 ab midn_ab_b vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmmn0 ab a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmp5 x int_zn yp vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp4 yp int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp3 int_zn x1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmmp2 ab a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmmp1 x1 b vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmmp0 x1 ab vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_ND2B_2




.subckt SAEDRVT14_ND2B_4 vdd vss vbp vbn x a b
xmn5 x int_zn yn vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn4 yn int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn3 int_zn x1 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmn2 ab a vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn1 midn_ab_b b vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn0 x1 ab midn_ab_b vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp5 x int_zn yp vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp4 yp int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp3 int_zn x1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp2 ab a vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp1 x1 ab vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmp0 x1 b vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
.ends SAEDRVT14_ND2B_4




.subckt SAEDRVT14_ND2B_U_0P5 vdd vss vbp vbn x a b
xmn2 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 midn_ab_b b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 x ab midn_ab_b vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 x ab vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 x b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ND2B_U_0P5




.subckt SAEDRVT14_ND2_CDC_0P5 vdd vss vbp vbn x a1 a2
xmn1 midn_a_b a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x a2 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ND2_CDC_0P5




.subckt SAEDRVT14_ND2_CDC_1 vdd vss vbp vbn x a1 a2
xmmn1 x a2 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn0 midn_a_b a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 x a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmmp0 x a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ND2_CDC_1




.subckt SAEDRVT14_ND2_CDC_2 vdd vss vbp vbn x a1 a2
xmmn11 x a2 midn_a_b1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn01 midn_a_b1 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn1 x a2 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn0 midn_a_b a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 x a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmmp0 x a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_ND2_CDC_2




.subckt SAEDRVT14_ND2_CDC_4 vdd vss vbp vbn x a1 a2
xmn13 midn_a_b3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 midn_a_b2 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn11 midn_a_b1 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn03 x a2 midn_a_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn02 x a2 midn_a_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn01 x a2 midn_a_b1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_a_b a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x a2 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x a2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp0 x a1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_ND2_CDC_4




.subckt SAEDRVT14_ND2_ECO_1 vdd vss vbp vbn x a1 a2
xmn1 midn_a_b a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x a1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 x a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ND2_ECO_1




.subckt SAEDRVT14_ND2_ECO_2 vdd vss vbp vbn x a1 a2
xmn11 midn_a_b1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn01 x a1 midn_a_b1 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 midn_a_b a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x a1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp0 x a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_ND2_ECO_2




.subckt SAEDRVT14_ND2_MM_0P5 vdd vss vbp vbn x a1 a2
xmn1 midn_en_ck a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn0 x a1 midn_en_ck vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp1 x a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 x a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ND2_MM_0P5




.subckt SAEDRVT14_ND2_MM_10 vdd vss vbp vbn x a1 a2
xmnfet x a1 midn_en_ck8 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn19 midn_en_ck9 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn18 midn_en_ck8 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn17 midn_en_ck7 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn16 midn_en_ck6 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn15 midn_en_ck5 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn14 midn_en_ck4 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn13 midn_en_ck3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 midn_en_ck2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn11 midn_en_ck1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn09 x a1 midn_en_ck9 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn07 x a1 midn_en_ck7 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn06 x a1 midn_en_ck6 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn05 x a1 midn_en_ck5 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn04 x a1 midn_en_ck4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn03 x a1 midn_en_ck3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn02 x a1 midn_en_ck2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn01 x a1 midn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_en_ck a2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn0 x a1 midn_en_ck vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 x a1 vdd vbp p08_rev l=0.014u nf=10 m=1 nfin=3
xmp0 x a2 vdd vbp p08_rev l=0.014u nf=10 m=1 nfin=3
.ends SAEDRVT14_ND2_MM_10




.subckt SAEDRVT14_ND2_MM_12 vdd vss vbp vbn x a1 a2
xmnfet x a1 midn_en_ck8 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn102 midn_en_ck02 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn101 midn_en_ck01 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn002 x a1 midn_en_ck02 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn001 x a1 midn_en_ck01 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn19 midn_en_ck9 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn18 midn_en_ck8 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn17 midn_en_ck7 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn16 midn_en_ck6 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn15 midn_en_ck5 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn14 midn_en_ck4 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn13 midn_en_ck3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 midn_en_ck2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn11 midn_en_ck1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn09 x a1 midn_en_ck9 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn07 x a1 midn_en_ck7 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn06 x a1 midn_en_ck6 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn05 x a1 midn_en_ck5 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn04 x a1 midn_en_ck4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn03 x a1 midn_en_ck3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn02 x a1 midn_en_ck2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn01 x a1 midn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_en_ck a2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn0 x a1 midn_en_ck vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 x a1 vdd vbp p08_rev l=0.014u nf=12 m=1 nfin=3
xmp0 x a2 vdd vbp p08_rev l=0.014u nf=12 m=1 nfin=3
.ends SAEDRVT14_ND2_MM_12




.subckt SAEDRVT14_ND2_MM_16 vdd vss vbp vbn x a1 a2
xmn115 midn_en_ck115 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn114 midn_en_ck114 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn113 midn_en_ck113 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn112 midn_en_ck112 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn111 midn_en_ck111 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn110 midn_en_ck110 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn109 midn_en_ck109 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn108 midn_en_ck108 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn107 midn_en_ck107 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn106 midn_en_ck106 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn105 midn_en_ck105 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn104 midn_en_ck104 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn103 midn_en_ck103 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn102 midn_en_ck102 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn101 midn_en_ck101 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn015 x a1 midn_en_ck115 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn014 x a1 midn_en_ck114 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn013 x a1 midn_en_ck113 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn012 x a1 midn_en_ck112 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn011 x a1 midn_en_ck111 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn010 x a1 midn_en_ck110 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn009 x a1 midn_en_ck109 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn008 x a1 midn_en_ck108 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn007 x a1 midn_en_ck107 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn006 x a1 midn_en_ck106 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn005 x a1 midn_en_ck105 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn004 x a1 midn_en_ck104 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn003 x a1 midn_en_ck103 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn002 x a1 midn_en_ck102 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn001 x a1 midn_en_ck101 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_en_ck a2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn0 x a1 midn_en_ck vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 x a1 vdd vbp p08_rev l=0.014u nf=16 m=1 nfin=3
xmp0 x a2 vdd vbp p08_rev l=0.014u nf=16 m=1 nfin=3
.ends SAEDRVT14_ND2_MM_16




.subckt SAEDRVT14_ND2_MM_1 vdd vss vbp vbn x a1 a2
xmn1 midn_en_ck a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn0 x a1 midn_en_ck vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 x a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ND2_MM_1




.subckt SAEDRVT14_ND2_MM_2 vdd vss vbp vbn x a1 a2
xmn11 midn_en_ck1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn01 x a1 midn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_en_ck a2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn0 x a1 midn_en_ck vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 x a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp0 x a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_ND2_MM_2




.subckt SAEDRVT14_ND2_MM_3 vdd vss vbp vbn x a1 a2
xmn1 midn_en_ck a2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn0 x a1 midn_en_ck vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 x a1 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmp0 x a2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
.ends SAEDRVT14_ND2_MM_3




.subckt SAEDRVT14_ND2_MM_4 vdd vss vbp vbn x a1 a2
xmn13 midn_en_ck3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 midn_en_ck2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn11 midn_en_ck1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn03 x a1 midn_en_ck3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn02 x a1 midn_en_ck2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn01 x a1 midn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_en_ck a2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn0 x a1 midn_en_ck vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 x a1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp0 x a2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
.ends SAEDRVT14_ND2_MM_4




.subckt SAEDRVT14_ND2_MM_6 vdd vss vbp vbn x a1 a2
xmn15 midn_en_ck5 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn14 midn_en_ck4 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn13 midn_en_ck3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 midn_en_ck2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn11 midn_en_ck1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn05 x a1 midn_en_ck5 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn04 x a1 midn_en_ck4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn03 x a1 midn_en_ck3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn02 x a1 midn_en_ck2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn01 x a1 midn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_en_ck a2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn0 x a1 midn_en_ck vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 x a1 vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=3
xmp0 x a2 vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=3
.ends SAEDRVT14_ND2_MM_6




.subckt SAEDRVT14_ND2_MM_8 vdd vss vbp vbn x a1 a2
xmn17 midn_en_ck7 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn16 midn_en_ck6 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn15 midn_en_ck5 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn14 midn_en_ck4 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn13 midn_en_ck3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 midn_en_ck2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn11 midn_en_ck1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn07 x a1 midn_en_ck7 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn06 x a1 midn_en_ck6 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn05 x a1 midn_en_ck5 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn04 x a1 midn_en_ck4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn03 x a1 midn_en_ck3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn02 x a1 midn_en_ck2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn01 x a1 midn_en_ck1 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_en_ck a2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn0 x a1 midn_en_ck vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 x a1 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=3
xmp0 x a2 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=3
.ends SAEDRVT14_ND2_MM_8




.subckt SAEDRVT14_ND3_0P5 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 midn_b_c a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ND3_0P5




.subckt SAEDRVT14_ND3_0P75 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 midn_b_c a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ND3_0P75




.subckt SAEDRVT14_ND3_1 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 midn_b_c a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ND3_1




.subckt SAEDRVT14_ND3_2 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn1_2 midn_a_b_2 a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0_2 x1 a1 midn_a_b_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 midn_b_c a3 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_ND3_2




.subckt SAEDRVT14_ND3_3 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmn2 midn_b_c a3 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=2
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
.ends SAEDRVT14_ND3_3




.subckt SAEDRVT14_ND3_4 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmn13 midn_a_b3 a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 midn_a_b2 a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn11 midn_a_b1 a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn03 x1 a1 midn_a_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn02 x1 a1 midn_a_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn01 x1 a1 midn_a_b1 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 midn_b_c a3 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
.ends SAEDRVT14_ND3_4




.subckt SAEDRVT14_ND3_8 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=2
xmn17 midn_a_b7 a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn16 midn_a_b6 a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn15 midn_a_b5 a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn14 midn_a_b4 a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn13 midn_a_b3 a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn12 midn_a_b2 a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn11 midn_a_b1 a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn07 x1 a1 midn_a_b7 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn06 x1 a1 midn_a_b6 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn05 x1 a1 midn_a_b5 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn04 x1 a1 midn_a_b4 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn03 x1 a1 midn_a_b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn02 x1 a1 midn_a_b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn01 x1 a1 midn_a_b1 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 midn_b_c a3 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=3
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=2
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=3
.ends SAEDRVT14_ND3_8




.subckt SAEDRVT14_ND3B_0P5 vdd vss vbp vbn x a b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 midn_b_c b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 midn_ab_b b1 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 x1 ab midn_ab_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x1 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 x1 ab vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 x1 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ND3B_0P5




.subckt SAEDRVT14_ND3B_0P75 vdd vss vbp vbn x a b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 midn_b_c b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 midn_ab_b b1 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 x1 ab midn_ab_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x1 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 x1 ab vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 x1 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ND3B_0P75




.subckt SAEDRVT14_ND3B_1 vdd vss vbp vbn x a b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 midn_b_c b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 midn_ab_b b1 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 x1 ab midn_ab_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x1 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 x1 ab vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 x1 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_ND3B_1




.subckt SAEDRVT14_ND3B_2 vdd vss vbp vbn x a b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn2_2 midn_b_c_2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1_2 midn_ab_b b1 midn_b_c_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 ab a vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn2 midn_b_c b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_ab_b b1 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x1 ab midn_ab_b vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp3 ab a vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp2 x1 b2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 x1 ab vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp0 x1 b1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_ND3B_2




.subckt SAEDRVT14_ND3B_4 vdd vss vbp vbn x a b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmn2_4 midn_b_c_4 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2_3 midn_b_c_3 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2_2 midn_b_c_2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1_4 midn_ab_b b1 midn_b_c_4 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1_3 midn_ab_b b1 midn_b_c_3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1_2 midn_ab_b b1 midn_b_c_2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 ab a vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn2 midn_b_c b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_ab_b b1 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x1 ab midn_ab_b vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp3 ab a vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp2 x1 b2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 x1 ab vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp0 x1 b1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_ND3B_4




.subckt SAEDRVT14_ND3_ECO_1 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 midn_b_c a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_ND3_ECO_1




.subckt SAEDRVT14_ND4_0P5 vdd vss vbp vbn x a1 a2 a3 a4
xmn6 x int_zn yn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn5 yn int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 int_zn x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_c_d a4 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn2 midn_b_c a3 midn_c_d vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp6 x int_zn yp vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp5 yp int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 int_zn x1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp3 x1 a4 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ND4_0P5




.subckt SAEDRVT14_ND4_0P75 vdd vss vbp vbn x a1 a2 a3 a4
xmn6 x int_zn yn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn5 yn int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 int_zn x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_c_d a4 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn2 midn_b_c a3 midn_c_d vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp6 x int_zn yp vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp5 yp int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 int_zn x1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp3 x1 a4 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ND4_0P75




.subckt SAEDRVT14_ND4_1 vdd vss vbp vbn x a1 a2 a3 a4
xmn6 x int_zn yn vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn5 yn int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn4 int_zn x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_c_d a4 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn2 midn_b_c a3 midn_c_d vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp6 x int_zn yp vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp5 yp int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp4 int_zn x1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp3 x1 a4 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_ND4_1




.subckt SAEDRVT14_ND4_2 vdd vss vbp vbn x a1 a2 a3 a4
xmn6 x int_zn yn vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn5 yn int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn4 int_zn x1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn3 midn_c_d a4 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn2 midn_b_c a3 midn_c_d vbn n08_rev l=0.014u nf=5 m=1 nfin=2
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp6 x int_zn yp vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp5 yp int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp4 int_zn x1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp3 x1 a4 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_ND4_2




.subckt SAEDRVT14_ND4_3 vdd vss vbp vbn x a1 a2 a3 a4
xmn6 x int_zn yn vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn5 yn int_zn vss vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn4 int_zn x1 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmn3 midn_c_d a4 vss vbn n08_rev l=0.014u nf=7 m=1 nfin=2
xmn2 midn_b_c a3 midn_c_d vbn n08_rev l=0.014u nf=7 m=1 nfin=2
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp6 x int_zn yp vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmp5 yp int_zn vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=3
xmp4 int_zn x1 vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=3
xmp3 x1 a4 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
.ends SAEDRVT14_ND4_3




.subckt SAEDRVT14_ND4_4 vdd vss vbp vbn x a1 a2 a3 a4
xmn6 x int_zn yn vbn n08_rev l=0.014u nf=8 m=1 nfin=3
xmn5 yn int_zn vss vbn n08_rev l=0.014u nf=8 m=1 nfin=3
xmn4 int_zn x1 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmn3 midn_c_d a4 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn2 midn_b_c a3 midn_c_d vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp6 x int_zn yp vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmp5 yp int_zn vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=3
xmp4 int_zn x1 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=3
xmp3 x1 a4 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
.ends SAEDRVT14_ND4_4




.subckt SAEDRVT14_ND4_8 vdd vss vbp vbn x a1 a2 a3 a4
xmn6 x int_zn yn vbn n08_rev l=0.014u nf=16 m=1 nfin=3
xmn5 yn int_zn vss vbn n08_rev l=0.014u nf=16 m=1 nfin=3
xmn4 int_zn x1 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=2
xmn3 midn_c_d a4 vss vbn n08_rev l=0.014u nf=10 m=1 nfin=4
xmn2 midn_b_c a3 midn_c_d vbn n08_rev l=0.014u nf=10 m=1 nfin=4
xmn1 midn_a_b a2 midn_b_c vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmn0 x1 a1 midn_a_b vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmp6 x int_zn yp vbp p08_rev l=0.014u nf=16 m=1 nfin=4
xmp5 yp int_zn vdd vbp p08_rev l=0.014u nf=16 m=1 nfin=3
xmp4 int_zn x1 vdd vbp p08_rev l=0.014u nf=16 m=1 nfin=3
xmp3 x1 a4 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=3
xmp2 x1 a3 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=3
xmp1 x1 a1 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=3
xmp0 x1 a2 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=3
.ends SAEDRVT14_ND4_8




.subckt SAEDRVT14_NR2_0P5 vdd vss vbp vbn x a1 a2
xmi0#2fn1 x a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 x a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp1 x a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_0P5




.subckt SAEDRVT14_NR2_16 vdd vss vbp vbn x a1 a2
xmi0#2fn1 x a1 vss vbn n08_rev l=0.014u nf=16 m=1 nfin=2
xmi0#2fn0 x a2 vss vbn n08_rev l=0.014u nf=16 m=1 nfin=2
xmi0#2fpfet x a1 i0#2fmidp_a_b8 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp115 i0#2fmidp_a_b15 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp114 i0#2fmidp_a_b14 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp113 i0#2fmidp_a_b13 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp112 i0#2fmidp_a_b12 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp111 i0#2fmidp_a_b11 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp110 i0#2fmidp_a_b10 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp015 x a1 i0#2fmidp_a_b15 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp014 x a1 i0#2fmidp_a_b14 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp013 x a1 i0#2fmidp_a_b13 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp012 x a1 i0#2fmidp_a_b12 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp011 x a1 i0#2fmidp_a_b11 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp010 x a1 i0#2fmidp_a_b10 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp19 i0#2fmidp_a_b9 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp18 i0#2fmidp_a_b8 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp17 i0#2fmidp_a_b7 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp16 i0#2fmidp_a_b6 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp15 i0#2fmidp_a_b5 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp14 i0#2fmidp_a_b4 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp13 i0#2fmidp_a_b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp12 i0#2fmidp_a_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp11 i0#2fmidp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp09 x a1 i0#2fmidp_a_b9 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp07 x a1 i0#2fmidp_a_b7 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp06 x a1 i0#2fmidp_a_b6 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp05 x a1 i0#2fmidp_a_b5 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp04 x a1 i0#2fmidp_a_b4 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp03 x a1 i0#2fmidp_a_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp02 x a1 i0#2fmidp_a_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp01 x a1 i0#2fmidp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp0 x a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_16




.subckt SAEDRVT14_NR2_1P5 vdd vss vbp vbn x a1 a2
xmi0#2fmn1 x a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn0 x a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp11 x a1 i0#2fmidp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp01 i0#2fmidp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp1 x a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fmp0 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_NR2_1P5




.subckt SAEDRVT14_NR2_1 vdd vss vbp vbn x a1 a2
xmi0#2fn1 x a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 x a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 x a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp0 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_NR2_1




.subckt SAEDRVT14_NR2_2 vdd vss vbp vbn x a1 a2
xmi0#2fmn1 x a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmn0 x a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp11 x a1 i0#2fmidp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp01 i0#2fmidp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fmp1 x a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fmp0 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_NR2_2




.subckt SAEDRVT14_NR2_3 vdd vss vbp vbn x a1 a2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 x1 a1 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmi0#2fn0 x1 a2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp1 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmi0#2fp0 x1 a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_NR2_3




.subckt SAEDRVT14_NR2_4 vdd vss vbp vbn x a1 a2
xmi0#2fn1 x a1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn0 x a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp13 i0#2fmidp_a_b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fmidp_a_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp11 i0#2fmidp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp03 x a1 i0#2fmidp_a_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp02 x a1 i0#2fmidp_a_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp01 x a1 i0#2fmidp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp0 x a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_4




.subckt SAEDRVT14_NR2_5 vdd vss vbp vbn x a1 a2
xm1 vss net21 x vbn n08_rev l=0.014u nf=5 m=1 nfin=4
xm0 vss net26 net21 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn1 net26 a1 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmi0#2fn0 net26 a2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xm3 vdd net21 x vbp p08_rev l=0.014u nf=5 m=1 nfin=4
xm2 vdd net26 net21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp1 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
xmi0#2fp0 net26 a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_NR2_5




.subckt SAEDRVT14_NR2_6 vdd vss vbp vbn x a1 a2
xmi0#2fn1 x a1 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=2
xmi0#2fn0 x a2 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=2
xmi0#2fp15 i0#2fmidp_a_b5 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp14 i0#2fmidp_a_b4 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp13 i0#2fmidp_a_b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp12 i0#2fmidp_a_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp11 i0#2fmidp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp05 x a1 i0#2fmidp_a_b5 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp04 x a1 i0#2fmidp_a_b4 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp03 x a1 i0#2fmidp_a_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp02 x a1 i0#2fmidp_a_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp01 x a1 i0#2fmidp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp0 x a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_6




.subckt SAEDRVT14_NR2_8 vdd vss vbp vbn x a1 a2
xmi0#2fn1 x a1 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=2
xmi0#2fn0 x a2 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=2
xmi0#2fp17 i0#2fmidp_a_b7 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp16 i0#2fmidp_a_b6 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp15 i0#2fmidp_a_b5 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp14 i0#2fmidp_a_b4 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp13 i0#2fmidp_a_b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp12 i0#2fmidp_a_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp11 i0#2fmidp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp07 x a1 i0#2fmidp_a_b7 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp06 x a1 i0#2fmidp_a_b6 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp05 x a1 i0#2fmidp_a_b5 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp04 x a1 i0#2fmidp_a_b4 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp03 x a1 i0#2fmidp_a_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp02 x a1 i0#2fmidp_a_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp01 x a1 i0#2fmidp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp0 x a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_8




.subckt SAEDRVT14_NR2B_0P75 vdd vss vbp vbn x a b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn2 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn1 x1 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn0 x1 ab vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp2 midp_ab_b b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 x1 ab midp_ab_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp0 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_NR2B_0P75




.subckt SAEDRVT14_NR2B_1P5 vdd vss vbp vbn x a b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn2 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn1 x1 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn0 x1 ab vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmmp2 midp_ab_b b vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmmp1 x1 ab midp_ab_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp0 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_NR2B_1P5




.subckt SAEDRVT14_NR2B_1 vdd vss vbp vbn x a b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn2 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn1 x1 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn0 x1 ab vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmmp2 midp_ab_b b vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmmp1 x1 ab midp_ab_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp0 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_NR2B_1




.subckt SAEDRVT14_NR2B_2 vdd vss vbp vbn x a b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn2 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn1 x1 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn0 x1 ab vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp2 midp_ab_b b vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmmp1 x1 ab midp_ab_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp0 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_NR2B_2




.subckt SAEDRVT14_NR2B_4 vdd vss vbp vbn x a b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn2 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn1 x1 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn0 x1 ab vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmmp2 midp_ab_b b vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmmp1 x1 ab midp_ab_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmmp0 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_NR2B_4




.subckt SAEDRVT14_NR2B_U_0P5 vdd vss vbp vbn x a b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 x1 ab vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 x1 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 midp_ab_b b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 x1 ab midp_ab_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_NR2B_U_0P5




.subckt SAEDRVT14_NR2_ECO_1 vdd vss vbp vbn x a1 a2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 x1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 x1 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 x1 a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_ECO_1




.subckt SAEDRVT14_NR2_ECO_2 vdd vss vbp vbn x a1 a2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 x1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 x1 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 x1 a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 midp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_ECO_2




.subckt SAEDRVT14_NR2_ISO_1 vdd vss vbp vbn x ck en
xmi0#2fn1 x en vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 x ck vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 x ck i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp0 i0#2fmidp_a_b en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_NR2_ISO_1




.subckt SAEDRVT14_NR2_ISO_4 vdd vss vbp vbn x ck en
xmi0#2fn1 x ck vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn0 x en vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp13 i0#2fmidp_a_b3 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp12 i0#2fmidp_a_b2 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp11 i0#2fmidp_a_b1 en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp03 x ck i0#2fmidp_a_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp02 x ck i0#2fmidp_a_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp01 x ck i0#2fmidp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1 i0#2fmidp_a_b en vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp0 x ck i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_ISO_4




.subckt SAEDRVT14_NR2_MM_0P5 vdd vss vbp vbn x a1 a2
xmmn1 x a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmn0 x a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmmp1 midp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmmp0 x a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_NR2_MM_0P5




.subckt SAEDRVT14_NR2_MM_10 vdd vss vbp vbn x a1 a2
xmmn1 x a2 vss vbn n08_rev l=0.014u nf=10 m=1 nfin=3
xmmn0 x a1 vss vbn n08_rev l=0.014u nf=10 m=1 nfin=3
xmmpfet x a1 midp_a_b8 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp19 midp_a_b9 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp18 midp_a_b8 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp17 midp_a_b7 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp16 midp_a_b6 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp15 midp_a_b5 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp14 midp_a_b4 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp13 midp_a_b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp12 midp_a_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp11 midp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp09 x a1 midp_a_b9 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp07 x a1 midp_a_b7 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp06 x a1 midp_a_b6 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp05 x a1 midp_a_b5 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp04 x a1 midp_a_b4 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp03 x a1 midp_a_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp02 x a1 midp_a_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp01 x a1 midp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 midp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 x a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_MM_10




.subckt SAEDRVT14_NR2_MM_12 vdd vss vbp vbn x a1 a2
xmmn1 x a2 vss vbn n08_rev l=0.014u nf=12 m=1 nfin=3
xmmn0 x a1 vss vbn n08_rev l=0.014u nf=12 m=1 nfin=3
xmmp111 midp_a_b011 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp110 midp_a_b010 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp109 midp_a_b009 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp108 midp_a_b008 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp107 midp_a_b007 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp106 midp_a_b006 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp105 midp_a_b005 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp104 midp_a_b004 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp103 midp_a_b003 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp102 midp_a_b002 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp101 midp_a_b001 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp011 x a1 midp_a_b011 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp010 x a1 midp_a_b010 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp009 x a1 midp_a_b009 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp008 x a1 midp_a_b008 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp007 x a1 midp_a_b007 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp006 x a1 midp_a_b006 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp005 x a1 midp_a_b005 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp004 x a1 midp_a_b004 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp003 x a1 midp_a_b003 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp002 x a1 midp_a_b002 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp001 x a1 midp_a_b001 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 midp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 x a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_MM_12




.subckt SAEDRVT14_NR2_MM_16 vdd vss vbp vbn x a1 a2
xmmn1 x a2 vss vbn n08_rev l=0.014u nf=16 m=1 nfin=3
xmmn0 x a1 vss vbn n08_rev l=0.014u nf=16 m=1 nfin=3
xmmp115 midp_a_b015 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp114 midp_a_b014 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp113 midp_a_b013 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp112 midp_a_b012 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp111 midp_a_b011 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp110 midp_a_b010 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp109 midp_a_b009 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp108 midp_a_b008 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp107 midp_a_b007 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp106 midp_a_b006 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp105 midp_a_b005 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp104 midp_a_b004 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp103 midp_a_b003 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp102 midp_a_b002 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp101 midp_a_b001 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp015 x a1 midp_a_b015 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp014 x a1 midp_a_b014 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp013 x a1 midp_a_b013 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp012 x a1 midp_a_b012 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp011 x a1 midp_a_b011 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp010 x a1 midp_a_b010 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp009 x a1 midp_a_b009 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp008 x a1 midp_a_b008 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp007 x a1 midp_a_b007 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp006 x a1 midp_a_b006 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp005 x a1 midp_a_b005 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp004 x a1 midp_a_b004 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp003 x a1 midp_a_b003 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp002 x a1 midp_a_b002 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp001 x a1 midp_a_b001 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 midp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 x a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_MM_16




.subckt SAEDRVT14_NR2_MM_1 vdd vss vbp vbn x a1 a2
xmmn1 x a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmn0 x a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmmp1 midp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 x a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_MM_1




.subckt SAEDRVT14_NR2_MM_2 vdd vss vbp vbn x a1 a2
xmmn1 x a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmmn0 x a1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmmp11 midp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp01 x a1 midp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 midp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 x a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_MM_2




.subckt SAEDRVT14_NR2_MM_3 vdd vss vbp vbn x a1 a2
xmmn1 x a2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmmn0 x a1 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=2
xmmp1 midp_a_b a2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmmp0 x a1 midp_a_b vbp p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_NR2_MM_3




.subckt SAEDRVT14_NR2_MM_4 vdd vss vbp vbn x a1 a2
xmmn1 x a2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmmn0 x a1 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmmp13 midp_a_b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp12 midp_a_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp11 midp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp03 x a1 midp_a_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp02 x a1 midp_a_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp01 x a1 midp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 midp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 x a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_MM_4




.subckt SAEDRVT14_NR2_MM_6 vdd vss vbp vbn x a1 a2
xmmn1 x a2 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmmn0 x a1 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmmp15 midp_a_b5 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp14 midp_a_b4 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp13 midp_a_b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp12 midp_a_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp11 midp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp05 x a1 midp_a_b5 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp04 x a1 midp_a_b4 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp03 x a1 midp_a_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp02 x a1 midp_a_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp01 x a1 midp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 midp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 x a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_MM_6




.subckt SAEDRVT14_NR2_MM_8 vdd vss vbp vbn x a1 a2
xmmn1 x a2 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=3
xmmn0 x a1 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=3
xmmp17 midp_a_b7 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp16 midp_a_b6 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp15 midp_a_b5 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp14 midp_a_b4 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp13 midp_a_b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp12 midp_a_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp11 midp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp07 x a1 midp_a_b7 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp06 x a1 midp_a_b6 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp05 x a1 midp_a_b5 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp04 x a1 midp_a_b4 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp03 x a1 midp_a_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp02 x a1 midp_a_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp01 x a1 midp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 midp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 x a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR2_MM_8




.subckt SAEDRVT14_NR3_0P5 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 x1 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x1 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 x1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_b_c a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_NR3_0P5




.subckt SAEDRVT14_NR3_0P75 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 x1 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 x1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_b_c a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 x1 a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR3_0P75




.subckt SAEDRVT14_NR3_1 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 x1 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 x1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_b_c a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 x1 a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR3_1




.subckt SAEDRVT14_NR3_2 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 x1 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 x1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_b_c a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 x1 a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR3_2




.subckt SAEDRVT14_NR3_3 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn2 x1 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 x1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp2 midp_b_c a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 x1 a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR3_3




.subckt SAEDRVT14_NR3_4 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmn2 x1 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x1 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 x1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=2
xmp2 midp_b_c a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 x1 a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR3_4




.subckt SAEDRVT14_NR3_8 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmn2 x1 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x1 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 x1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=2
xmp2 midp_b_c a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 x1 a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR3_8




.subckt SAEDRVT14_NR3B_0P75 vdd vss vbp vbn x a b1 b2
xm2 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xm3 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 x1 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 x1 ab vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 x1 b1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xm0 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xm1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_b_c b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_ab_b b1 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 ab midp_ab_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_NR3B_0P75




.subckt SAEDRVT14_NR3B_1P5 vdd vss vbp vbn x a b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x1 b2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn1 x1 ab vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn0 x1 b1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp21 midp_b_c1 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp11 midp_ab_b b1 midp_b_c1 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_b_c b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_ab_b b1 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 ab midp_ab_b vbp p08_rev l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_NR3B_1P5




.subckt SAEDRVT14_NR3B_4 vdd vss vbp vbn x a b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 x1 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 x1 ab vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 x1 b1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 midp_b_c b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_ab_b b1 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 x1 ab midp_ab_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR3B_1




.subckt SAEDRVT14_NR3B_2 vdd vss vbp vbn x a b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x1 b2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn1 x1 ab vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn0 x1 b1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp21 midp_b_c1 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp11 midp_ab_b b1 midp_b_c1 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_b_c b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_ab_b b1 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 ab midp_ab_b vbp p08_rev l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_NR3B_2




.subckt SAEDRVT14_NR3B_4 vdd vss vbp vbn x a b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn3 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x1 b2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmn1 x1 ab vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmn0 x1 b1 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp23 midp_b_c3 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp22 midp_b_c2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp21 midp_b_c1 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp13 midp_ab_b b1 midp_b_c3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp12 midp_ab_b b1 midp_b_c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp11 midp_ab_b b1 midp_b_c1 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_b_c b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_ab_b b1 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 ab midp_ab_b vbp p08_rev l=0.014u nf=4 m=1 nfin=2
.ends SAEDRVT14_NR3B_4




.subckt SAEDRVT14_NR3B_U_0P5 vdd vss vbp vbn x a b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 ab a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x1 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 x1 ab vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 x1 b1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 ab a vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_b_c b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 midp_ab_b b1 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 x1 ab midp_ab_b vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_NR3B_U_0P5




.subckt SAEDRVT14_NR3_ECO_1 vdd vss vbp vbn x a1 a2 a3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 x1 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 x1 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn0 x1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_b_c a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 x1 a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR3_ECO_1




.subckt SAEDRVT14_NR4_0P75 vdd vss vbp vbn x a1 a2 a3 a4
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 x1 a4 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x1 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 x1 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 x1 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_c_d a4 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 midp_b_c a3 midp_c_d vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_NR4_0P75




.subckt SAEDRVT14_NR4_2 vdd vss vbp vbn x a1 a2 a3 a4
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 x1 a4 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn2 x1 a3 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn1 x1 a1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn0 x1 a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp32 midp_c_d2 a4 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp22 midp_b_c a3 midp_c_d2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp12 midp_a_b2 a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp02 x1 a1 midp_a_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 midp_c_d a4 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 midp_b_c a3 midp_c_d vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 x1 a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_NR4_2




.subckt SAEDRVT14_OA211_1 vdd vss vbp vbn x a1 a2 b1 b2
xn5 x int_zn vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn4 vss a2 midn_a1a2_b vbn n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 midn_b_c b1 int_zn vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn1 vss a1 midn_a1a2_b vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn0 midn_a1a2_b b2 midn_b_c vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xp7 midp_a1_a2 a2 vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=3
xp6 x int_zn vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp5 int_zn a1 midp_a1_a2 vbp p08_rev2 l=0.014u nf=2 m=1 nfin=3
xp4 int_zn b2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 int_zn b1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OA211_1




.subckt SAEDRVT14_OA211_2 vdd vss vbp vbn x a1 a2 b1 b2
xn5 x int_zn vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn4 vss a2 midn_a1a2_b vbn n08_rev2 l=0.014u nf=6 m=1 nfin=3
xn2 midn_b_c b1 int_zn vbn n08_rev2 l=0.014u nf=2 m=1 nfin=3
xn1 vss a1 midn_a1a2_b vbn n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn0 midn_a1a2_b b2 midn_b_c vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xp7 midp_a1_a2 a2 vdd vbp p08_rev2 l=0.014u nf=4 m=1 nfin=3
xp6 x int_zn vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp5 int_zn a1 midp_a1_a2 vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 int_zn b2 vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=2
xp3 int_zn b1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA211_2




.subckt SAEDRVT14_OA211_4 vdd vss vbp vbn x a1 a2 b1 b2
xn5 x int_zn vss vbn n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn4 vss a2 midn_a1a2_b vbn n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn2 midn_b_c b1 int_zn vbn n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn1 vss a1 midn_a1a2_b vbn n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn0 midn_a1a2_b b2 midn_b_c vbn n08_rev2 l=0.014u nf=4 m=1 nfin=4
xp7 midp_a1_a2 a2 vdd vbp p08_rev2 l=0.014u nf=6 m=1 nfin=3
xp6 x int_zn vdd vbp p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp5 int_zn a1 midp_a1_a2 vbp p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp4 int_zn b2 vdd vbp p08_rev2 l=0.014u nf=4 m=1 nfin=2
xp3 int_zn b1 vdd vbp p08_rev2 l=0.014u nf=3 m=1 nfin=2
.ends SAEDRVT14_OA211_4




.subckt SAEDRVT14_OA21_1 vdd vss vbp vbn x a1 a2 b
xmn4 vss a2 midn_a1a2_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn3 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 vss a1 midn_a1a2_b vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_a1a2_b b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp4 int_zn a1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 int_zn b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA21_1




.subckt SAEDRVT14_OA211_U_0P5 vdd vss vbp vbn x a1 a2 b1 b2
xn5 x int_zn vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn4 vss a2 midn_a1a2_b vbn n08_rev2 l=0.014u nf=5 m=1 nfin=2
xn2 midn_b_c b1 int_zn vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn1 vss a1 midn_a1a2_b vbn n08_rev2 l=0.014u nf=2 m=1 nfin=3
xn0 midn_a1a2_b b2 midn_b_c vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xp7 midp_a1_a2 a2 vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=3
xp6 x int_zn vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp5 int_zn a1 midp_a1_a2 vbp p08_rev2 l=0.014u nf=2 m=1 nfin=3
xp4 int_zn b2 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 int_zn b1 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OA211_U_0P5




.subckt SAEDRVT14_OA21_2 vdd vss vbp vbn x a1 a2 b
xmn4 vss a2 midn_a1a2_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn3 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 vss a1 midn_a1a2_b vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_a1a2_b b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp4 int_zn a1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp0 int_zn b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA21_2




.subckt SAEDRVT14_OA21_4 vdd vss vbp vbn x a1 a2 b
xmn4 vss a2 midn_a1a2_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 x int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn1 vss a1 midn_a1a2_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 midn_a1a2_b b int_zn vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp52 midp_a1_a22 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp42 int_zn a1 midp_a1_a22 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 int_zn a1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 x int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp0 int_zn b vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_OA21_4




.subckt SAEDRVT14_OA21B_1 vdd vss vbp vbn x a1 a2 b
xmn4 x b1ndb2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 b1ndb2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 b1ndb2 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 x b midp_a_b1ndb2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 midp_a_b1ndb2 b1ndb2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 b1ndb2 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_b1_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OA21B_1




.subckt SAEDRVT14_OA21B_2 vdd vss vbp vbn x a1 a2 b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 x1 b1ndb2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn3 x1 b vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 b1ndb2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 b1ndb2 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp42 x1 b midp_a_b1ndb22 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp32 midp_a_b1ndb22 b1ndb2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x1 b midp_a_b1ndb2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 midp_a_b1ndb2 b1ndb2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 b1ndb2 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_b1_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OA21B_2




.subckt SAEDRVT14_OA21B_4 vdd vss vbp vbn x a1 a2 b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 x1 b1ndb2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn3 x1 b vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn1 b1ndb2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 b1ndb2 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp44 x1 b midp_a_b1ndb24 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp43 x1 b midp_a_b1ndb23 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp42 x1 b midp_a_b1ndb22 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp34 midp_a_b1ndb24 b1ndb2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp33 midp_a_b1ndb23 b1ndb2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp32 midp_a_b1ndb22 b1ndb2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x1 b midp_a_b1ndb2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 midp_a_b1ndb2 b1ndb2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 b1ndb2 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 midp_b1_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OA21B_4




.subckt SAEDRVT14_OA21B_U_0P5 vdd vss vbp vbn x a1 a2 b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn4 x1 b1ndb2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 x1 b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 b1ndb2 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 b1ndb2 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 x1 b midp_a_b1ndb2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_a_b1ndb2 b1ndb2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 b1ndb2 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 midp_b1_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OA21B_U_0P5




.subckt SAEDRVT14_OA21_MM_1 vdd vss vbp vbn x a1 a2 b
xmn5 int_zn a2 midn_a1a2_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 int_zn a1 midn_a1a2_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn3 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_a1a2_b b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 int_zn a1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp4 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 int_zn b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA21_MM_1




.subckt SAEDRVT14_OA21_MM_2 vdd vss vbp vbn x a1 a2 b
xmn5 int_zn a2 midn_a1a2_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 int_zn a1 midn_a1a2_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn3 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 midn_a1a2_b b vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 int_zn a1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp4 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 int_zn b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA21_MM_2




.subckt SAEDRVT14_OA21_MM_4 vdd vss vbp vbn x a1 a2 b
xmn5 int_zn a2 midn_a1a2_b vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn4 int_zn a1 midn_a1a2_b vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn3 x int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn1 midn_a1a2_b b vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmp51 int_zn a1 midp_a1_a21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp41 midp_a1_a21 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 int_zn a1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp4 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 x int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 int_zn b vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_OA21_MM_4




.subckt SAEDRVT14_OA21_MM_6 vdd vss vbp vbn x a1 a2 b
xmn5 int_zn a2 midn_a1a2_b vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn4 int_zn a1 midn_a1a2_b vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn3 x int_zn vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmn1 midn_a1a2_b b vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp5 int_zn a1 midp_a1_a2 vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp4 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp3 x int_zn vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmp1 int_zn b vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_OA21_MM_6




.subckt SAEDRVT14_OA21_U_0P5 vdd vss vbp vbn x a1 a2 b
xmn4 vss a2 midn_a1a2_b vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn3 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 vss a1 midn_a1a2_b vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 midn_a1a2_b b int_zn vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp4 int_zn a1 midp_a1_a2 vbp p08_rev l=0.014u nf=2 m=1 nfin=2
xmp3 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 int_zn b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OA21_U_0P5




.subckt SAEDRVT14_OA22_0P75 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmn7 int_zn A1 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn6 int_zn A2 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn5 midn_a1a2_b1b2 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn4 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn1 midn_a1a2_b1b2 B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp8 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp7 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp6 midp_a1_a2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp5 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp4 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA22_0P75




.subckt SAEDRVT14_OA221_1 VDD VSS VBP VBN X A1 A2 B1 B2 C
Mxn9 midn_a1a2_b1b2 B2 midn_b1b2_c VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxn8 VSS A2 midn_a1a2_b1b2 VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxn7 VSS A1 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn6 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn1 midn_a1a2_b1b2 B1 midn_b1b2_c VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn0 midn_b1b2_c C int_zn VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxp10 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxp9 midp_a1_a2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxp8 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxp7 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp6 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxp3 int_zn C VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_OA221_1




.subckt SAEDRVT14_OA221_2 VDD VSS VBP VBN X A1 A2 B1 B2 C
Mxn9 midn_a1a2_b1b2 B2 midn_b1b2_c VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxn8 VSS A2 midn_a1a2_b1b2 VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxn7 VSS A1 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxn6 X int_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxn1 midn_a1a2_b1b2 B1 midn_b1b2_c VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxn0 midn_b1b2_c C int_zn VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxp10 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp9 midp_a1_a2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp8 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxp7 X int_zn VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxp6 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp3 int_zn C VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_OA221_2




.subckt SAEDRVT14_OA221_4 VDD VSS VBP VBN X A1 A2 B1 B2 C
Mxn9 midn_a1a2_b1b2 B2 midn_b1b2_c VBN n08 l=0.014u nf=2 m=2 nfin=4
Mxn8 VSS A2 midn_a1a2_b1b2 VBN n08 l=0.014u nf=2 m=2 nfin=4
Mxn7 VSS A1 midn_a1a2_b1b2 VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxn6 X int_zn VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxn1 midn_a1a2_b1b2 B1 midn_b1b2_c VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxn0 midn_b1b2_c C int_zn VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxp102 int_zn A1 midp_a1_a22 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp92 midp_a1_a22 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp82 midp_b1_b22 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp62 int_zn B1 midp_b1_b22 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp10 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp9 midp_a1_a2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp8 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp7 X int_zn VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxp6 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxp3 int_zn C VDD VBP p08 l=0.014u nf=2 m=2 nfin=4
.ends SAEDRVT14_OA221_4




.subckt SAEDRVT14_OA22_1 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmn7 int_zn A1 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn6 int_zn A2 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn5 midn_a1a2_b1b2 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn4 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn1 midn_a1a2_b1b2 B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp8 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp7 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp6 midp_a1_a2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp5 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp4 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA22_1




.subckt SAEDRVT14_OA221_U_0P5 VDD VSS VBP VBN X A1 A2 B1 B2 C
Mxn9 midn_a1a2_b1b2 B2 midn_b1b2_c VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn8 VSS A2 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn7 VSS A1 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn6 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxn1 midn_a1a2_b1b2 B1 midn_b1b2_c VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn0 midn_b1b2_c C int_zn VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxp10 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxp9 midp_a1_a2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxp8 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxp7 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxp6 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxp3 int_zn C VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OA221_U_0P5




.subckt SAEDRVT14_OA222_1 VDD VSS VBP VBN X A1 A2 B1 B2 C1 C2
Mxn13 midn_b1b2_c1c2 C2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxn12 midn_a1a2_b1b2 B2 midn_b1b2_c1c2 VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxn11 int_zn A2 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn10 int_zn A1 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxn9 midn_a1a2_b1b2 B1 midn_b1b2_c1c2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn8 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn1 midn_b1b2_c1c2 C1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxp13 midp_c1_c2 C2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp12 int_zn C1 midp_c1_c2 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp11 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxp10 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxp9 midp_a1_a2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxp8 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp6 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OA222_1




.subckt SAEDRVT14_OA222_2 VDD VSS VBP VBN X A1 A2 B1 B2 C1 C2
Mxn13 midn_b1b2_c1c2 C2 VSS VBN n08 l=0.014u nf=5 m=1 nfin=2
Mxn12 midn_a1a2_b1b2 B2 midn_b1b2_c1c2 VBN n08 l=0.014u nf=3 m=1 nfin=3
Mxn11 int_zn A2 midn_a1a2_b1b2 VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxn10 int_zn A1 midn_a1a2_b1b2 VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxn9 midn_a1a2_b1b2 B1 midn_b1b2_c1c2 VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxn8 X int_zn VSS VBN n08 l=0.014u nf=3 m=1 nfin=3
Mxn1 midn_b1b2_c1c2 C1 VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxp13 midp_c1_c2 C2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxp12 int_zn C1 midp_c1_c2 VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxp11 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxp10 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxp9 midp_a1_a2 A2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=2
Mxp8 X int_zn VDD VBP p08 l=0.014u nf=3 m=1 nfin=4
Mxp6 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_OA222_2




.subckt SAEDRVT14_OA222_4 VDD VSS VBP VBN X A1 A2 B1 B2 C1 C2
Mxn13 midn_b1b2_c1c2 C2 VSS VBN n08 l=0.014u nf=5 m=1 nfin=4
Mxn12 midn_a1a2_b1b2 B2 midn_b1b2_c1c2 VBN n08 l=0.014u nf=5 m=1 nfin=4
Mxn11 int_zn A2 midn_a1a2_b1b2 VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxn10 int_zn A1 midn_a1a2_b1b2 VBN n08 l=0.014u nf=4 m=1 nfin=2
Mxn9 midn_a1a2_b1b2 B1 midn_b1b2_c1c2 VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxn8 X int_zn VSS VBN n08 l=0.014u nf=8 m=1 nfin=3
Mxn1 midn_b1b2_c1c2 C1 VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxp13 midp_c1_c2 C2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxp12 int_zn C1 midp_c1_c2 VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxp11 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxp10 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxp9 midp_a1_a2 A2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=2
Mxp8 X int_zn VDD VBP p08 l=0.014u nf=8 m=1 nfin=4
Mxp6 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=4 m=1 nfin=2
.ends SAEDRVT14_OA222_4




.subckt SAEDRVT14_OA22_2 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmn7 int_zn A1 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn6 int_zn A2 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn5 midn_a1a2_b1b2 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn4 X int_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn1 midn_a1a2_b1b2 B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp8 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp7 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp6 midp_a1_a2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp5 X int_zn VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp4 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA22_2




.subckt SAEDRVT14_OA222_U_0P5 VDD VSS VBP VBN X A1 A2 B1 B2 C1 C2
Mxn13 midn_b1b2_c1c2 C2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxn12 midn_a1a2_b1b2 B2 midn_b1b2_c1c2 VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxn11 int_zn A2 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn10 int_zn A1 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxn9 midn_a1a2_b1b2 B1 midn_b1b2_c1c2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn8 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxn1 midn_b1b2_c1c2 C1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxp13 midp_c1_c2 C2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp12 int_zn C1 midp_c1_c2 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp11 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxp10 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxp9 midp_a1_a2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxp8 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxp6 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OA222_U_0P5




.subckt SAEDRVT14_OA22_4 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmn7 int_zn A1 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn6 int_zn A2 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn5 midn_a1a2_b1b2 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn4 X int_zn VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmn1 midn_a1a2_b1b2 B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp8 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp7 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp6 midp_a1_a2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp5 X int_zn VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxmp4 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA22_4




.subckt SAEDRVT14_OA22_U_0P5 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmn7 int_zn A1 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn6 int_zn A2 midn_a1a2_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn5 midn_a1a2_b1b2 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn4 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn1 midn_a1a2_b1b2 B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp8 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp7 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp6 midp_a1_a2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp5 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp4 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OA22_U_0P5




.subckt SAEDRVT14_OA2BB2_0P5 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmn8 X int_zn yn VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn7 yn int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn6 int_zn x1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn5 midn_a1_a2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn4 x1 b1ndb2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn3 x1 A1 midn_a1_a2 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn1 b1ndb2 B2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn0 b1ndb2 B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmp8 X int_zn yp VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp7 yp int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp6 int_zn x1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp5 x1 A2 midp_a1a2_b1ndb2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp3 x1 A1 midp_a1a2_b1ndb2 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp2 midp_a1a2_b1ndb2 b1ndb2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp1 b1ndb2 B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_OA2BB2_0P5




.subckt SAEDRVT14_OA2BB2_1 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmn8 X int_zn yn VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn7 yn int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn6 int_zn x1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn5 midn_a1_a2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn4 x1 b1ndb2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn3 x1 A1 midn_a1_a2 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn1 b1ndb2 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 b1ndb2 B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmp8 X int_zn yp VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp7 yp int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp6 int_zn x1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp5 x1 A2 midp_a1a2_b1ndb2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp3 x1 A1 midp_a1a2_b1ndb2 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp2 midp_a1a2_b1ndb2 b1ndb2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp1 b1ndb2 B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OA2BB2_1




.subckt SAEDRVT14_OA2BB2_2 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmn8 X int_zn yn VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn7 yn int_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn6 int_zn x1 VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmn5 midn_a1_a2 A2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmn4 x1 b1ndb2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmn3 x1 A1 midn_a1_a2 VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmn1 b1ndb2 B2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmn0 b1ndb2 B1 VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmp8 X int_zn yp VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp7 yp int_zn VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp6 int_zn x1 VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp5 x1 A2 midp_a1a2_b1ndb2 VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp3 x1 A1 midp_a1a2_b1ndb2 VBP p08 l=0.014u nf=2 m=1 nfin=2
Mxmp2 midp_a1a2_b1ndb2 b1ndb2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=2
Mxmp1 b1ndb2 B1 midp_b1_b2 VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp0 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_OA2BB2_2




.subckt SAEDRVT14_OA2BB2_4 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmn8 X int_zn yn VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmn7 yn int_zn VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmn6 int_zn x1 VSS VBN n08 l=0.014u nf=4 m=1 nfin=2
Mxmn5 midn_a1_a2 A2 VSS VBN n08 l=0.014u nf=4 m=1 nfin=2
Mxmn4 x1 b1ndb2 VSS VBN n08 l=0.014u nf=4 m=1 nfin=2
Mxmn3 x1 A1 midn_a1_a2 VBN n08 l=0.014u nf=4 m=1 nfin=2
Mxmn1 b1ndb2 B2 VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmn0 b1ndb2 B1 VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmp8 X int_zn yp VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp7 yp int_zn VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxmp6 int_zn x1 VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxmp5 x1 A2 midp_a1a2_b1ndb2 VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxmp3 x1 A1 midp_a1a2_b1ndb2 VBP p08 l=0.014u nf=4 m=1 nfin=2
Mxmp2 midp_a1a2_b1ndb2 b1ndb2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=2
Mxmp1 b1ndb2 B1 midp_b1_b2 VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxmp0 midp_b1_b2 B2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_OA2BB2_4




.subckt SAEDRVT14_OA2BB2_V1_0P5 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmp5 net13 A2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=2
Mxmp4 net13 A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp3 X net15 net13 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp1 net16 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmn0 net15 B1 net16 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmn5 net15 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn4 net15 B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn3 X net15 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn2 X A1 midn_a1a2 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn1 midn_a1a2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OA2BB2_V1_0P5




.subckt SAEDRVT14_OA2BB2_V1_0P75 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmp5 net13 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp4 net13 A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp3 X net15 net13 VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp1 net16 B2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmn0 net15 B1 net16 VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmn5 net15 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn4 net15 B1 VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn3 X net15 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn2 X A1 midn_a1a2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn1 midn_a1a2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA2BB2_V1_0P75




.subckt SAEDRVT14_OA2BB2_V1_1 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmp5 net13 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp4 net13 A1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp3 X net15 net13 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 net16 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 net15 B1 net16 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmn5 net15 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn4 net15 B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn3 X net15 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn2 X A1 midn_a1a2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn1 midn_a1a2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OA2BB2_V1_1




.subckt SAEDRVT14_OA2BB2_V1_2 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmp5 net13 A2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp4 net13 A1 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp3 X net15 net13 VBP p08 l=0.014u nf=6 m=1 nfin=4
Mxmp1 net16 B2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmn0 net15 B1 net16 VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmn22 X A1 midn_a1a22 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn12 midn_a1a22 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn5 net15 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn4 net15 B1 VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmn3 X net15 VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmn2 X A1 midn_a1a2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn1 midn_a1a2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OA2BB2_V1_2




.subckt SAEDRVT14_OA2BB2_V1_4 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmp5 net13 A2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp4 net13 A1 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp3 X net15 net13 VBP p08 l=0.014u nf=8 m=1 nfin=4
Mxmp1 net16 B2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmn0 net15 B1 net16 VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmn5 net15 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn4 net15 B1 VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmn3 X net15 VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmn2 X A1 midn_a1a2 VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmn1 midn_a1a2 A2 VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_OA2BB2_V1_4




.subckt SAEDRVT14_OA31_1P5 VDD VSS VBP VBN X A1 A2 A3 B
Mxmn6 midn_a_b1b2b3 A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn5 midn_a_b1b2b3 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn4 X int_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn1 midn_a_b1b2b3 A1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 int_zn B midn_a_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmp7 midp_b2_b3 A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp6 int_zn B VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp5 X int_zn VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp4 midp_b1_b2 A2 midp_b2_b3 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp1 int_zn A1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA31_1P5




.subckt SAEDRVT14_OA31_1 VDD VSS VBP VBN X A1 A2 A3 B
Mxmn6 midn_a_b1b2b3 A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn5 midn_a_b1b2b3 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn4 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn1 midn_a_b1b2b3 A1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 int_zn B midn_a_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmp7 midp_b2_b3 A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp6 int_zn B VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp5 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp4 midp_b1_b2 A2 midp_b2_b3 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp1 int_zn A1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA31_1




.subckt SAEDRVT14_OA31_2 VDD VSS VBP VBN X A1 A2 A3 B
Mxmn6 midn_a_b1b2b3 A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn5 midn_a_b1b2b3 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn4 X int_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmn1 midn_a_b1b2b3 A1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 int_zn B midn_a_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmp7 midp_b2_b3 A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp6 int_zn B VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp5 X int_zn VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp4 midp_b1_b2 A2 midp_b2_b3 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp1 int_zn A1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA31_2




.subckt SAEDRVT14_OA31_4 VDD VSS VBP VBN X A1 A2 A3 B
Mxmn6 midn_a_b1b2b3 A3 VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn5 midn_a_b1b2b3 A2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn4 X int_zn VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmn1 midn_a_b1b2b3 A1 VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn0 int_zn B midn_a_b1b2b3 VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmp42 midp_b1_b22 A2 midp_b2_b3 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp12 int_zn A1 midp_b1_b22 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp7 midp_b2_b3 A3 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp6 int_zn B VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp5 X int_zn VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxmp4 midp_b1_b2 A2 midp_b2_b3 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 int_zn A1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OA31_4




.subckt SAEDRVT14_OA31_U_0P5 VDD VSS VBP VBN X A1 A2 A3 B
Mxmn6 midn_a_b1b2b3 A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn5 midn_a_b1b2b3 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn4 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn1 midn_a_b1b2b3 A1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn0 int_zn B midn_a_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp7 midp_b2_b3 A3 VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp6 int_zn B VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp5 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp4 midp_b1_b2 A2 midp_b2_b3 VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp1 int_zn A1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OA31_U_0P5




.subckt SAEDRVT14_OA32_0P75 VDD VSS VBP VBN X A1 A2 A3 B1 B2
Mxmn9 int_zn B1 midn_a1a2_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn8 int_zn B2 midn_a1a2_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn7 midn_a1a2_b1b2b3 A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn6 midn_a1a2_b1b2b3 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn5 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn1 midn_a1a2_b1b2b3 A1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp10 midp_b2_b3 A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp9 midp_a1_a2 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp8 midp_b1_b2 A2 midp_b2_b3 VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp7 int_zn A1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp6 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp4 int_zn B1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA32_0P75




.subckt SAEDRVT14_OA32_1 VDD VSS VBP VBN X A1 A2 A3 B1 B2
Mxmn9 int_zn B1 midn_a1a2_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn8 int_zn B2 midn_a1a2_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn7 midn_a1a2_b1b2b3 A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn6 midn_a1a2_b1b2b3 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn5 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn1 midn_a1a2_b1b2b3 A1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp10 midp_b2_b3 A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp9 midp_a1_a2 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp8 midp_b1_b2 A2 midp_b2_b3 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp7 int_zn A1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp6 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp4 int_zn B1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OA32_1




.subckt SAEDRVT14_OA32_2 VDD VSS VBP VBN X A1 A2 A3 B1 B2
Mxmn9 int_zn B1 midn_a1a2_b1b2b3 VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn8 int_zn B2 midn_a1a2_b1b2b3 VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmn7 midn_a1a2_b1b2b3 A3 VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn6 midn_a1a2_b1b2b3 A2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn5 X int_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmn1 midn_a1a2_b1b2b3 A1 VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmp10 midp_b2_b3 A3 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp9 midp_a1_a2 B2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=2
Mxmp8 midp_b1_b2 A2 midp_b2_b3 VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp7 int_zn A1 midp_b1_b2 VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp6 X int_zn VDD VBP p08 l=0.014u nf=2 m=1 nfin=2
Mxmp4 int_zn B1 midp_a1_a2 VBP p08 l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_OA32_2




.subckt SAEDRVT14_OA32_4 VDD VSS VBP VBN X A1 A2 A3 B1 B2
Mxmn9 int_zn B1 midn_a1a2_b1b2b3 VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmn8 int_zn B2 midn_a1a2_b1b2b3 VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmn7 midn_a1a2_b1b2b3 A3 VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmn6 midn_a1a2_b1b2b3 A2 VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmn5 X int_zn VSS VBN n08 l=0.014u nf=4 m=1 nfin=2
Mxmn1 midn_a1a2_b1b2b3 A1 VSS VBN n08 l=0.014u nf=4 m=1 nfin=2
Mxmp10 midp_b2_b3 A3 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp9 midp_a1_a2 B2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxmp8 midp_b1_b2 A2 midp_b2_b3 VBP p08 l=0.014u nf=5 m=1 nfin=4
Mxmp7 int_zn A1 midp_b1_b2 VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp6 X int_zn VDD VBP p08 l=0.014u nf=4 m=1 nfin=2
Mxmp4 int_zn B1 midp_a1_a2 VBP p08 l=0.014u nf=4 m=1 nfin=3
.ends SAEDRVT14_OA32_4




.subckt SAEDRVT14_OA32_U_0P5 VDD VSS VBP VBN X A1 A2 A3 B1 B2
Mxmn9 int_zn B1 midn_a1a2_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn8 int_zn B2 midn_a1a2_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn7 midn_a1a2_b1b2b3 A3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn6 midn_a1a2_b1b2b3 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn5 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn1 midn_a1a2_b1b2b3 A1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp10 midp_b2_b3 A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp9 midp_a1_a2 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp8 midp_b1_b2 A2 midp_b2_b3 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp7 int_zn A1 midp_b1_b2 VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp6 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp4 int_zn B1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA32_U_0P5




.subckt SAEDRVT14_OA33_1 VDD VSS VBP VBN X A1 A2 A3 B1 B2 B3
Mxmmn18 midn_a1a2a3_b1b2b3 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmmn17 midn_a1a2a3_b1b2b3 B3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmmn16 int_zn A3 midn_a1a2a3_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmmn15 int_zn A2 midn_a1a2a3_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmmn14 int_zn A1 midn_a1a2a3_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmmn8 midn_a1a2a3_b1b2b3 B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmmn7 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmmp17 midp_b2_b3 B3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp16 midp_a2_a3 A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmmp15 midp_a1_a2 A2 midp_a2_a3 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp14 midp_b1_b2 B2 midp_b2_b3 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp13 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp12 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmmp6 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OA33_1




.subckt SAEDRVT14_OA33_2 VDD VSS VBP VBN X A1 A2 A3 B1 B2 B3
Mxmmn18 midn_a1a2a3_b1b2b3 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmmn17 midn_a1a2a3_b1b2b3 B3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmmn16 int_zn A3 midn_a1a2a3_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmmn15 int_zn A2 midn_a1a2a3_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmmn14 int_zn A1 midn_a1a2a3_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmmn8 midn_a1a2a3_b1b2b3 B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmmn7 X int_zn VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmmp17 midp_b2_b3 B3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp16 midp_a2_a3 A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmmp15 midp_a1_a2 A2 midp_a2_a3 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp14 midp_b1_b2 B2 midp_b2_b3 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp13 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp12 X int_zn VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmmp6 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OA33_2




.subckt SAEDRVT14_OA33_4 VDD VSS VBP VBN X A1 A2 A3 B1 B2 B3
Mxmnbuf2 X d1g2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmnbuf1 d1g2 x1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmmn18 midn_a1a2a3_b1b2b3 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmmn17 midn_a1a2a3_b1b2b3 B3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmmn16 int_zn A3 midn_a1a2a3_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmmn15 int_zn A2 midn_a1a2a3_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmmn14 int_zn A1 midn_a1a2a3_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmmn8 midn_a1a2a3_b1b2b3 B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmmn7 x1 int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmpbuf2 X d1g2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmpbuf1 d1g2 x1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp17 midp_b2_b3 B3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp16 midp_a2_a3 A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmmp15 midp_a1_a2 A2 midp_a2_a3 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp14 midp_b1_b2 B2 midp_b2_b3 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp13 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmmp12 x1 int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmmp6 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OA33_4




.subckt SAEDRVT14_OA33_U_0P5 VDD VSS VBP VBN X A1 A2 A3 B1 B2 B3
Mxmn11 midn_a1a2a3_b1b2b3 B2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn10 midn_a1a2a3_b1b2b3 B3 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn9 int_zn A3 midn_a1a2a3_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn8 int_zn A2 midn_a1a2a3_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn7 int_zn A1 midn_a1a2a3_b1b2b3 VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn6 X int_zn VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmn1 midn_a1a2a3_b1b2b3 B1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmp12 int_zn B1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp11 midp_b1_b2 B2 midp_b2_b3 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp10 midp_b2_b3 B3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp9 midp_a2_a3 A3 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp8 midp_a1_a2 A2 midp_a2_a3 VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp7 X int_zn VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp4 int_zn A1 midp_a1_a2 VBP p08 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OA33_U_0P5




.subckt SAEDRVT14_OAI21_0P5 VDD VSS VBP VBN X A1 A2 B
Mxmn2 X B midn_a_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn1 midn_a_b1b2 A1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 midn_a_b1b2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp2 midp_b1_b2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 X A1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp0 X B VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI21_0P5




.subckt SAEDRVT14_OAI21_0P75 VDD VSS VBP VBN X A1 A2 B
Mxmn2 X B midn_a_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn1 midn_a_b1b2 A1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 midn_a_b1b2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmp2 midp_b1_b2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 X A1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp0 X B VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI21_0P75




.subckt SAEDRVT14_OAI211_0P5 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmnbuf2 X d1g2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmnbuf1 d1g2 x1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn3 midn_a_b B2 midn_b_c1c2 VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn2 x1 B1 midn_a_b VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn1 midn_b_c1c2 A1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=3
Mxmn0 midn_b_c1c2 A2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmpbuf2 X d1g2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmpbuf1 d1g2 x1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp3 x1 B1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmp2 midp_c1_c2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp1 x1 A1 midp_c1_c2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 x1 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI211_0P5




.subckt SAEDRVT14_OAI211_1 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmnbuf2 X d1g2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=2
Mxmnbuf1 d1g2 x1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 midn_a_b B2 midn_b_c1c2 VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn2 x1 B1 midn_a_b VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmn1 midn_b_c1c2 A1 VSS VBN n08 l=0.014u nf=2 m=1 nfin=2
Mxmn0 midn_b_c1c2 A2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmpbuf2 X d1g2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
Mxmpbuf1 d1g2 x1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp3 x1 B1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp2 midp_c1_c2 A2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp1 x1 A1 midp_c1_c2 VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp0 x1 B2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OAI211_1




.subckt SAEDRVT14_OAI211_2 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmnbuf2 X d1g2 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmnbuf1 d1g2 x1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 midn_a_b B2 midn_b_c1c2 VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmn2 x1 B1 midn_a_b VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmn1 midn_b_c1c2 A1 VSS VBN n08 l=0.014u nf=4 m=1 nfin=2
Mxmn0 midn_b_c1c2 A2 VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmpbuf2 X d1g2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmpbuf1 d1g2 x1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp3 x1 B1 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmp2 midp_c1_c2 A2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp1 x1 A1 midp_c1_c2 VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxmp0 x1 B2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_OAI211_2




.subckt SAEDRVT14_OAI211_4 VDD VSS VBP VBN X A1 A2 B1 B2
Mxmnbuf2 X d1g2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmnbuf1 d1g2 x1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn3 midn_a_b B2 midn_b_c1c2 VBN n08 l=0.014u nf=8 m=1 nfin=3
Mxmn2 x1 B1 midn_a_b VBN n08 l=0.014u nf=8 m=1 nfin=4
Mxmn1 midn_b_c1c2 A1 VSS VBN n08 l=0.014u nf=8 m=1 nfin=2
Mxmn0 midn_b_c1c2 A2 VSS VBN n08 l=0.014u nf=8 m=1 nfin=4
Mxmpbuf2 X d1g2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=4
Mxmpbuf1 d1g2 x1 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp3 x1 B1 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp2 midp_c1_c2 A2 VDD VBP p08 l=0.014u nf=8 m=1 nfin=4
Mxmp1 x1 A1 midp_c1_c2 VBP p08 l=0.014u nf=8 m=1 nfin=3
Mxmp0 x1 B2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_OAI211_4




.subckt SAEDRVT14_OAI21_1P5 VDD VSS VBP VBN X A1 A2 B
Mxmn2 X B midn_a_b1b2 VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn1 midn_a_b1b2 A1 VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn0 midn_a_b1b2 A2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmp22 midp_b1_b22 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp12 X A1 midp_b1_b22 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp2 midp_b1_b2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp1 X A1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp0 X B VDD VBP p08 l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_OAI21_1P5




.subckt SAEDRVT14_OAI21_1 VDD VSS VBP VBN X A1 A2 B
Mxmn2 X B midn_a_b1b2 VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn1 midn_a_b1b2 A1 VSS VBN n08 l=0.014u nf=1 m=1 nfin=4
Mxmn0 midn_a_b1b2 A2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmp2 midp_b1_b2 A2 VDD VBP p08 l=0.014u nf=2 m=1 nfin=3
Mxmp1 X A1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp0 X B VDD VBP p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI21_1




.subckt SAEDRVT14_OAI21_2 VDD VSS VBP VBN X A1 A2 B
Mxmn2 X B midn_a_b1b2 VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn1 midn_a_b1b2 A1 VSS VBN n08 l=0.014u nf=2 m=1 nfin=3
Mxmn0 midn_a_b1b2 A2 VSS VBN n08 l=0.014u nf=2 m=1 nfin=4
Mxmp22 midp_b1_b22 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp12 X A1 midp_b1_b22 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp2 midp_b1_b2 A2 VDD VBP p08 l=0.014u nf=1 m=1 nfin=4
Mxmp1 X A1 midp_b1_b2 VBP p08 l=0.014u nf=1 m=1 nfin=3
Mxmp0 X B VDD VBP p08 l=0.014u nf=2 m=1 nfin=2
.ends SAEDRVT14_OAI21_2




.subckt SAEDRVT14_OAI21_3 VDD VSS VBP VBN X A1 A2 B
Mxmn2 X B midn_a_b1b2 VBN n08 l=0.014u nf=3 m=1 nfin=3
Mxmn1 midn_a_b1b2 A1 VSS VBN n08 l=0.014u nf=3 m=1 nfin=3
Mxmn0 midn_a_b1b2 A2 VSS VBN n08 l=0.014u nf=3 m=1 nfin=4
Mxmp2 midp_b1_b2 A2 VDD VBP p08 l=0.014u nf=3 m=1 nfin=4
Mxmp1 X A1 midp_b1_b2 VBP p08 l=0.014u nf=3 m=1 nfin=3
Mxmp0 X B VDD VBP p08 l=0.014u nf=3 m=1 nfin=2
.ends SAEDRVT14_OAI21_3




.subckt SAEDRVT14_OAI21_4 VDD VSS VBP VBN X A1 A2 B
Mxmn2 X B midn_a_b1b2 VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmn1 midn_a_b1b2 A1 VSS VBN n08 l=0.014u nf=4 m=1 nfin=3
Mxmn0 midn_a_b1b2 A2 VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmp2 midp_b1_b2 A2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp1 X A1 midp_b1_b2 VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxmp0 X B VDD VBP p08 l=0.014u nf=4 m=1 nfin=2
.ends SAEDRVT14_OAI21_4




.subckt SAEDRVT14_OAI21_V1_4 VDD VSS VBP VBN X A1 A2 B
Mxmn2 midn_a_b1b2 B VSS VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmn1 X A1 midn_a_b1b2 VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmn0 X A2 midn_a_b1b2 VBN n08 l=0.014u nf=4 m=1 nfin=4
Mxmp2 midp_b1_b2 A2 VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
Mxmp1 X A1 midp_b1_b2 VBP p08 l=0.014u nf=4 m=1 nfin=4
Mxmp0 X B VDD VBP p08 l=0.014u nf=4 m=1 nfin=3
.ends SAEDRVT14_OAI21_V1_4




.subckt SAEDRVT14_OAI21_V1_6 VDD VSS VBP VBN X A1 A2 B
Mxmn2 midn_a_b1b2 B VSS VBN n08 l=0.014u nf=6 m=1 nfin=4
Mxmn1 X A1 midn_a_b1b2 VBN n08 l=0.014u nf=6 m=1 nfin=4
Mxmn0 X A2 midn_a_b1b2 VBN n08 l=0.014u nf=6 m=1 nfin=4
Mxmp2 midp_b1_b2 A2 VDD VBP p08 l=0.014u nf=6 m=1 nfin=4
Mxmp1 X A1 midp_b1_b2 VBP p08 l=0.014u nf=6 m=1 nfin=4
Mxmp0 X B VDD VBP p08 l=0.014u nf=6 m=1 nfin=3
.ends SAEDRVT14_OAI21_V1_6




.subckt SAEDRVT14_OAI21_V1_8 VDD VSS VBP VBN X A1 A2 B
Mxmn2 midn_a_b1b2 B VSS VBN n08 l=0.014u nf=8 m=1 nfin=4
Mxmn1 X A1 midn_a_b1b2 VBN n08 l=0.014u nf=8 m=1 nfin=4
Mxmn0 X A2 midn_a_b1b2 VBN n08 l=0.014u nf=8 m=1 nfin=4
Mxmp2 midp_b1_b2 A2 VDD VBP p08 l=0.014u nf=8 m=1 nfin=4
Mxmp1 X A1 midp_b1_b2 VBP p08 l=0.014u nf=8 m=1 nfin=4
Mxmp0 X B VDD VBP p08 l=0.014u nf=8 m=1 nfin=3
.ends SAEDRVT14_OAI21_V1_8




.subckt SAEDRVT14_OAI22_0P5 vdd vss vbp vbn x a1 a2 b1 b2
xmn3 x a1 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x a2 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 midn_a1a2_b1b2 b1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_a1a2_b1b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 x a1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_b1_b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 x b1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI22_0P5





.subckt SAEDRVT14_SRRDPQ_1 ck d nrestore q qn save vdd vddr vss
xm13 net8 net1556 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn15 jk jk2 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm0 net28 nrestore _n766 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn21 netn102 saven vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn20 jk2 jk netn102 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn19 netn10 restore vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn18 _n766 jk netn10 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn22 saven save vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn32 netn103 save vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn33 jk2 net8 netn103 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn26 restore nrestore vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm5 net2 ckn vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm7 net1556 net8 net2 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn03 hjf d vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm11 net29 net28 net7 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn13 q net8 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm3 net28 net29 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm12 net7 ckp vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm15 qn net1556 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn011 ckn ck vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn1 net29 ckn hjf vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn012 ckp ckn vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn7 net1556 ckp _n766 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp11 net28 restore _n766 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp15 jk jk2 vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp19 _n766 jk netp10 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp18 netp10 nrestore vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp1 net29 ckp hjf vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp7 net1556 ckn _n766 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp21 jk2 jk netp102 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp26 restore nrestore vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp22 saven save vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp33 jk2 net8 netp103 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm17 qn net1556 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm4 net3 ckp vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm6 net1556 net8 net3 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm1 netp102 save vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm8 netp103 saven vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp03 hjf d vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm18 q net8 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm9 net29 net28 net9 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp011 ckn ck vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm10 net9 ckn vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp012 ckp ckn vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm14 net8 net1556 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm2 net28 net29 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
.ends SAEDRVT14_SRRDPQ_1




.subckt SAEDRVT14_OAI221_0P5 vdd vss vbp vbn x a1 a2 b1 b2 c
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 midn_a_b1b2 a1 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 midn_a_b1b2 a2 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x1 c midn_a_b1b2 vbn n08_rev l=0.014u nf=4 m=1 nfin=2
xmn1 midn_b1b2_c1c2 b1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_b1b2_c1c2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 midp_b1_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 x1 c vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_c1_c2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 x1 b1 midp_c1_c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI221_0P5




.subckt SAEDRVT14_OAI221_1 vdd vss vbp vbn x a1 a2 b1 b2 c
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 midn_a_b1b2 a1 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 midn_a_b1b2 a2 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 x1 c midn_a_b1b2 vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn1 midn_b1b2_c1c2 b1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 midn_b1b2_c1c2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 midp_b1_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 x1 c vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 midp_c1_c2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 b1 midp_c1_c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OAI221_1




.subckt SAEDRVT14_OAI221_2 vdd vss vbp vbn x a1 a2 b1 b2 c
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 midn_a_b1b2 a1 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn4 midn_a_b1b2 a2 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn2 x1 c midn_a_b1b2 vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 midn_b1b2_c1c2 b1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn0 midn_b1b2_c1c2 b2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp52 x1 a1 midp_b1_b22 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp42 midp_b1_b22 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp22 midp_c1_c22 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp12 x1 b1 midp_c1_c22 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp5 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 midp_b1_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 x1 c vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 midp_c1_c2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 b1 midp_c1_c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OAI221_2




.subckt SAEDRVT14_OAI221_4 vdd vss vbp vbn x a1 a2 b1 b2 c
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn5 midn_a_b1b2 a1 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn4 midn_a_b1b2 a2 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn2 x1 c midn_a_b1b2 vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn1 midn_b1b2_c1c2 b1 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn0 midn_b1b2_c1c2 b2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=5 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp54 x1 a1 midp_b1_b24 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp53 x1 a1 midp_b1_b23 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp52 x1 a1 midp_b1_b22 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp44 midp_b1_b24 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp43 midp_b1_b23 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp42 midp_b1_b22 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp24 midp_c1_c24 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp23 midp_c1_c23 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp22 midp_c1_c22 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp14 x1 b1 midp_c1_c24 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp13 x1 b1 midp_c1_c23 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp12 x1 b1 midp_c1_c22 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp5 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 midp_b1_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 x1 c vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp2 midp_c1_c2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 b1 midp_c1_c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OAI221_4




.subckt SAEDRVT14_OAI22_1P5 vdd vss vbp vbn x a1 a2 b1 b2
xmn3 x a1 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn2 x a2 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn1 midn_a1a2_b1b2 b1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn0 midn_a1a2_b1b2 b2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmp21 midp_b1_b21 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp11 x b1 midp_b1_b21 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x a1 midp_a1_a2 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp3 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp2 midp_b1_b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x b1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OAI22_1P5




.subckt SAEDRVT14_OAI22_1 vdd vss vbp vbn x a1 a2 b1 b2
xmn3 x a1 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 x a2 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_a1a2_b1b2 b1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 midn_a1a2_b1b2 b2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x a1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 midp_b1_b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x b1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OAI22_1




.subckt SAEDRVT14_OAI222_0P5 vdd vss vbp vbn x a1 a2 b1 b2 c1 c2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn7 x1 a2 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn6 x1 a1 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn5 midn_a1a2_b1b2 b1 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn4 midn_a1a2_b1b2 b2 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 midn_b1b2_c1c2 c1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_b1b2_c1c2 c2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp7 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 x1 a1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 x1 b1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp4 midp_b1_b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_c1_c2 c2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x1 c1 midp_c1_c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OAI222_0P5




.subckt SAEDRVT14_OAI222_1 vdd vss vbp vbn x a1 a2 b1 b2 c1 c2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn7 x1 a2 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn6 x1 a1 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn5 midn_a1a2_b1b2 b1 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn4 midn_a1a2_b1b2 b2 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 midn_b1b2_c1c2 c1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_b1b2_c1c2 c2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp7 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 x1 a1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 x1 b1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp4 midp_b1_b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_c1_c2 c2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x1 c1 midp_c1_c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OAI222_1




.subckt SAEDRVT14_OAI222_2 vdd vss vbp vbn x a1 a2 b1 b2 c1 c2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn7 x1 a2 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn6 x1 a1 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn5 midn_a1a2_b1b2 b1 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn4 midn_a1a2_b1b2 b2 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 midn_b1b2_c1c2 c1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_b1b2_c1c2 c2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp7 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 x1 a1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 x1 b1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp4 midp_b1_b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_c1_c2 c2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x1 c1 midp_c1_c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OAI222_2




.subckt SAEDRVT14_OAI222_4 vdd vss vbp vbn x a1 a2 b1 b2 c1 c2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn7 x1 a2 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn6 x1 a1 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn5 midn_a1a2_b1b2 b1 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn4 midn_a1a2_b1b2 b2 midn_b1b2_c1c2 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 midn_b1b2_c1c2 c1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_b1b2_c1c2 c2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp7 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp6 x1 a1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp5 x1 b1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp4 midp_b1_b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_c1_c2 c2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x1 c1 midp_c1_c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OAI222_4




.subckt SAEDRVT14_OAI22_2 vdd vss vbp vbn x a1 a2 b1 b2
xmn3 x a1 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn2 x a2 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn1 midn_a1a2_b1b2 b1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn0 midn_a1a2_b1b2 b2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmp21 midp_b1_b21 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp11 x b1 midp_b1_b21 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp4 x a1 midp_a1_a2 vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp3 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmp2 midp_b1_b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x b1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OAI22_2




.subckt SAEDRVT14_OAI22_3 vdd vss vbp vbn x a1 a2 b1 b2
xmn3 x a1 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn2 x a2 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn1 midn_a1a2_b1b2 b1 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn0 midn_a1a2_b1b2 b2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmp4 x a1 midp_a1_a2 vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp3 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp2 midp_b1_b2 b2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 x b1 midp_b1_b2 vbp p08_rev l=0.014u nf=3 m=1 nfin=4
.ends SAEDRVT14_OAI22_3




.subckt SAEDRVT14_OAI22_4 vdd vss vbp vbn x a1 a2 b1 b2
xmn3 x a1 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn2 x a2 midn_a1a2_b1b2 vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn1 midn_a1a2_b1b2 b1 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn0 midn_a1a2_b1b2 b2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp23 midp_b1_b23 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp22 midp_b1_b22 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp21 midp_b1_b21 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp13 x b1 midp_b1_b23 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp12 x b1 midp_b1_b22 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp11 x b1 midp_b1_b21 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x a1 midp_a1_a2 vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp3 midp_a1_a2 a2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp2 midp_b1_b2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x b1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OAI22_4




.subckt SAEDRVT14_OAI31_0P5 vdd vss vbp vbn x a1 a2 a3 b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_a_b1b2b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 x1 b midn_a_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 midn_a_b1b2b3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_a_b1b2b3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_b2_b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 midp_b1_b2 a2 midp_b2_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 x1 b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI31_0P5




.subckt SAEDRVT14_OAI31_0P75 vdd vss vbp vbn x a1 a2 a3 b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_a_b1b2b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 x1 b midn_a_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 midn_a_b1b2b3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_a_b1b2b3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_b2_b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 midp_b1_b2 a2 midp_b2_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 x1 b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI31_0P75




.subckt SAEDRVT14_OAI311_0P5 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 midn_b_c1c2c3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_a_b b2 midn_b_c1c2c3 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x1 b1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 midn_b_c1c2c3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_b_c1c2c3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 x1 a1 midp_c1_c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 x1 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_c1_c2 a2 midp_c2_c3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_c2_c3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 x1 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI311_0P5




.subckt SAEDRVT14_OAI311_0P75 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 midn_b_c1c2c3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_a_b b2 midn_b_c1c2c3 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x1 b1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 midn_b_c1c2c3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_b_c1c2c3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 x1 a1 midp_c1_c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 x1 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_c1_c2 a2 midp_c2_c3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_c2_c3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 x1 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI311_0P75




.subckt SAEDRVT14_OAI311_1 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 midn_b_c1c2c3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_a_b b2 midn_b_c1c2c3 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x1 b1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 midn_b_c1c2c3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_b_c1c2c3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 x1 a1 midp_c1_c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 x1 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_c1_c2 a2 midp_c2_c3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_c2_c3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 x1 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI311_1




.subckt SAEDRVT14_OAI311_2 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 midn_b_c1c2c3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_a_b b2 midn_b_c1c2c3 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x1 b1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 midn_b_c1c2c3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_b_c1c2c3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 x1 a1 midp_c1_c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 x1 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_c1_c2 a2 midp_c2_c3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_c2_c3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 x1 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI311_2




.subckt SAEDRVT14_OAI311_4 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 midn_b_c1c2c3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_a_b b2 midn_b_c1c2c3 vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x1 b1 midn_a_b vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 midn_b_c1c2c3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_b_c1c2c3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 x1 a1 midp_c1_c2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 x1 b1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 midp_c1_c2 a2 midp_c2_c3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_c2_c3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp0 x1 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI311_4




.subckt SAEDRVT14_OAI31_1 vdd vss vbp vbn x a1 a2 a3 b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_a_b1b2b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 x1 b midn_a_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 midn_a_b1b2b3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_a_b1b2b3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_b2_b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 midp_b1_b2 a2 midp_b2_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 x1 b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI31_1




.subckt SAEDRVT14_OAI31_2 vdd vss vbp vbn x a1 a2 a3 b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_a_b1b2b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 x1 b midn_a_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_a_b1b2b3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_a_b1b2b3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_b2_b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 midp_b1_b2 a2 midp_b2_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OAI31_2




.subckt SAEDRVT14_OAI31_4 vdd vss vbp vbn x a1 a2 a3 b
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 midn_a_b1b2b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 x1 b midn_a_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_a_b1b2b3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_a_b1b2b3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_b2_b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 midp_b1_b2 a2 midp_b2_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x1 b vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OAI31_4




.subckt SAEDRVT14_OAI32_0P5 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 midn_a1a2_b1b2b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 x1 b1 midn_a1a2_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 x1 b2 midn_a1a2_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_a1a2_b1b2b3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_a1a2_b1b2b3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 midp_b2_b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x1 b1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 midp_a1_a2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 midp_b1_b2 a2 midp_b2_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OAI32_0P5




.subckt SAEDRVT14_OAI32_0P75 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 midn_a1a2_b1b2b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 x1 b1 midn_a1a2_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 x1 b2 midn_a1a2_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_a1a2_b1b2b3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_a1a2_b1b2b3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 midp_b2_b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x1 b1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 midp_a1_a2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 midp_b1_b2 a2 midp_b2_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OAI32_0P75




.subckt SAEDRVT14_OAI32_1 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 midn_a1a2_b1b2b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 x1 b1 midn_a1a2_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 x1 b2 midn_a1a2_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_a1a2_b1b2b3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_a1a2_b1b2b3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 midp_b2_b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x1 b1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 midp_a1_a2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 midp_b1_b2 a2 midp_b2_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OAI32_1




.subckt SAEDRVT14_OAI32_2 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 midn_a1a2_b1b2b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 x1 b1 midn_a1a2_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 x1 b2 midn_a1a2_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_a1a2_b1b2b3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_a1a2_b1b2b3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 midp_b2_b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x1 b1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 midp_a1_a2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 midp_b1_b2 a2 midp_b2_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OAI32_2




.subckt SAEDRVT14_OAI32_4 vdd vss vbp vbn x a1 a2 a3 b1 b2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 midn_a1a2_b1b2b3 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 x1 b1 midn_a1a2_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 x1 b2 midn_a1a2_b1b2b3 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 midn_a1a2_b1b2b3 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 midn_a1a2_b1b2b3 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 midp_b2_b3 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 x1 b1 midp_a1_a2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 midp_a1_a2 b2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 midp_b1_b2 a2 midp_b2_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 x1 a1 midp_b1_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OAI32_4




.subckt SAEDRVT14_OAI33_0P5 vdd vss vbp vbn x a1 a2 a3 b1 b2 b3
xn5 x1 a3 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn4 midn_a1a2a3_b1b2b3 b3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn3 x1 a1 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 x1 a2 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn1 midn_a1a2a3_b1b2b3 b1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 midn_a1a2a3_b1b2b3 b2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xp6 midp_a2_a3 a3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp5 midp_b2_b3 b3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp4 x1 a1 midp_a1_a2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp3 midp_a1_a2 a2 midp_a2_a3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 midp_b1_b2 b2 midp_b2_b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 x1 b1 midp_b1_b2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI33_0P5




.subckt SAEDRVT14_OAI33_0P75 vdd vss vbp vbn x a1 a2 a3 b1 b2 b3
xn5 x1 a3 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn4 midn_a1a2a3_b1b2b3 b3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn3 x1 a1 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 x1 a2 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn1 midn_a1a2a3_b1b2b3 b1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 midn_a1a2a3_b1b2b3 b2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xp6 midp_a2_a3 a3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp5 midp_b2_b3 b3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp4 x1 a1 midp_a1_a2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp3 midp_a1_a2 a2 midp_a2_a3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp2 midp_b1_b2 b2 midp_b2_b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 x1 b1 midp_b1_b2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI33_0P75




.subckt SAEDRVT14_OAI33_1 vdd vss vbp vbn x a1 a2 a3 b1 b2 b3
xn5 x1 a3 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn4 midn_a1a2a3_b1b2b3 b3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn3 x1 a1 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 x1 a2 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn1 midn_a1a2a3_b1b2b3 b1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 midn_a1a2a3_b1b2b3 b2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xp6 midp_a2_a3 a3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp5 midp_b2_b3 b3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp4 x1 a1 midp_a1_a2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp3 midp_a1_a2 a2 midp_a2_a3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 midp_b1_b2 b2 midp_b2_b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 x1 b1 midp_b1_b2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI33_1




.subckt SAEDRVT14_OAI33_2 vdd vss vbp vbn x a1 a2 a3 b1 b2 b3
xn5 x1 a3 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn4 midn_a1a2a3_b1b2b3 b3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn3 x1 a1 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 x1 a2 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn1 midn_a1a2a3_b1b2b3 b1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 midn_a1a2a3_b1b2b3 b2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xp6 midp_a2_a3 a3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp5 midp_b2_b3 b3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp4 x1 a1 midp_a1_a2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp3 midp_a1_a2 a2 midp_a2_a3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 midp_b1_b2 b2 midp_b2_b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 x1 b1 midp_b1_b2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI33_2




.subckt SAEDRVT14_OAI33_4 vdd vss vbp vbn x a1 a2 a3 b1 b2 b3
xn5 x1 a3 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn4 midn_a1a2a3_b1b2b3 b3 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn3 x1 a1 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 x1 a2 midn_a1a2a3_b1b2b3 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn1 midn_a1a2a3_b1b2b3 b1 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 midn_a1a2a3_b1b2b3 b2 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xmnbuf2 x d1g2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmnbuf1 d1g2 x1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xp6 midp_a2_a3 a3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp5 midp_b2_b3 b3 vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp4 x1 a1 midp_a1_a2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp3 midp_a1_a2 a2 midp_a2_a3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp2 midp_b1_b2 b2 midp_b2_b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 x1 b1 midp_b1_b2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmpbuf2 x d1g2 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmpbuf1 d1g2 x1 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_OAI33_4




.subckt SAEDRVT14_OR2_0P5 vdd vss vbp vbn x a1 a2
xmi0#2fn3 i0#2fint_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fint_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 i0#2fint_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2_0P5




.subckt SAEDRVT14_OR2_0P75 vdd vss vbp vbn x a1 a2
xmi0#2fn2 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn1 i0#2fint_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fint_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp2 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp1 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp0 i0#2fint_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2_0P75




.subckt SAEDRVT14_OR2_1 vdd vss vbp vbn x a1 a2
xmi0#2fn2 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn1 i0#2fint_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 i0#2fint_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp2 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp0 i0#2fint_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2_1




.subckt SAEDRVT14_OR2_2 vdd vss vbp vbn x a1 a2
xmi0#2fn2 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn1 i0#2fint_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 i0#2fint_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp1 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0 i0#2fint_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OR2_2




.subckt SAEDRVT14_OR2_4 vdd vss vbp vbn x a1 a2
xmi0#2fn2 x i0#2fint_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fn1 i0#2fint_zn a1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi0#2fn0 i0#2fint_zn a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp1_1 i0#2fmidp_a_b_1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0_1 i0#2fint_zn a1 i0#2fmidp_a_b_1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 x i0#2fint_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fp1 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp0 i0#2fint_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OR2_4




.subckt SAEDRVT14_OR2B_PMM_2 vdd vss vddr vbp vbn x a b
xn3 int_zn isonb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=3
xn0 int_zn b vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xmn3 isonb a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xp3 midp_a_b isonb vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x int_zn vddr vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp1 int_zn b midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp3 isonb a vddr vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2B_PMM_2




.subckt SAEDRVT14_OR2B_PMM_8 vdd vss vddr vbp vbn x a b
xn3 int_zn isonb vss vbn n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn0 int_zn b vss vbn n08_rev2 l=0.014u nf=4 m=1 nfin=3
xmn3 isonb a vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xp33 midp_a_b3 isonb vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp32 midp_a_b2 isonb vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp31 midp_a_b1 isonb vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp13 int_zn b midp_a_b3 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp12 int_zn b midp_a_b2 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp11 int_zn b midp_a_b1 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 midp_a_b isonb vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x int_zn vddr vbp p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp1 int_zn b midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp3 isonb a vddr vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OR2B_PMM_8




.subckt SAEDRVT14_OR2B_PSECO_1 vdd vss vddr x a b
xn3 int_zn isonb vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 x int_zn vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 int_zn b vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=3
xmn5 vss int_zn vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 isonb a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp3 midp_a_b isonb vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x int_zn vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 int_zn b midp_a_b vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp5 vddr int_zn vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 isonb a vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2B_PSECO_1




.subckt SAEDRVT14_OR2B_PSECO_2 vdd vss vddr x a b
xn3 int_zn isonb vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 x int_zn vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn0 int_zn b vss vss n08_rev2 l=0.014u nf=1 m=1 nfin=3
xmn3 isonb a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp3 midp_a_b isonb vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x int_zn vddr vddr p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp1 int_zn b midp_a_b vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp3 isonb a vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2B_PSECO_2




.subckt SAEDRVT14_OR2B_PSECO_4 vdd vss vddr x a b
xn3 int_zn isonb vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn2 x int_zn vss vss n08_rev2 l=0.014u nf=4 m=1 nfin=4
xn0 int_zn b vss vss n08_rev2 l=0.014u nf=2 m=1 nfin=3
xmn3 isonb a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp31 midp_a_b1 isonb vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp11 int_zn b midp_a_b1 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 midp_a_b isonb vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x int_zn vddr vddr p08_rev2 l=0.014u nf=4 m=1 nfin=4
xp1 int_zn b midp_a_b vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp3 isonb a vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2B_PSECO_4




.subckt SAEDRVT14_OR2B_PSECO_8 vdd vss vddr x a b
xn3 int_zn isonb vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=4
xn2 x int_zn vss vss n08_rev2 l=0.014u nf=8 m=1 nfin=4
xn0 int_zn b vss vss n08_rev2 l=0.014u nf=3 m=1 nfin=3
xmn3 isonb a vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xp32 midp_a_b2 isonb vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp31 midp_a_b1 isonb vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp12 int_zn b midp_a_b2 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp11 int_zn b midp_a_b1 vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp3 midp_a_b isonb vddr vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp2 x int_zn vddr vddr p08_rev2 l=0.014u nf=8 m=1 nfin=4
xp1 int_zn b midp_a_b vddr p08_rev2 l=0.014u nf=1 m=1 nfin=4
xmp3 isonb a vddr vddr p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2B_PSECO_8




.subckt SAEDRVT14_OR2_ECO_2 vdd vss vbp vbn x a1 a2
xmn3 int_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 x int_zn vss vbn n08_rev l=0.014u nf=2 m=2 nfin=4
xmn0 int_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 midp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=2 nfin=4
xmp1 int_zn a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OR2_ECO_2




.subckt SAEDRVT14_OR2_ISO_1 ck en vbn vbp vdd vss x
xp3 midp_a_b en vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp2 x int_zn vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 int_zn ck midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 int_zn en vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 int_zn ck vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2_ISO_1




.subckt SAEDRVT14_OR2_ISO_4 ck en vbn vbp vdd vss x
xp3 midp_a_b en vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp2 x int_zn vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 int_zn ck midp_a_b vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xn3 int_zn en vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn2 x int_zn vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 int_zn ck vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2_ISO_4




.subckt SAEDRVT14_OR2_MM_0P5 vdd vss vbp vbn x a1 a2
xmi0#2fn3 int_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn0 int_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp1 int_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2_MM_0P5




.subckt SAEDRVT14_OR2_MM_0P75 vdd vss vbp vbn x a1 a2
xmi0#2fn3 int_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn0 int_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp1 int_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2_MM_0P75




.subckt SAEDRVT14_OR2_MM_12 vdd vss vbp vbn x a1 a2
xmi0#2fn3 int_zn a2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmi0#2fn2 x int_zn vss vbn n08_rev l=0.014u nf=12 m=1 nfin=4
xmi0#2fn0 int_zn a1 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmi0#2fp33 i0#2fmidp_a_b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp32 i0#2fmidp_a_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp31 i0#2fmidp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp13 int_zn a1 i0#2fmidp_a_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp12 int_zn a1 i0#2fmidp_a_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp11 int_zn a1 i0#2fmidp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 x int_zn vdd vbp p08_rev l=0.014u nf=12 m=1 nfin=4
xmi0#2fp1 int_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OR2_MM_12




.subckt SAEDRVT14_OR2_MM_16 vdd vss vbp vbn x a1 a2
xmi0#2fn3 int_zn a2 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmi0#2fn2 x int_zn vss vbn n08_rev l=0.014u nf=16 m=1 nfin=4
xmi0#2fn0 int_zn a1 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=3
xmi0#2fp33 i0#2fmidp_a_b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp32 i0#2fmidp_a_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp31 i0#2fmidp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp13 int_zn a1 i0#2fmidp_a_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp12 int_zn a1 i0#2fmidp_a_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp11 int_zn a1 i0#2fmidp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 x int_zn vdd vbp p08_rev l=0.014u nf=16 m=1 nfin=4
xmi0#2fp1 int_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OR2_MM_16




.subckt SAEDRVT14_OR2_MM_1P5 vdd vss vbp vbn x a1 a2
xmi0#2fn3 int_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi0#2fn0 int_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
xmi0#2fp1 int_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2_MM_1P5




.subckt SAEDRVT14_OR2_MM_1 vdd vss vbp vbn x a1 a2
xmi0#2fn3 int_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fn0 int_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp2 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp1 int_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2_MM_1




.subckt SAEDRVT14_OR2_MM_20 vdd vss vbp vbn x a1 a2
xmi0#2fn3 int_zn a2 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=3
xmi0#2fn2 x int_zn vss vbn n08_rev l=0.014u nf=20 m=1 nfin=4
xmi0#2fn0 int_zn a1 vss vbn n08_rev l=0.014u nf=5 m=1 nfin=3
xmi0#2fp34 i0#2fmidp_a_b4 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp33 i0#2fmidp_a_b3 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp32 i0#2fmidp_a_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp31 i0#2fmidp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp14 int_zn a1 i0#2fmidp_a_b4 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp13 int_zn a1 i0#2fmidp_a_b3 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp12 int_zn a1 i0#2fmidp_a_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp11 int_zn a1 i0#2fmidp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 x int_zn vdd vbp p08_rev l=0.014u nf=20 m=1 nfin=4
xmi0#2fp1 int_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OR2_MM_20




.subckt SAEDRVT14_OR2_MM_2 vdd vss vbp vbn x a1 a2
xmi0#2fn3 int_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fn2 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fn0 int_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp2 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmi0#2fp1 int_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2_MM_2




.subckt SAEDRVT14_OR2_MM_3 vdd vss vbp vbn x a1 a2
xmi0#2fn3 int_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fn2 x int_zn vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmi0#2fn0 int_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 x int_zn vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmi0#2fp1 int_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OR2_MM_3




.subckt SAEDRVT14_OR2_MM_4 vdd vss vbp vbn x a1 a2
xmi0#2fn3 int_zn a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fn2 x int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fn0 int_zn a1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmi0#2fp31 i0#2fmidp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp11 int_zn a1 i0#2fmidp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmi0#2fp2 x int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmi0#2fp1 int_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR2_MM_4




.subckt SAEDRVT14_OR2_MM_6 vdd vss vbp vbn x a1 a2
xmi0#2fn3 int_zn a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi0#2fn2 x int_zn vss vbn n08_rev l=0.014u nf=6 m=1 nfin=4
xmi0#2fn0 int_zn a1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmi0#2fp31 i0#2fmidp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp11 int_zn a1 i0#2fmidp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 x int_zn vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=4
xmi0#2fp1 int_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OR2_MM_6




.subckt SAEDRVT14_OR2_MM_8 vdd vss vbp vbn x a1 a2
xmi0#2fn3 int_zn a2 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmi0#2fn2 x int_zn vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmi0#2fn0 int_zn a1 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmi0#2fp32 i0#2fmidp_a_b2 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp31 i0#2fmidp_a_b1 a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp12 int_zn a1 i0#2fmidp_a_b2 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp11 int_zn a1 i0#2fmidp_a_b1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp3 i0#2fmidp_a_b a2 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmi0#2fp2 x int_zn vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
xmi0#2fp1 int_zn a1 i0#2fmidp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OR2_MM_8




.subckt SAEDRVT14_OR3_0P5 vdd vss vbp vbn x a1 a2 a3
xmn3 int_zn a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn1 int_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 int_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_b_c a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp2 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 int_zn a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR3_0P5




.subckt SAEDRVT14_OR3_0P75 vdd vss vbp vbn x a1 a2 a3
xmn3 int_zn a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn2 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 int_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 int_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_b_c a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 int_zn a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OR3_0P75




.subckt SAEDRVT14_OR3_1 vdd vss vbp vbn x a1 a2 a3
xmn3 int_zn a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x int_zn vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 int_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 int_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_b_c a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x int_zn vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 int_zn a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_OR3_1




.subckt SAEDRVT14_OR3_2 vdd vss vbp vbn x a1 a2 a3
xmn3 int_zn a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x int_zn vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 int_zn a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 int_zn a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp3 midp_b_c a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x int_zn vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 int_zn a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OR3_2




.subckt SAEDRVT14_OR3_4 vdd vss vbp vbn x a1 a2 a3
xmn3 int_zn a3 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmn2 x int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn1 int_zn a1 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmn0 int_zn a2 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=2
xmp3_1 midp_b_c_1 a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1_1 midp_a_b a2 midp_b_c_1 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 midp_b_c a3 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 int_zn a1 midp_a_b vbp p08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_OR3_4




.subckt SAEDRVT14_OR4_1 vdd vss vbp vbn x a1 a2 a3 a4
xmn4 net17 a4 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 net17 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x net17 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 net17 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 net17 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 midp_c_d a4 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 midp_b_c a3 midp_c_d vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp2 x net17 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 net17 a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OR4_1




.subckt SAEDRVT14_OR4_2 vdd vss vbp vbn x a1 a2 a3 a4
xmn4 net17 a4 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn3 net17 a3 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn2 x net17 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 net17 a1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn0 net17 a2 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmp4 midp_c_d a4 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 midp_b_c a3 midp_c_d vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 x net17 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=4
xmp1 midp_a_b a2 midp_b_c vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 net17 a1 midp_a_b vbp p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_OR4_2




.subckt SAEDRVT14_PGATDRV_V1_8 vddp vdd vss vbp vbn vddc enxb
xn1 vss enxb vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xp1 vddc enxb vddp vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_PGATDRV_V1_8




.subckt SAEDRVT14_SRLD_3 vdd vss vbp vbn q qn s r
xmp9 qn qf vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp8 sx s vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp7 q qf_x vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp6 net21 rx vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp5 qf_x s net21 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp4 rx r vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 net025 qf_x vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 net021 qf vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp1 qf sx vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp1 qf r net025 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 qf_x s net021 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmn8 qn qf vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn7 q qf_x vss vbn n08_rev l=0.014u nf=3 m=1 nfin=4
xmn6 sx s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn5 qf_x s vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn4 rx r vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 qf qf_x vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn2 qf_x qf vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 qf sx net22 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 net22 r vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_SRLD_3




.subckt SAEDRVT14_SRRDPQ_1 ck d nrestore q qn save vdd vddr vss
xm13 net8 net1556 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn15 jk jk2 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm0 net28 nrestore _n766 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn21 netn102 saven vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn20 jk2 jk netn102 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn19 netn10 restore vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn18 _n766 jk netn10 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn22 saven save vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn32 netn103 save vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn33 jk2 net8 netn103 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn26 restore nrestore vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm5 net2 ckn vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm7 net1556 net8 net2 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn03 hjf d vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm11 net29 net28 net7 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn13 q net8 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm3 net28 net29 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm12 net7 ckp vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm15 qn net1556 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn011 ckn ck vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn1 net29 ckn hjf vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn012 ckp ckn vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn7 net1556 ckp _n766 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp11 net28 restore _n766 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp15 jk jk2 vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp19 _n766 jk netp10 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp18 netp10 nrestore vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp1 net29 ckp hjf vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp7 net1556 ckn _n766 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp21 jk2 jk netp102 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp26 restore nrestore vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp22 saven save vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp33 jk2 net8 netp103 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm17 qn net1556 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm4 net3 ckp vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm6 net1556 net8 net3 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm1 netp102 save vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm8 netp103 saven vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp03 hjf d vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm18 q net8 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm9 net29 net28 net9 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp011 ckn ck vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm10 net9 ckn vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp012 ckp ckn vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm14 net8 net1556 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm2 net28 net29 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
.ends SAEDRVT14_SRRDPQ_1




.subckt SAEDRVT14_SRRDPQ_2 ck d nrestore q qn save vdd vddr vss
xm13 net8 net1556 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn15 jk jk2 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm0 net28 nrestore _n766 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn21 netn102 saven vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn20 jk2 jk netn102 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn19 netn10 restore vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn18 _n766 jk netn10 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn22 saven save vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xmn32 netn103 save vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn33 jk2 net8 netn103 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn26 restore nrestore vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm5 net2 ckn vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm7 net1556 net8 net2 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn03 hjf d vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm11 net29 net28 net7 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn13 q net8 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm3 net28 net29 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm12 net7 ckp vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm15 qn net1556 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn011 ckn ck vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xmn1 net29 ckn hjf vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn012 ckp ckn vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xmn7 net1556 ckp _n766 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp11 net28 restore _n766 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp15 jk jk2 vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp19 _n766 jk netp10 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp18 netp10 nrestore vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp1 net29 ckp hjf vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp7 net1556 ckn _n766 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp21 jk2 jk netp102 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp26 restore nrestore vdd vdd p08_rev l=0.014u nf=2 m=1 nfin=4
xmp22 saven save vddr vdd p08_rev l=0.014u nf=2 m=1 nfin=4
xmp33 jk2 net8 netp103 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm17 qn net1556 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm4 net3 ckp vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm6 net1556 net8 net3 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm1 netp102 save vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm8 netp103 saven vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp03 hjf d vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm18 q net8 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm9 net29 net28 net9 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp011 ckn ck vdd vdd p08_rev l=0.014u nf=2 m=1 nfin=4
xm10 net9 ckn vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp012 ckp ckn vdd vdd p08_rev l=0.014u nf=2 m=1 nfin=4
xm14 net8 net1556 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm2 net28 net29 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
.ends SAEDRVT14_SRRDPQ_2




.subckt SAEDRVT14_SRRDPQ4_1 ck d1 d2 d3 d4 nrestore q1 q2 q3 q4 qn1 qn2 qn3 qn4 save vdd vddr vss
xm177 net282 nrestore _n7662 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn7 net15561 ckp _n7661 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn1 net291 ckn hjf1 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm180 jk2 jk212 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm182 net82 net15562 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm15 qn1 net15561 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm12 net71 ckp vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm183 net15563 ckp _n7663 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm184 net293 ckn hjf3 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm3 net281 net291 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn13 q1 net81 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm142 net291 net281 net71 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn03 hjf1 d1 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm187 qn3 net15563 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm188 net731 ckp vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm190 net283 net293 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm191 q3 net83 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm192 net293 net283 net731 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm253 net284 nrestore _n7664 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm7 net15561 net81 net69 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm195 hjf3 d3 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm5 net69 ckn vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn33 jk211 net81 netn1031 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm201 net15563 net83 net23 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn32 netn1031 save vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn18 _n7661 jk1 netn101 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm202 net23 ckn vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn19 netn101 restore vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn20 jk211 jk1 netn1021 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn21 netn1021 saven vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm205 jk213 net83 netn1033 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm206 netn1033 save vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm207 _n7663 jk3 netn103 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm0 net281 nrestore _n7661 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm208 netn103 restore vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm209 jk213 jk3 netn1023 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm210 netn1023 saven vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm256 jk4 jk214 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn15 jk1 jk211 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm13 net81 net15561 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm145 net15562 ckp _n7662 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm215 net283 nrestore _n7663 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm218 jk3 jk213 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm220 net83 net15563 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm146 net292 ckn hjf2 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm149 qn2 net15562 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm150 net72 ckp vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm152 net282 net292 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm153 q2 net82 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm154 net292 net282 net72 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm221 net15564 ckp _n7664 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm222 net294 ckn hjf4 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm225 qn4 net15564 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm157 hjf2 d2 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm226 net85 ckp vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm228 net284 net294 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm229 q4 net84 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm230 net294 net284 net85 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm163 net15562 net82 net79 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm164 net79 ckn vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm233 hjf4 d4 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm167 jk212 net82 netn1032 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm168 netn1032 save vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm169 _n7662 jk2 netn102 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm170 netn102 restore vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm171 jk212 jk2 netn1022 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm239 net15564 net84 net24 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm172 netn1022 saven vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm240 net24 ckn vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm243 jk214 net84 netn1034 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm244 netn1034 save vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm245 _n7664 jk4 netn104 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm246 netn104 restore vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm248 netn1024 saven vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm247 jk214 jk4 netn1024 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm9 ckp ckn vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm258 net84 net15564 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm26 saven save vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm25 restore nrestore vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm11 ckn ck vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm178 _n7662 jk2 netp102 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm179 jk2 jk212 vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm2 net281 net291 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm14 net81 net15561 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm181 net282 restore _n7662 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm141 net91 ckn vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm143 net291 net281 net91 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm185 net283 net293 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm18 q1 net81 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm186 net83 net15563 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp03 hjf1 d1 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm189 net93 ckn vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm144 netp1031 saven vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm1 netp1021 save vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm254 _n7664 jk4 netp104 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm255 jk4 jk214 vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm193 net293 net283 net93 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm6 net15561 net81 net70 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm194 q3 net83 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm4 net70 ckp vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm17 qn1 net15561 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp33 jk211 net81 netp1031 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm196 hjf3 d3 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm197 netp1033 saven vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm198 netp1023 save vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm199 net15563 net83 net33 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm200 net33 ckp vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm203 qn3 net15563 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp21 jk211 jk1 netp1021 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp7 net15561 ckn _n7661 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm204 jk213 net83 netp1033 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp1 net291 ckp hjf1 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp18 netp101 nrestore vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp19 _n7661 jk1 netp101 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp15 jk1 jk211 vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm211 jk213 jk3 netp1023 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm252 netp104 nrestore vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm251 net294 ckp hjf4 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm212 net15563 ckn _n7663 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm213 net293 ckp hjf3 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp11 net281 restore _n7661 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm214 netp103 nrestore vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm216 _n7663 jk3 netp103 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm217 jk3 jk213 vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm219 net283 restore _n7663 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm147 net282 net292 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm148 net82 net15562 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm151 net92 ckn vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm223 net284 net294 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm155 net292 net282 net92 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm224 net84 net15564 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm156 q2 net82 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm227 net94 ckn vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm250 net15564 ckn _n7664 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm249 jk214 jk4 netp1024 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm257 net284 restore _n7664 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm158 hjf2 d2 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm159 netp1032 saven vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm160 netp1022 save vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm161 net15562 net82 net745 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm162 net745 ckp vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm231 net294 net284 net94 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm232 q4 net84 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm234 hjf4 d4 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm235 netp1034 saven vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm236 netp1024 save vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm165 qn2 net15562 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm166 jk212 net82 netp1032 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm237 net15564 net84 net34 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm238 net34 ckp vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm173 jk212 jk2 netp1022 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm241 qn4 net15564 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm242 jk214 net84 netp1034 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm174 net15562 ckn _n7662 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm175 net292 ckp hjf2 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm176 netp102 nrestore vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm8 ckp ckn vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm24 restore nrestore vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm27 saven save vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm10 ckn ck vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_SRRDPQ4_1




.subckt SAEDRVT14_SRRDPQ4_2 ck d1 d2 d3 d4 nrestore q1 q2 q3 q4 qn1 qn2 qn3 qn4 save vdd vddr vss
xm418 net282 nrestore _n7662 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn7 net15561 ckp _n7661 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn1 net291 ckn hjf1 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm415 jk2 jk212 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm413 net82 net15562 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm15 qn1 net15561 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn33 jk211 net81 netn1031 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm349 net294 net284 net183 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm352 q4 net84 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm5 net184 ckn vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm397 hjf3 d3 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm7 net15561 net81 net184 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm354 net284 net294 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm359 net183 ckp vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm360 hjf2 d2 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm401 net284 nrestore _n7664 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm403 net293 net283 net731 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm404 q3 net83 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm146 net292 ckn hjf2 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm369 net83 net15563 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm371 jk3 jk213 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm374 net283 nrestore _n7663 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm145 net15562 ckp _n7662 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm312 net84 net15564 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm13 net81 net15561 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm315 jk214 jk4 netn1024 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm316 netn1024 saven vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm317 netn104 restore vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm318 _n7664 jk4 netn104 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn15 jk1 jk211 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm378 jk4 jk214 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm321 netn1034 save vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm322 jk214 net84 netn1034 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm382 netn1023 saven vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm411 net293 ckn hjf3 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm383 jk213 jk3 netn1023 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm326 net24 ckn vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm328 netn1022 saven vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm329 net15564 net84 net24 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm384 netn103 restore vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm0 net281 nrestore _n7661 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm385 _n7663 jk3 netn103 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm386 netn1033 save vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm387 jk213 net83 netn1033 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm330 jk212 jk2 netn1022 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm331 netn102 restore vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm332 _n7662 jk2 netn102 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm333 netn1032 save vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm334 jk212 net82 netn1032 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn21 netn1021 saven vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn20 jk211 jk1 netn1021 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn19 netn101 restore vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm390 net23 ckn vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn18 _n7661 jk1 netn101 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn32 netn1031 save vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm362 qn4 net15564 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm405 net283 net293 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm342 hjf4 d4 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm366 net294 ckn hjf4 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm407 net731 ckp vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm408 qn3 net15563 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn03 hjf1 d1 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm367 net15564 ckp _n7664 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm368 net292 net282 net72 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm153 q2 net82 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm152 net282 net292 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm150 net72 ckp vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm391 net15563 net83 net23 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm345 net186 ckn vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm149 qn2 net15562 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm142 net291 net281 net71 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xmn13 q1 net81 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm3 net281 net291 vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm346 net15562 net82 net186 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm9 ckp ckn vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm412 net15563 ckp _n7663 vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm12 net71 ckp vss vss n08_rev l=0.014u nf=1.0 m=1 nfin=4
xm26 saven save vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm25 restore nrestore vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm11 ckn ck vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm417 _n7662 jk2 netp102 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm416 jk2 jk212 vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm2 net281 net291 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm14 net81 net15561 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm414 net282 restore _n7662 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm396 hjf3 d3 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm348 net15562 net82 net745 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm350 netp1022 save vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp33 jk211 net81 netp1031 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm351 netp1032 saven vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm353 hjf2 d2 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm17 qn1 net15561 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm4 net185 ckp vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm398 q3 net83 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm355 net284 restore _n7664 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm6 net15561 net81 net185 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm399 net293 net283 net93 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm356 jk214 jk4 netp1024 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm357 net15564 ckn _n7664 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm358 net94 ckn vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm400 jk4 jk214 vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm402 _n7664 jk4 netp104 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm361 q2 net82 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm1 netp1021 save vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm144 netp1031 saven vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm147 net282 net292 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm141 net91 ckn vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm370 net283 restore _n7663 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm372 jk3 jk213 vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm373 _n7663 jk3 netp103 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm375 netp103 nrestore vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp11 net281 restore _n7661 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm376 net293 ckp hjf3 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm319 netp102 nrestore vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm377 net15563 ckn _n7663 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm320 net292 ckp hjf2 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm379 net294 ckp hjf4 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm380 netp104 nrestore vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm381 jk213 jk3 netp1023 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp15 jk1 jk211 vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm323 net15562 ckn _n7662 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp19 _n7661 jk1 netp101 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm324 jk214 net84 netp1034 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm325 qn4 net15564 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm327 jk212 jk2 netp1022 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp18 netp101 nrestore vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp1 net291 ckp hjf1 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm388 jk213 net83 netp1033 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm335 net34 ckp vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm336 net15564 net84 net34 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp7 net15561 ckn _n7661 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm337 jk212 net82 netp1032 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm338 qn2 net15562 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp21 jk211 jk1 netp1021 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm339 netp1024 save vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm389 qn3 net15563 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm340 netp1034 saven vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm341 hjf4 d4 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm363 net84 net15564 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm364 net292 net282 net92 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm406 net93 ckn vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm365 net284 net294 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm343 q4 net84 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xmp03 hjf1 d1 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm409 net83 net15563 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm18 q1 net81 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm410 net283 net293 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm143 net291 net281 net91 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm151 net92 ckn vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm344 net294 net284 net94 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm392 net33 ckp vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm393 net15563 net83 net33 vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm148 net82 net15562 vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm8 ckp ckn vdd vdd p08_rev l=0.014u nf=2 m=1 nfin=4
xm394 netp1023 save vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm24 restore nrestore vdd vdd p08_rev l=0.014u nf=2 m=1 nfin=4
xm27 saven save vddr vdd p08_rev l=0.014u nf=2 m=1 nfin=4
xm10 ckn ck vdd vdd p08_rev l=0.014u nf=2 m=1 nfin=4
xm347 net745 ckp vdd vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
xm395 netp1033 saven vddr vdd p08_rev l=0.014u nf=1.0 m=1 nfin=4
.ends SAEDRVT14_SRRDPQ4_2




.subckt SAEDRVT14_SSRRDPQ_1
xm27 qn ckp net3 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm25 qn q vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm23 q net3 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm21 net33 ckn net3 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm19 net4 ckn net28 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm17 net4 net33 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm15 net33 net28 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm13 d ckp net28 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm9 ckp ckn vdd vdd p08_rev l=0.014u nf=2 m=1 nfin=4
xm1 ckn sr vdd vdd p08_rev l=0.014u nf=2 m=1 nfin=4
xm0 ckn ck vdd vdd p08_rev l=0.014u nf=2 m=1 nfin=4
xm28 qn ckn net3 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm26 qn q vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm24 q net3 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm22 net33 ckp net3 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm20 net4 ckp net28 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm18 net4 net33 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm16 net33 net28 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm14 d ckn net28 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm10 ckp ckn vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm3 net22 ck vss vss n08_rev l=0.014u nf=2 m=1 nfin=4
xm2 ckn sr net22 vss n08_rev l=0.014u nf=2 m=1 nfin=4
.ends SAEDRVT14_SSRRDPQ_1




.subckt SAEDRVT14_SSRRDPQ_2
xm27 qn ckp net3 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm25 qn q vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm23 q net3 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm21 net33 ckn net3 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm19 net4 ckn net28 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm17 net4 net33 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm15 net33 net28 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm13 d ckp net28 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm9 ckp ckn vdd vdd p08_rev l=0.014u nf=4 m=1 nfin=4
xm1 ckn sr vdd vdd p08_rev l=0.014u nf=4 m=1 nfin=4
xm0 ckn ck vdd vdd p08_rev l=0.014u nf=4 m=1 nfin=4
xm28 qn ckn net3 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm26 qn q vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm24 q net3 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm22 net33 ckp net3 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm20 net4 ckp net28 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm18 net4 net33 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm16 net33 net28 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm14 d ckn net28 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm10 ckp ckn vss vss n08_rev l=0.014u nf=4 m=1 nfin=4
xm3 net22 ck vss vss n08_rev l=0.014u nf=4 m=1 nfin=4
xm2 ckn sr net22 vss n08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_SSRRDPQ_2




.subckt SAEDRVT14_SSRRDPQ4_1 d1 d2 d3 d4 q1 q2 q3 q4 qn1 qn2 qn3 qn4 sr vdd vddr vss ck
xm21 net139 ckn net150 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm13 d1 ckp net140 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm15 net139 net140 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm23 q1 net150 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm19 net138 ckn net140 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm17 net138 net139 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm25 qn1 q1 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm27 qn1 ckp net150 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm89 d3 ckp net146 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm98 q3 net151 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm90 net145 net146 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm91 net144 ckn net146 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm100 qn3 q3 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm93 net144 net145 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm96 net145 ckn net151 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm102 qn3 ckp net151 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm80 net142 ckn net152 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm73 d2 ckp net143 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm74 net142 net143 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm82 q2 net152 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm75 net141 ckn net143 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm77 net141 net142 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm84 qn2 q2 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm86 qn2 ckp net152 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm105 d4 ckp net149 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm114 q4 net153 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm106 net148 net149 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm107 net147 ckn net149 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm116 qn4 q4 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm9 ckp ckn vdd vdd p08_rev l=0.014u nf=4 m=1 nfin=4
xm109 net147 net148 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm112 net148 ckn net153 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm1 ckn sr vdd vdd p08_rev l=0.014u nf=4 m=1 nfin=4
xm0 ckn ck vdd vdd p08_rev l=0.014u nf=4 m=1 nfin=4
xm118 qn4 ckp net153 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm14 d1 ckn net140 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm22 net139 ckp net150 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm24 q1 net150 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm18 net138 net139 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm16 net139 net140 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm26 qn1 q1 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm28 qn1 ckn net150 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm20 net138 ckp net140 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm97 net145 ckp net151 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm88 d3 ckn net146 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm99 q3 net151 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm92 net144 net145 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm94 net145 net146 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm101 qn3 q3 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm103 qn3 ckn net151 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm72 d2 ckn net143 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm81 net142 ckp net152 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm83 q2 net152 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm76 net141 net142 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm78 net142 net143 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm85 qn2 q2 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm87 qn2 ckn net152 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm79 net141 ckp net143 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm104 d4 ckn net149 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm113 net148 ckp net153 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm115 q4 net153 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm108 net147 net148 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm95 net144 ckp net146 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm10 ckp ckn vss vss n08_rev l=0.014u nf=4 m=1 nfin=4
xm3 net22 ck vss vss n08_rev l=0.014u nf=4 m=1 nfin=4
xm2 ckn sr net22 vss n08_rev l=0.014u nf=4 m=1 nfin=4
xm110 net148 net149 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm117 qn4 q4 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm119 qn4 ckn net153 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm111 net147 ckp net149 vss n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_SSRRDPQ4_1




.subckt SAEDRVT14_SSRRDPQ4_2 d1 d2 d3 d4 q1 q2 q3 q4 qn1 qn2 qn3 qn4 sr vdd vddr vss ck
xm62 net146 ckn net148 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm70 qn4 ckp net149 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm60 net146 net147 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm68 qn4 q4 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm58 net147 net148 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm66 q4 net149 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm64 net147 ckn net149 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm56 d4 ckp net148 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm54 qn3 ckp net145 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm46 net142 ckn net144 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm52 qn3 q3 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm44 net142 net143 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm42 net143 net144 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm50 q3 net145 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm48 net143 ckn net145 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm30 net138 ckn net140 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm38 qn2 ckp net141 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm28 net138 net139 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm36 qn2 q2 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm26 net139 net140 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm34 q2 net141 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm32 net139 ckn net141 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm24 d2 ckp net140 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm19 net134 ckn net136 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm27 qn1 ckp net137 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm25 qn1 q1 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm17 net134 net135 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm23 q1 net137 vddr vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm9 ckp ckn vdd vdd p08_rev l=0.014u nf=8 m=1 nfin=4
xm40 d3 ckp net144 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm1 ckn sr vdd vdd p08_rev l=0.014u nf=8 m=1 nfin=4
xm0 ckn ck vdd vdd p08_rev l=0.014u nf=8 m=1 nfin=4
xm21 net135 ckn net137 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm15 net135 net136 vdd vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm13 d1 ckp net136 vdd p08_rev l=0.014u nf=1 m=1 nfin=4
xm63 net146 ckp net148 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm71 qn4 ckn net149 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm61 net146 net147 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm69 qn4 q4 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm59 net147 net148 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm67 q4 net149 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm57 d4 ckn net148 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm65 net147 ckp net149 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm45 net142 net143 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm47 net142 ckp net144 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm53 qn3 q3 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm51 q3 net145 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm43 net143 net144 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm55 qn3 ckn net145 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm41 d3 ckn net144 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm49 net143 ckp net145 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm31 net138 ckp net140 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm39 qn2 ckn net141 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm29 net138 net139 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm37 qn2 q2 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm27_1 net139 net140 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm35 q2 net141 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm25_1 d2 ckn net140 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm33 net139 ckp net141 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm20 net134 ckp net136 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm26_1 qn1 q1 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm18 net134 net135 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm24_1 q1 net137 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm22 net135 ckp net137 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm10 ckp ckn vss vss n08_rev l=0.014u nf=8 m=1 nfin=4
xm16 net135 net136 vss vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm3 net22 ck vss vss n08_rev l=0.014u nf=8 m=1 nfin=4
xm2 ckn sr net22 vss n08_rev l=0.014u nf=8 m=1 nfin=4
xm14 d1 ckn net136 vss n08_rev l=0.014u nf=1 m=1 nfin=4
xm28_1 qn1 ckn net137 vss n08_rev l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_SSRRDPQ4_1




.subckt SAEDRVT14_SYNC2CDCMSFQ_1 vdd vss vbp vbn q qsrc ckdst cksrc dsrc sdidst sdisrc sendst sensrc
xsrcdff#2fn1 srcdff#2fckbb srcdff#2fckb vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fn0 srcdff#2fckb cksrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn13 srcdff#2fibase#2fnet046 srcdff#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn12 srcdff#2fmq srcdff#2fckbb srcdff#2fibase#2fnet048 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn11 srcdff#2fibase#2fnet048 srcdff#2fmq_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn10 srcdff#2fmq_x srcdff#2fmq vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn9 srcdff#2fqf_x srcdff#2fckb srcdff#2fibase#2fnet046 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn8 srcdff#2fqf srcdff#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn6 srcdff#2fmq srcdff#2fckb srcdff#2fibase#2fnet028 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn5 srcdff#2fmq_x srcdff#2fckbb srcdff#2fqf_x vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn0 srcdff#2fibase#2fnet028 srcdff#2fnet050 vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi3#2fn0 ddst srcdff#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi2#2fn0 srcdff_qb srcdff#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi0#2fn17 srcdff#2fi0#2fseb sensrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn3 srcdff#2fnet050 srcdff#2fi0#2fseb srcdff#2fi0#2fnet22 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn2 srcdff#2fi0#2fnet22 dsrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn1 srcdff#2fnet050 sensrc srcdff#2fi0#2fnet19 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn0 srcdff#2fi0#2fnet19 sdisrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xn20 qsrc srcdff_qb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xi9#2fn20 q i9#2fd4lat vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fn19 i9#2fckbb i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fn18 i9#2fckb ckdst vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi9#2fi31#2fn17 i9#2fi31#2fseb sendst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn3 i9#2fdb i9#2fi31#2fseb i9#2fi31#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn2 i9#2fi31#2fnet22 ddst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn1 i9#2fdb sendst i9#2fi31#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn0 i9#2fi31#2fnet19 sdidst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi3#2fn12 i9#2fi3#2fmq_x i9#2fd4lat i9#2fi3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fn11 i9#2fi3#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fn10 i9#2fd4lat i9#2fi3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fn7 i9#2fi3#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fn6 i9#2fi3#2fmq_x i9#2fd3lat i9#2fi3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn12 i9#2fi2#2fmq_x i9#2fd3lat i9#2fi2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fn11 i9#2fi2#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn10 i9#2fd3lat i9#2fi2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fn7 i9#2fi2#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn6 i9#2fi2#2fmq_x i9#2fd2lat i9#2fi2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn12 i9#2fi1#2fmq_x i9#2fd2lat i9#2fi1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fn11 i9#2fi1#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn10 i9#2fd2lat i9#2fi1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fn7 i9#2fi1#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn6 i9#2fi1#2fmq_x i9#2fd1lat i9#2fi1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn12 i9#2fi0#2fmq_x i9#2fd1lat i9#2fi0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fn11 i9#2fi0#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn10 i9#2fd1lat i9#2fi0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fn7 i9#2fi0#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn6 i9#2fi0#2fmq_x i9#2fdb i9#2fi0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xsrcdff#2fp1 srcdff#2fckbb srcdff#2fckb vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fp0 srcdff#2fckb cksrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp11 srcdff#2fibase#2fnet045 srcdff#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp10 srcdff#2fmq srcdff#2fckb srcdff#2fibase#2fnet047 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp9 srcdff#2fibase#2fnet047 srcdff#2fmq_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp8 srcdff#2fmq_x srcdff#2fmq vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp7 srcdff#2fqf_x srcdff#2fckbb srcdff#2fibase#2fnet045 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp6 srcdff#2fqf srcdff#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp4 srcdff#2fmq srcdff#2fckbb srcdff#2fibase#2fnet027 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp3 srcdff#2fqf_x srcdff#2fckb srcdff#2fmq_x vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp1 srcdff#2fibase#2fnet027 srcdff#2fnet050 vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi3#2fp1 ddst srcdff#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi2#2fp1 srcdff_qb srcdff#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi0#2fp15 srcdff#2fi0#2fseb sensrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp3 srcdff#2fnet050 sensrc srcdff#2fi0#2fnet21 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp2 srcdff#2fi0#2fnet21 dsrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp1 srcdff#2fnet050 srcdff#2fi0#2fseb srcdff#2fi0#2fnet20 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp0 srcdff#2fi0#2fnet20 sdisrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xp18 qsrc srcdff_qb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xi9#2fp18 q i9#2fd4lat vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fp17 i9#2fckbb i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fp16 i9#2fckb ckdst vdd vbp p08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi9#2fi31#2fp15 i9#2fi31#2fseb sendst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp3 i9#2fdb sendst i9#2fi31#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp2 i9#2fi31#2fnet21 ddst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp1 i9#2fdb i9#2fi31#2fseb i9#2fi31#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp0 i9#2fi31#2fnet20 sdidst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi3#2fp10 i9#2fi3#2fmq_x i9#2fd4lat i9#2fi3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp9 i9#2fi3#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp8 i9#2fd4lat i9#2fi3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fp5 i9#2fi3#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp4 i9#2fi3#2fmq_x i9#2fd3lat i9#2fi3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp10 i9#2fi2#2fmq_x i9#2fd3lat i9#2fi2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp9 i9#2fi2#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp8 i9#2fd3lat i9#2fi2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fp5 i9#2fi2#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp4 i9#2fi2#2fmq_x i9#2fd2lat i9#2fi2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp10 i9#2fi1#2fmq_x i9#2fd2lat i9#2fi1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp9 i9#2fi1#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp8 i9#2fd2lat i9#2fi1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fp5 i9#2fi1#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp4 i9#2fi1#2fmq_x i9#2fd1lat i9#2fi1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp10 i9#2fi0#2fmq_x i9#2fd1lat i9#2fi0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp9 i9#2fi0#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp8 i9#2fd1lat i9#2fi0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fp5 i9#2fi0#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp4 i9#2fi0#2fmq_x i9#2fdb i9#2fi0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC2CDCMSFQ_1




.subckt SAEDRVT14_SYNC2FLSH2MSFQ_1 vdd vss vbp vbn q sdo ck d flsh park_hi sc1 sdi
xn12 cka ckab vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn10 midn_a_b1b2 ck vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn9 ckab ck vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn4 q d4lat vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 ckab flsh vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn20 sdo d4lat vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 ckb bhix midn_a_b1b2 vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn2 bhix flsh vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmn1 bhix sc1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 midn_a_b1b2 park_hi vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
ximux#2fn17 imux#2fseb park_hi vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmn3 db imux#2fseb imux#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmn2 imux#2fnet22 d vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmn1 db park_hi imux#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmn0 imux#2fnet19 sdi vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn11 i3#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn11 i2#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn11 i1#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn11 i0#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn6 i0#2fmq_x db i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xp10 cka ckab vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp7 ckab ck net61 vbp p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 q d4lat vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 net61 flsh vdd vbp p08_rev2 l=0.014u nf=3 m=1 nfin=4
xmp23 sdo d4lat vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 midp_b1_b2 ck vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp4 net041 flsh vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
xmp3 ckb bhix vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 ckb park_hi midp_b1_b2 vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 bhix sc1 net041 vbp p08_rev l=0.014u nf=1 m=1 nfin=3
ximux#2fp15 imux#2fseb park_hi vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmp3 db park_hi imux#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmp2 imux#2fnet21 d vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmp1 db imux#2fseb imux#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmp0 imux#2fnet20 sdi vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp4 i0#2fmq_x db i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC2FLSH2MSFQ_1




.subckt SAEDRVT14_SYNC2FLSHMSFQNS_1 vdd vss vbp vbn q ck d flsh
xn0 flshb flsh vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xi43#2fn2 ckbb ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi43#2fn1 i43#2fmidn_a_b flshb vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi43#2fn0 ckb ck i43#2fmidn_a_b vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi42#2fmn2 cka ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmn1 ckab flsh vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmn0 ckab ck vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=2   
xi3#2fn12 i3#2fmq_x i3#2fnet013 i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn11 i3#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 i3#2fnet013 i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn7 i3#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fmn4 q i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn11 i2#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn11 i1#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn11 i0#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn6 i0#2fmq_x d i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xp0 flshb flsh vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xi43#2fp2 ckbb ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi43#2fp1 ckb ck vdd vbp p08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi43#2fp0 ckb flshb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp12 i42#2fmidp_a_b2 flsh vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp11 i42#2fmidp_a_b1 flsh vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp02 ckab ck i42#2fmidp_a_b2 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp01 ckab ck i42#2fmidp_a_b1 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp2 cka ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp1 i42#2fmidp_a_b flsh vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp0 ckab ck i42#2fmidp_a_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp10 i3#2fmq_x i3#2fnet013 i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 i3#2fnet013 i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp5 i3#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fmp4 q i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp4 i0#2fmq_x d i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC2FLSHMSFQNS_1




.subckt SAEDRVT14_SYNC2FLSHMSFQNS_6 vdd vss vbp vbn q ck d flsh
xn4 q qb vss vbn n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn3 qb d4lat vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn0 flshb flsh vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xi43#2fn2 ckbb ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi43#2fn1 i43#2fmidn_a_b flshb vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi43#2fn0 ckb ck i43#2fmidn_a_b vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi42#2fmn2 cka ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmn1 ckab flsh vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmn0 ckab ck vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=2   
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn11 i3#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn11 i2#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn11 i1#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn11 i0#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn6 i0#2fmq_x d i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xp4 qb d4lat vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp2 q qb vdd vbp p08_rev2 l=0.014u nf=6 m=1 nfin=4
xp0 flshb flsh vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xi43#2fp2 ckbb ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi43#2fp1 ckb ck vdd vbp p08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi43#2fp0 ckb flshb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp12 i42#2fmidp_a_b2 flsh vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp11 i42#2fmidp_a_b1 flsh vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp02 ckab ck i42#2fmidp_a_b2 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp01 ckab ck i42#2fmidp_a_b1 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp2 cka ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp1 i42#2fmidp_a_b flsh vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp0 ckab ck i42#2fmidp_a_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp4 i0#2fmq_x d i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC2FLSHMSFQNS_6




.subckt SAEDRVT14_SYNC2MSFQ_1 vdd vss vbp vbn q ck d sdi sen
xn20 q d4lat vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn19 ckbb ckb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn18 ckb ck vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xi31#2fn17 i31#2fseb sen vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmn3 db i31#2fseb i31#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmn2 i31#2fnet22 d vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmn1 db sen i31#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmn0 i31#2fnet19 sdi vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn11 i3#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn11 i2#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn11 i1#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn11 i0#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn6 i0#2fmq_x db i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xp18 q d4lat vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp17 ckbb ckb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp16 ckb ck vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xi31#2fp15 i31#2fseb sen vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmp3 db sen i31#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmp2 i31#2fnet21 d vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmp1 db i31#2fseb i31#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmp0 i31#2fnet20 sdi vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp4 i0#2fmq_x db i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC2MSFQ_1




.subckt SAEDRVT14_SYNC2MSFQNS_6 vdd vss vbp vbn q ck d
xn19 ckbb ckb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn18 ckb ck vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn4 q qb vss vbn n08_rev2 l=0.014u nf=6 m=1 nfin=4
xn3 qb d4lat vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn11 i3#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn11 i2#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn11 i1#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn11 i0#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn6 i0#2fmq_x d i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xp17 ckbb ckb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp16 ckb ck vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp4 qb d4lat vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp2 q qb vdd vbp p08_rev2 l=0.014u nf=6 m=1 nfin=4
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp4 i0#2fmq_x d i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC2MSFQNS_6




.subckt SAEDRVT14_SYNC2P5CDCMSFQ_1 vdd vss vbp vbn q qsrc ckdst cksrc dsrc sdidst sdisrc sendst sensrc
xsrcdff#2fn1 srcdff#2fckbb srcdff#2fckb vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fn0 srcdff#2fckb cksrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn13 srcdff#2fibase#2fnet046 srcdff#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn12 srcdff#2fmq srcdff#2fckbb srcdff#2fibase#2fnet048 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn11 srcdff#2fibase#2fnet048 srcdff#2fmq_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn10 srcdff#2fmq_x srcdff#2fmq vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn9 srcdff#2fqf_x srcdff#2fckb srcdff#2fibase#2fnet046 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn8 srcdff#2fqf srcdff#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn6 srcdff#2fmq srcdff#2fckb srcdff#2fibase#2fnet028 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn5 srcdff#2fmq_x srcdff#2fckbb srcdff#2fqf_x vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn0 srcdff#2fibase#2fnet028 srcdff#2fnet050 vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi3#2fn0 ddst srcdff#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi2#2fn0 srcdff_qb srcdff#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi0#2fn17 srcdff#2fi0#2fseb sensrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn3 srcdff#2fnet050 srcdff#2fi0#2fseb srcdff#2fi0#2fnet22 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn2 srcdff#2fi0#2fnet22 dsrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn1 srcdff#2fnet050 sensrc srcdff#2fi0#2fnet19 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn0 srcdff#2fi0#2fnet19 sdisrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xn20 qsrc srcdff_qb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xi9#2fsdi_latch#2fn24 i9#2fsdi_latch#2fdb sdidst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fn19 i9#2fsdi_latch#2fckbb i9#2fsdi_latch#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fn18 i9#2fsdi_latch#2fckb ckdst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fn14 i9#2fsdil_q i9#2fsdi_latch#2fqf_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fsdi_latch#2fi31#2fn23 i9#2fsdi_latch#2fi31#2fnet61 i9#2fsdi_latch#2fqf vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fi31#2fn20 i9#2fsdi_latch#2fdb i9#2fsdi_latch#2fckb i9#2fsdi_latch#2fqf_x vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fi31#2fn12 i9#2fsdi_latch#2fqf_x i9#2fsdi_latch#2fckbb i9#2fsdi_latch#2fi31#2fnet61 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fi31#2fn10 i9#2fsdi_latch#2fqf i9#2fsdi_latch#2fqf_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fn20 q i9#2fd5lat vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fn19 i9#2fckbb i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fn18 i9#2fckb ckdst vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi9#2fi4#2fn12 i9#2fi4#2fmq_x i9#2fd5lat i9#2fi4#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fn11 i9#2fi4#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fn10 i9#2fd5lat i9#2fi4#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fn7 i9#2fi4#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fn6 i9#2fi4#2fmq_x i9#2fd4lat i9#2fi4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi30#2fn17 i9#2fi30#2fseb sendst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi30#2fmn3 i9#2fdb i9#2fi30#2fseb i9#2fi30#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi30#2fmn2 i9#2fi30#2fnet22 ddst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi30#2fmn1 i9#2fdb sendst i9#2fi30#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi30#2fmn0 i9#2fi30#2fnet19 i9#2fsdil_q vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi3#2fn12 i9#2fi3#2fmq_x i9#2fd4lat i9#2fi3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fn11 i9#2fi3#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fn10 i9#2fd4lat i9#2fi3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fn7 i9#2fi3#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fn6 i9#2fi3#2fmq_x i9#2fd3lat i9#2fi3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn12 i9#2fi2#2fmq_x i9#2fd3lat i9#2fi2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fn11 i9#2fi2#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn10 i9#2fd3lat i9#2fi2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fn7 i9#2fi2#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn6 i9#2fi2#2fmq_x i9#2fd2lat i9#2fi2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn12 i9#2fi1#2fmq_x i9#2fd2lat i9#2fi1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fn11 i9#2fi1#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn10 i9#2fd2lat i9#2fi1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fn7 i9#2fi1#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn6 i9#2fi1#2fmq_x i9#2fd1lat i9#2fi1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn12 i9#2fi0#2fmq_x i9#2fd1lat i9#2fi0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fn11 i9#2fi0#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn10 i9#2fd1lat i9#2fi0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fn7 i9#2fi0#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn6 i9#2fi0#2fmq_x i9#2fdb i9#2fi0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xsrcdff#2fp1 srcdff#2fckbb srcdff#2fckb vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fp0 srcdff#2fckb cksrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp11 srcdff#2fibase#2fnet045 srcdff#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp10 srcdff#2fmq srcdff#2fckb srcdff#2fibase#2fnet047 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp9 srcdff#2fibase#2fnet047 srcdff#2fmq_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp8 srcdff#2fmq_x srcdff#2fmq vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp7 srcdff#2fqf_x srcdff#2fckbb srcdff#2fibase#2fnet045 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp6 srcdff#2fqf srcdff#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp4 srcdff#2fmq srcdff#2fckbb srcdff#2fibase#2fnet027 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp3 srcdff#2fqf_x srcdff#2fckb srcdff#2fmq_x vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp1 srcdff#2fibase#2fnet027 srcdff#2fnet050 vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi3#2fp1 ddst srcdff#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi2#2fp1 srcdff_qb srcdff#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi0#2fp15 srcdff#2fi0#2fseb sensrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp3 srcdff#2fnet050 sensrc srcdff#2fi0#2fnet21 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp2 srcdff#2fi0#2fnet21 dsrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp1 srcdff#2fnet050 srcdff#2fi0#2fseb srcdff#2fi0#2fnet20 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp0 srcdff#2fi0#2fnet20 sdisrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xp18 qsrc srcdff_qb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xi9#2fsdi_latch#2fp23 i9#2fsdi_latch#2fdb sdidst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fp17 i9#2fsdi_latch#2fckbb i9#2fsdi_latch#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fsdi_latch#2fp16 i9#2fsdi_latch#2fckb ckdst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fsdi_latch#2fp11 i9#2fsdil_q i9#2fsdi_latch#2fqf_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fsdi_latch#2fi31#2fp21 i9#2fsdi_latch#2fqf_x i9#2fsdi_latch#2fckb i9#2fsdi_latch#2fi31#2fnet98 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fi31#2fp18 i9#2fsdi_latch#2fqf_x i9#2fsdi_latch#2fckbb i9#2fsdi_latch#2fdb vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fi31#2fp9 i9#2fsdi_latch#2fi31#2fnet98 i9#2fsdi_latch#2fqf vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fi31#2fp8 i9#2fsdi_latch#2fqf i9#2fsdi_latch#2fqf_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fp18 q i9#2fd5lat vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fp17 i9#2fckbb i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fp16 i9#2fckb ckdst vdd vbp p08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi9#2fi4#2fp10 i9#2fi4#2fmq_x i9#2fd5lat i9#2fi4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp9 i9#2fi4#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp8 i9#2fd5lat i9#2fi4#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fp5 i9#2fi4#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp4 i9#2fi4#2fmq_x i9#2fd4lat i9#2fi4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi30#2fp15 i9#2fi30#2fseb sendst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi30#2fmp3 i9#2fdb sendst i9#2fi30#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi30#2fmp2 i9#2fi30#2fnet21 ddst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi30#2fmp1 i9#2fdb i9#2fi30#2fseb i9#2fi30#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi30#2fmp0 i9#2fi30#2fnet20 i9#2fsdil_q vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi3#2fp10 i9#2fi3#2fmq_x i9#2fd4lat i9#2fi3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp9 i9#2fi3#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp8 i9#2fd4lat i9#2fi3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fp5 i9#2fi3#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp4 i9#2fi3#2fmq_x i9#2fd3lat i9#2fi3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp10 i9#2fi2#2fmq_x i9#2fd3lat i9#2fi2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp9 i9#2fi2#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp8 i9#2fd3lat i9#2fi2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fp5 i9#2fi2#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp4 i9#2fi2#2fmq_x i9#2fd2lat i9#2fi2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp10 i9#2fi1#2fmq_x i9#2fd2lat i9#2fi1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp9 i9#2fi1#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp8 i9#2fd2lat i9#2fi1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fp5 i9#2fi1#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp4 i9#2fi1#2fmq_x i9#2fd1lat i9#2fi1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp10 i9#2fi0#2fmq_x i9#2fd1lat i9#2fi0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp9 i9#2fi0#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp8 i9#2fd1lat i9#2fi0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fp5 i9#2fi0#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp4 i9#2fi0#2fmq_x i9#2fdb i9#2fi0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC2P5CDCMSFQ_1




.subckt SAEDRVT14_SYNC2P5FLSHMSFQ_1 vdd vss vbp vbn q ck d flsh sdi sen
xsdi_latch#2fn24 sdi_latch#2fdb sdi vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn19 sdi_latch#2fckbb sdi_latch#2fckb vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn18 sdi_latch#2fckb ck vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn14 sdil_q sdi_latch#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fi31#2fn23 sdi_latch#2fi31#2fnet61 sdi_latch#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn20 sdi_latch#2fdb sdi_latch#2fckb sdi_latch#2fqf_x vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn12 sdi_latch#2fqf_x sdi_latch#2fckbb sdi_latch#2fi31#2fnet61 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn10 sdi_latch#2fqf sdi_latch#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xn16 sebb seb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn15 seb flshb net58 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn14 net58 sen vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn4 q d5lat vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 flshb flsh vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xi44#2fn4 i44#2fnet20 sebb db vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi44#2fn3 i44#2fnet18 seb db vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi44#2fn2 i44#2fnet20 sdil_q vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi44#2fn0 i44#2fnet18 d vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi43#2fn2 ckbb ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi43#2fn1 i43#2fmidn_a_b flshb vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi43#2fn0 ckb ck i43#2fmidn_a_b vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi42#2fmn2 cka ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmn1 ckab flsh vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmn0 ckab ck vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi4#2fn12 i4#2fmq_x d5lat i4#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn11 i4#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn10 d5lat i4#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn7 i4#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn6 i4#2fmq_x d4lat i4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn11 i3#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn11 i2#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn11 i1#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn11 i0#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn6 i0#2fmq_x db i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fp23 sdi_latch#2fdb sdi vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fp17 sdi_latch#2fckbb sdi_latch#2fckb vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fp16 sdi_latch#2fckb ck vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fp11 sdil_q sdi_latch#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fi31#2fp21 sdi_latch#2fqf_x sdi_latch#2fckb sdi_latch#2fi31#2fnet98 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp18 sdi_latch#2fqf_x sdi_latch#2fckbb sdi_latch#2fdb vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp9 sdi_latch#2fi31#2fnet98 sdi_latch#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp8 sdi_latch#2fqf sdi_latch#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xp14 seb sen vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp13 seb flshb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp12 sebb seb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp2 q d5lat vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp0 flshb flsh vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xi44#2fp4 i44#2fnet21 seb db vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi44#2fp3 i44#2fnet19 sebb db vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi44#2fp2 i44#2fnet21 sdil_q vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi44#2fp0 i44#2fnet19 d vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi43#2fp2 ckbb ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi43#2fp1 ckb ck vdd vbp p08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi43#2fp0 ckb flshb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp12 i42#2fmidp_a_b2 flsh vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp11 i42#2fmidp_a_b1 flsh vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp02 ckab ck i42#2fmidp_a_b2 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp01 ckab ck i42#2fmidp_a_b1 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp2 cka ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp1 i42#2fmidp_a_b flsh vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp0 ckab ck i42#2fmidp_a_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fp10 i4#2fmq_x d5lat i4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp9 i4#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp8 d5lat i4#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fp5 i4#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp4 i4#2fmq_x d4lat i4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp4 i0#2fmq_x db i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC2P5FLSHMSFQ_1




.subckt SAEDRVT14_SYNC2P5RMSFQ_1 vdd vss vbp vbn q ck d reseth sdi sen
xsdi_latch#2fn24 sdi_latch#2fdb sdi vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn19 sdi_latch#2fckbb sdi_latch#2fckb vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn18 sdi_latch#2fckb ck vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn14 sdil_q sdi_latch#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fi31#2fn23 sdi_latch#2fi31#2fnet61 sdi_latch#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn20 sdi_latch#2fdb sdi_latch#2fckb sdi_latch#2fqf_x vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn12 sdi_latch#2fqf_x sdi_latch#2fckbb sdi_latch#2fi31#2fnet61 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn10 sdi_latch#2fqf sdi_latch#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xn20 q d5lat vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn19 ckbb ckb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn18 ckb ck vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn17 seb sen vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn4 db seb net69 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn3 net69 d vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 net72 sdil_q vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 db sen net72 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xmn7 resetb reseth vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xi4#2fn12 i4#2fmq_x d5lat i4#2fnet018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn11 i4#2fnet018 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn10 d5lat i4#2fmq_x i4#2fnet014 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn7 i4#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi4#2fn6 i4#2fmq_x d4lat i4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi4#2fmn4 i4#2fnet014 resetb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn11 i3#2fnet018 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x i3#2fnet014 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fmn4 i3#2fnet014 resetb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn11 i2#2fnet018 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x i2#2fnet014 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fmn4 i2#2fnet014 resetb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn11 i1#2fnet018 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x i1#2fnet014 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fmn4 i1#2fnet014 resetb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn11 i0#2fnet018 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x i0#2fnet014 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn6 i0#2fmq_x db i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmn4 i0#2fnet014 resetb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xsdi_latch#2fp23 sdi_latch#2fdb sdi vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fp17 sdi_latch#2fckbb sdi_latch#2fckb vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fp16 sdi_latch#2fckb ck vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fp11 sdil_q sdi_latch#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fi31#2fp21 sdi_latch#2fqf_x sdi_latch#2fckb sdi_latch#2fi31#2fnet98 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp18 sdi_latch#2fqf_x sdi_latch#2fckbb sdi_latch#2fdb vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp9 sdi_latch#2fi31#2fnet98 sdi_latch#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp8 sdi_latch#2fqf sdi_latch#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xp18 q d5lat vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp17 ckbb ckb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp16 ckb ck vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp15 seb sen vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp2 db sen net70 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net70 d vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net71 sdil_q vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xn1 db seb net71 vbp p08 l=0.014u nf=1 m=1 nfin=2
xmp7 resetb reseth vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xi4#2fp10 i4#2fmq_x d5lat i4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp9 i4#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp8 d5lat i4#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fp5 i4#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi4#2fp4 i4#2fmq_x d4lat i4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi4#2fmp4 d5lat resetb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fmp4 d4lat resetb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fmp4 d3lat resetb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fmp4 d2lat resetb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp4 i0#2fmq_x db i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmp4 d1lat resetb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
.ends SAEDRVT14_SYNC2P5RMSFQ_1




.subckt SAEDRVT14_SYNC2P5SMSFQ_1 vdd vss vbp vbn q ck d seth sdi sen
xsdi_latch#2fn24 sdi_latch#2fdb sdi vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn19 sdi_latch#2fckbb sdi_latch#2fckb vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn18 sdi_latch#2fckb ck vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn14 sdil_q sdi_latch#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fi31#2fn23 sdi_latch#2fi31#2fnet61 sdi_latch#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn20 sdi_latch#2fdb sdi_latch#2fckb sdi_latch#2fqf_x vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn12 sdi_latch#2fqf_x sdi_latch#2fckbb sdi_latch#2fi31#2fnet61 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn10 sdi_latch#2fqf sdi_latch#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xn20 q d5lat vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn19 ckbb ckb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn18 ckb ck vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn17 seb sen vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn4 db seb net69 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn3 net69 d vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 net72 sdil_q vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 db sen net72 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xi4#2fn12 i4#2fmq_x d5lat i4#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn11 i4#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn10 d5lat i4#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn7 i4#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi4#2fn6 i4#2fmq_x d4lat i4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi4#2fmn4 d5lat seth vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn11 i3#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fmn4 d4lat seth vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn11 i2#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fmn4 d3lat seth vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn11 i1#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fmn4 d2lat seth vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn11 i0#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn6 i0#2fmq_x db i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmn4 d1lat seth vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xsdi_latch#2fp23 sdi_latch#2fdb sdi vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fp17 sdi_latch#2fckbb sdi_latch#2fckb vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fp16 sdi_latch#2fckb ck vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fp11 sdil_q sdi_latch#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fi31#2fp21 sdi_latch#2fqf_x sdi_latch#2fckb sdi_latch#2fi31#2fnet98 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp18 sdi_latch#2fqf_x sdi_latch#2fckbb sdi_latch#2fdb vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp9 sdi_latch#2fi31#2fnet98 sdi_latch#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp8 sdi_latch#2fqf sdi_latch#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xp18 q d5lat vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp17 ckbb ckb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp16 ckb ck vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp15 seb sen vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp2 db sen net70 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net70 d vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net71 sdil_q vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xn1 db seb net71 vbp p08 l=0.014u nf=1 m=1 nfin=2
xi4#2fp10 i4#2fmq_x d5lat i4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp9 i4#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp8 d5lat i4#2fmq_x i4#2fnet014 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fp5 i4#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi4#2fp4 i4#2fmq_x d4lat i4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi4#2fmp4 i4#2fnet014 seth vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x i3#2fnet014 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fmp4 i3#2fnet014 seth vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x i2#2fnet014 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fmp4 i2#2fnet014 seth vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x i1#2fnet014 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fmp4 i1#2fnet014 seth vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x i0#2fnet014 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp4 i0#2fmq_x db i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmp4 i0#2fnet014 seth vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
.ends SAEDRVT14_SYNC2P5SMSFQ_1




.subckt SAEDRVT14_SYNC2RMSFQ_1 vdd vss vbp vbn q ck d reseth sdi sen
xn20 q d4lat vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn19 ckbb ckb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn18 ckb ck vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn17 seb sen vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn4 db seb net69 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn3 net69 d vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 net72 sdi vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 db sen net72 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xmn7 resetb reseth vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn11 i3#2fnet018 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x i3#2fnet014 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fmn4 i3#2fnet014 resetb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn11 i2#2fnet018 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x i2#2fnet014 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fmn4 i2#2fnet014 resetb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn11 i1#2fnet018 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x i1#2fnet014 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fmn4 i1#2fnet014 resetb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet018 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn11 i0#2fnet018 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x i0#2fnet014 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn6 i0#2fmq_x db i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmn4 i0#2fnet014 resetb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xp18 q d4lat vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp17 ckbb ckb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp16 ckb ck vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp15 seb sen vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp2 db sen net70 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net70 d vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net71 sdi vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xn1 db seb net71 vbp p08 l=0.014u nf=1 m=1 nfin=2
xmp7 resetb reseth vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fmp4 d4lat resetb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fmp4 d3lat resetb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fmp4 d2lat resetb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp4 i0#2fmq_x db i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmp4 d1lat resetb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
.ends SAEDRVT14_SYNC2RMSFQ_1




.subckt SAEDRVT14_SYNC2SMSFQ_1 vdd vss vbp vbn q ck d seth sdi sen
xn20 q d4lat vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn19 ckbb ckb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn18 ckb ck vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn17 seb sen vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn4 db seb net69 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn3 net69 d vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn2 net72 sdi vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 db sen net72 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn11 i3#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fmn4 d4lat seth vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn11 i2#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fmn4 d3lat seth vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn11 i1#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fmn4 d2lat seth vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn11 i0#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fn6 i0#2fmq_x db i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmn4 d1lat seth vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xp18 q d4lat vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp17 ckbb ckb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp16 ckb ck vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp15 seb sen vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp2 db sen net70 vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp1 net70 d vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xp0 net71 sdi vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xn1 db seb net71 vbp p08 l=0.014u nf=1 m=1 nfin=2
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x i3#2fnet014 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fmp4 i3#2fnet014 seth vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x i2#2fnet014 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi2#2fmp4 i2#2fnet014 seth vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x i1#2fnet014 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi1#2fmp4 i1#2fnet014 seth vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x i0#2fnet014 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fp4 i0#2fmq_x db i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi0#2fmp4 i0#2fnet014 seth vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
.ends SAEDRVT14_SYNC2SMSFQ_1




.subckt SAEDRVT14_SYNC3CDCMSFQ_1 vdd vss vbp vbn q qsrc ckdst cksrc dsrc sdidst sdisrc sendst sensrc
xsrcdff#2fn1 srcdff#2fckbb srcdff#2fckb vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fn0 srcdff#2fckb cksrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn13 srcdff#2fibase#2fnet046 srcdff#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn12 srcdff#2fmq srcdff#2fckbb srcdff#2fibase#2fnet048 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn11 srcdff#2fibase#2fnet048 srcdff#2fmq_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn10 srcdff#2fmq_x srcdff#2fmq vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn9 srcdff#2fqf_x srcdff#2fckb srcdff#2fibase#2fnet046 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn8 srcdff#2fqf srcdff#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn6 srcdff#2fmq srcdff#2fckb srcdff#2fibase#2fnet028 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn5 srcdff#2fmq_x srcdff#2fckbb srcdff#2fqf_x vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn0 srcdff#2fibase#2fnet028 srcdff#2fnet050 vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi3#2fn0 ddst srcdff#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi2#2fn0 srcdff_qb srcdff#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi0#2fn17 srcdff#2fi0#2fseb sensrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn3 srcdff#2fnet050 srcdff#2fi0#2fseb srcdff#2fi0#2fnet22 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn2 srcdff#2fi0#2fnet22 dsrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn1 srcdff#2fnet050 sensrc srcdff#2fi0#2fnet19 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn0 srcdff#2fi0#2fnet19 sdisrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xn20 qsrc srcdff_qb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xi9#2fn20 q i9#2fd6lat vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fn19 i9#2fckbb i9#2fckb vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi9#2fn18 i9#2fckb ckdst vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi9#2fi5#2fn12 i9#2fi5#2fmq_x i9#2fd6lat i9#2fi5#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi5#2fn11 i9#2fi5#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fn10 i9#2fd6lat i9#2fi5#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi5#2fn7 i9#2fi5#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fn6 i9#2fi5#2fmq_x i9#2fd5lat i9#2fi5#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fn12 i9#2fi4#2fmq_x i9#2fd5lat i9#2fi4#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fn11 i9#2fi4#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fn10 i9#2fd5lat i9#2fi4#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fn7 i9#2fi4#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fn6 i9#2fi4#2fmq_x i9#2fd4lat i9#2fi4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi31#2fn17 i9#2fi31#2fseb sendst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn3 i9#2fdb i9#2fi31#2fseb i9#2fi31#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn2 i9#2fi31#2fnet22 ddst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn1 i9#2fdb sendst i9#2fi31#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn0 i9#2fi31#2fnet19 sdidst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi3#2fn12 i9#2fi3#2fmq_x i9#2fd4lat i9#2fi3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fn11 i9#2fi3#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fn10 i9#2fd4lat i9#2fi3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fn7 i9#2fi3#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fn6 i9#2fi3#2fmq_x i9#2fd3lat i9#2fi3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn12 i9#2fi2#2fmq_x i9#2fd3lat i9#2fi2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fn11 i9#2fi2#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn10 i9#2fd3lat i9#2fi2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fn7 i9#2fi2#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn6 i9#2fi2#2fmq_x i9#2fd2lat i9#2fi2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn12 i9#2fi1#2fmq_x i9#2fd2lat i9#2fi1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fn11 i9#2fi1#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn10 i9#2fd2lat i9#2fi1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fn7 i9#2fi1#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn6 i9#2fi1#2fmq_x i9#2fd1lat i9#2fi1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn12 i9#2fi0#2fmq_x i9#2fd1lat i9#2fi0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fn11 i9#2fi0#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn10 i9#2fd1lat i9#2fi0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fn7 i9#2fi0#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn6 i9#2fi0#2fmq_x i9#2fdb i9#2fi0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xsrcdff#2fp1 srcdff#2fckbb srcdff#2fckb vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fp0 srcdff#2fckb cksrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp11 srcdff#2fibase#2fnet045 srcdff#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp10 srcdff#2fmq srcdff#2fckb srcdff#2fibase#2fnet047 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp9 srcdff#2fibase#2fnet047 srcdff#2fmq_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp8 srcdff#2fmq_x srcdff#2fmq vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp7 srcdff#2fqf_x srcdff#2fckbb srcdff#2fibase#2fnet045 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp6 srcdff#2fqf srcdff#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp4 srcdff#2fmq srcdff#2fckbb srcdff#2fibase#2fnet027 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp3 srcdff#2fqf_x srcdff#2fckb srcdff#2fmq_x vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp1 srcdff#2fibase#2fnet027 srcdff#2fnet050 vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi3#2fp1 ddst srcdff#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi2#2fp1 srcdff_qb srcdff#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi0#2fp15 srcdff#2fi0#2fseb sensrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp3 srcdff#2fnet050 sensrc srcdff#2fi0#2fnet21 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp2 srcdff#2fi0#2fnet21 dsrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp1 srcdff#2fnet050 srcdff#2fi0#2fseb srcdff#2fi0#2fnet20 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp0 srcdff#2fi0#2fnet20 sdisrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xp18 qsrc srcdff_qb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xi9#2fp18 q i9#2fd6lat vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fp17 i9#2fckbb i9#2fckb vdd vbp p08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi9#2fp16 i9#2fckb ckdst vdd vbp p08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi9#2fi5#2fp10 i9#2fi5#2fmq_x i9#2fd6lat i9#2fi5#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp9 i9#2fi5#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp8 i9#2fd6lat i9#2fi5#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi5#2fp5 i9#2fi5#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp4 i9#2fi5#2fmq_x i9#2fd5lat i9#2fi5#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp10 i9#2fi4#2fmq_x i9#2fd5lat i9#2fi4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp9 i9#2fi4#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp8 i9#2fd5lat i9#2fi4#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fp5 i9#2fi4#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp4 i9#2fi4#2fmq_x i9#2fd4lat i9#2fi4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi31#2fp15 i9#2fi31#2fseb sendst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp3 i9#2fdb sendst i9#2fi31#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp2 i9#2fi31#2fnet21 ddst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp1 i9#2fdb i9#2fi31#2fseb i9#2fi31#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp0 i9#2fi31#2fnet20 sdidst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi3#2fp10 i9#2fi3#2fmq_x i9#2fd4lat i9#2fi3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp9 i9#2fi3#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp8 i9#2fd4lat i9#2fi3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fp5 i9#2fi3#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp4 i9#2fi3#2fmq_x i9#2fd3lat i9#2fi3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp10 i9#2fi2#2fmq_x i9#2fd3lat i9#2fi2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp9 i9#2fi2#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp8 i9#2fd3lat i9#2fi2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fp5 i9#2fi2#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp4 i9#2fi2#2fmq_x i9#2fd2lat i9#2fi2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp10 i9#2fi1#2fmq_x i9#2fd2lat i9#2fi1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp9 i9#2fi1#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp8 i9#2fd2lat i9#2fi1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fp5 i9#2fi1#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp4 i9#2fi1#2fmq_x i9#2fd1lat i9#2fi1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp10 i9#2fi0#2fmq_x i9#2fd1lat i9#2fi0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp9 i9#2fi0#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp8 i9#2fd1lat i9#2fi0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fp5 i9#2fi0#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp4 i9#2fi0#2fmq_x i9#2fdb i9#2fi0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC3CDCMSFQ_1




.subckt SAEDRVT14_SYNC3FLSH2MSFQ_1 vdd vss vbp vbn q sdo ck d flsh park_hi sc1 sdi
xn12 cka ckab vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn10 midn_a_b1b2 ck vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn9 ckab ck vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn4 q d6lat vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn2 ckab flsh vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xmn20 sdo d6lat vss vbn n08_rev l=0.014u nf=1 m=1 nfin=2
xmn4 ckbb ckb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn3 ckb bhix midn_a_b1b2 vbn n08_rev l=0.014u nf=2 m=1 nfin=4
xmn2 bhix flsh vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn1 bhix sc1 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 midn_a_b1b2 park_hi vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
ximux#2fn17 imux#2fseb park_hi vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmn3 db imux#2fseb imux#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmn2 imux#2fnet22 d vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmn1 db park_hi imux#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmn0 imux#2fnet19 sdi vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi5#2fn12 i5#2fmq_x d6lat i5#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fn11 i5#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn10 d6lat i5#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fn7 i5#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn6 i5#2fmq_x d5lat i5#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn12 i4#2fmq_x d5lat i4#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn11 i4#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn10 d5lat i4#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn7 i4#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn6 i4#2fmq_x d4lat i4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn11 i3#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn11 i2#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn11 i1#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn11 i0#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn6 i0#2fmq_x db i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xp10 cka ckab vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp7 ckab ck net61 vbp p08_rev2 l=0.014u nf=3 m=1 nfin=4
xp2 q d6lat vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp1 net61 flsh vdd vbp p08_rev2 l=0.014u nf=3 m=1 nfin=4
xmp23 sdo d6lat vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=2
xmp5 midp_b1_b2 ck vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp4 net041 flsh vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp3 ckb bhix vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp2 ckb park_hi midp_b1_b2 vbp p08_rev l=0.014u nf=3 m=1 nfin=4
xmp1 ckbb ckb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 bhix sc1 net041 vbp p08_rev l=0.014u nf=1 m=1 nfin=4
ximux#2fp15 imux#2fseb park_hi vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmp3 db park_hi imux#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmp2 imux#2fnet21 d vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmp1 db imux#2fseb imux#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
ximux#2fmp0 imux#2fnet20 sdi vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi5#2fp10 i5#2fmq_x d6lat i5#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp9 i5#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp8 d6lat i5#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fp5 i5#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp4 i5#2fmq_x d5lat i5#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp10 i4#2fmq_x d5lat i4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp9 i4#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp8 d5lat i4#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fp5 i4#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp4 i4#2fmq_x d4lat i4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp4 i0#2fmq_x db i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC3FLSH2MSFQ_1




.subckt SAEDRVT14_SYNC3MSFQ_1 vdd vss vbp vbn q ck d sdi sen
xn20 q d6lat vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn19 ckbb ckb vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn18 ckb ck vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xi5#2fn12 i5#2fmq_x d6lat i5#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fn11 i5#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn10 d6lat i5#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fn7 i5#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn6 i5#2fmq_x d5lat i5#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn12 i4#2fmq_x d5lat i4#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn11 i4#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn10 d5lat i4#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn7 i4#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn6 i4#2fmq_x d4lat i4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi31#2fn17 i31#2fseb sen vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmn3 db i31#2fseb i31#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmn2 i31#2fnet22 d vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmn1 db sen i31#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmn0 i31#2fnet19 sdi vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn11 i3#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn11 i2#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn11 i1#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn11 i0#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn6 i0#2fmq_x db i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xp18 q d6lat vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp17 ckbb ckb vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp16 ckb ck vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xi5#2fp10 i5#2fmq_x d6lat i5#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp9 i5#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp8 d6lat i5#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fp5 i5#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp4 i5#2fmq_x d5lat i5#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp10 i4#2fmq_x d5lat i4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp9 i4#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp8 d5lat i4#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fp5 i4#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp4 i4#2fmq_x d4lat i4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi31#2fp15 i31#2fseb sen vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmp3 db sen i31#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmp2 i31#2fnet21 d vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmp1 db i31#2fseb i31#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmp0 i31#2fnet20 sdi vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp4 i0#2fmq_x db i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC3MSFQ_1




.subckt SAEDRVT14_SYNC3ORMSFQNS_1 vdd vss vbp vbn q ck d en setb te
xn19 ckb ckbb vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=3
xn3 db d vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xmn8 net031 setb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn7 q d6lat net031 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xi5#2fn12 i5#2fmq_x d6lat i5#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fn11 i5#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn10 d6lat i5#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fn7 i5#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn6 i5#2fmq_x d5lat i5#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn12 i4#2fmq_x d5lat i4#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn11 i4#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn10 d5lat i4#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn7 i4#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn6 i4#2fmq_x d4lat i4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn11 i3#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn11 i2#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn11 i1#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn11 i0#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn6 i0#2fmq_x db i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xck_gater#2fn24 ck_gater#2fe_nr_te te vss vbn n08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fn10 ck_gater#2fe_nr_te en vss vbn n08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fn1 ck_gater#2fckbb ck_gater#2fckb vss vbn n08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fn0 ck_gater#2fckb ck vss vbn n08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi31#2fn2 ckbb ck_gater#2fzn vss vbn n08 l=0.014u nf=2 m=1 nfin=4
xck_gater#2fi31#2fn1 ck_gater#2fi31#2fmidn_en_ck ck_gater#2fqf vss vbn n08 l=0.014u nf=1 m=1 nfin=3
xck_gater#2fi31#2fn0 ck_gater#2fzn ck ck_gater#2fi31#2fmidn_en_ck vbn n08 l=0.014u nf=1 m=1 nfin=3
xck_gater#2fi1#2fn23 ck_gater#2fi1#2fnet61 ck_gater#2fqf vss vbn n08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi1#2fn20 ck_gater#2fe_nr_te ck_gater#2fckb ck_gater#2fqf_x vbn n08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi1#2fn12 ck_gater#2fqf_x ck_gater#2fckbb ck_gater#2fi1#2fnet61 vbn n08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi1#2fn10 ck_gater#2fqf ck_gater#2fqf_x vss vbn n08 l=0.014u nf=1 m=1 nfin=2
xp17 ckb ckbb vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=3
xp1 db d vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xmp8 q setb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp7 q d6lat vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xi5#2fp10 i5#2fmq_x d6lat i5#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp9 i5#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp8 d6lat i5#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fp5 i5#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp4 i5#2fmq_x d5lat i5#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp10 i4#2fmq_x d5lat i4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp9 i4#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp8 d5lat i4#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fp5 i4#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp4 i4#2fmq_x d4lat i4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp4 i0#2fmq_x db i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xck_gater#2fp23 ck_gater#2fe_nr_te te ck_gater#2fnet42 vbp p08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fp22 ck_gater#2fnet42 en vdd vbp p08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fp1 ck_gater#2fckbb ck_gater#2fckb vdd vbp p08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fp0 ck_gater#2fckb ck vdd vbp p08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi31#2fp2 ckbb ck_gater#2fzn vdd vbp p08 l=0.014u nf=2 m=1 nfin=4
xck_gater#2fi31#2fp1 ck_gater#2fzn ck vdd vbp p08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi31#2fp0 ck_gater#2fzn ck_gater#2fqf vdd vbp p08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi1#2fp21 ck_gater#2fqf_x ck_gater#2fckb ck_gater#2fi1#2fnet98 vbp p08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi1#2fp18 ck_gater#2fqf_x ck_gater#2fckbb ck_gater#2fe_nr_te vbp p08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi1#2fp9 ck_gater#2fi1#2fnet98 ck_gater#2fqf vdd vbp p08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi1#2fp8 ck_gater#2fqf ck_gater#2fqf_x vdd vbp p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_SYNC3ORMSFQNS_1




.subckt SAEDRVT14_SYNC3P5CDCMSFQ_1 vdd vss vbp vbn q qsrc ckdst cksrc dsrc sdidst sdisrc sendst sensrc
xsrcdff#2fn1 srcdff#2fckbb srcdff#2fckb vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fn0 srcdff#2fckb cksrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn13 srcdff#2fibase#2fnet046 srcdff#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn12 srcdff#2fmq srcdff#2fckbb srcdff#2fibase#2fnet048 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn11 srcdff#2fibase#2fnet048 srcdff#2fmq_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn10 srcdff#2fmq_x srcdff#2fmq vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn9 srcdff#2fqf_x srcdff#2fckb srcdff#2fibase#2fnet046 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn8 srcdff#2fqf srcdff#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn6 srcdff#2fmq srcdff#2fckb srcdff#2fibase#2fnet028 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn5 srcdff#2fmq_x srcdff#2fckbb srcdff#2fqf_x vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn0 srcdff#2fibase#2fnet028 srcdff#2fnet050 vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi3#2fn0 ddst srcdff#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi2#2fn0 srcdff_qb srcdff#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi0#2fn17 srcdff#2fi0#2fseb sensrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn3 srcdff#2fnet050 srcdff#2fi0#2fseb srcdff#2fi0#2fnet22 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn2 srcdff#2fi0#2fnet22 dsrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn1 srcdff#2fnet050 sensrc srcdff#2fi0#2fnet19 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn0 srcdff#2fi0#2fnet19 sdisrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xn20 qsrc srcdff_qb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xi9#2fsdi_latch#2fn24 i9#2fsdi_latch#2fdb sdidst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fn19 i9#2fsdi_latch#2fckbb i9#2fsdi_latch#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fn18 i9#2fsdi_latch#2fckb ckdst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fn14 i9#2fsdil_q i9#2fsdi_latch#2fqf_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fsdi_latch#2fi31#2fn23 i9#2fsdi_latch#2fi31#2fnet61 i9#2fsdi_latch#2fqf vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fi31#2fn20 i9#2fsdi_latch#2fdb i9#2fsdi_latch#2fckb i9#2fsdi_latch#2fqf_x vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fi31#2fn12 i9#2fsdi_latch#2fqf_x i9#2fsdi_latch#2fckbb i9#2fsdi_latch#2fi31#2fnet61 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fi31#2fn10 i9#2fsdi_latch#2fqf i9#2fsdi_latch#2fqf_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fn20 q i9#2fd7lat vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fn19 i9#2fckbb i9#2fckb vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi9#2fn18 i9#2fckb ckdst vss vbn n08_rev3 l=0.014u nf=3 m=1 nfin=4   
xi9#2fi6#2fn12 i9#2fi6#2fmq_x i9#2fd7lat i9#2fi6#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi6#2fn11 i9#2fi6#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fn10 i9#2fd7lat i9#2fi6#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi6#2fn7 i9#2fi6#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fn6 i9#2fi6#2fmq_x i9#2fd6lat i9#2fi6#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fn12 i9#2fi5#2fmq_x i9#2fd6lat i9#2fi5#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi5#2fn11 i9#2fi5#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fn10 i9#2fd6lat i9#2fi5#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi5#2fn7 i9#2fi5#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fn6 i9#2fi5#2fmq_x i9#2fd5lat i9#2fi5#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fn12 i9#2fi4#2fmq_x i9#2fd5lat i9#2fi4#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fn11 i9#2fi4#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fn10 i9#2fd5lat i9#2fi4#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fn7 i9#2fi4#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fn6 i9#2fi4#2fmq_x i9#2fd4lat i9#2fi4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi32#2fn17 i9#2fi32#2fseb sendst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi32#2fmn3 i9#2fdb i9#2fi32#2fseb i9#2fi32#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi32#2fmn2 i9#2fi32#2fnet22 ddst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi32#2fmn1 i9#2fdb sendst i9#2fi32#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi32#2fmn0 i9#2fi32#2fnet19 i9#2fsdil_q vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi3#2fn12 i9#2fi3#2fmq_x i9#2fd4lat i9#2fi3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fn11 i9#2fi3#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fn10 i9#2fd4lat i9#2fi3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fn7 i9#2fi3#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fn6 i9#2fi3#2fmq_x i9#2fd3lat i9#2fi3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn12 i9#2fi2#2fmq_x i9#2fd3lat i9#2fi2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fn11 i9#2fi2#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn10 i9#2fd3lat i9#2fi2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fn7 i9#2fi2#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn6 i9#2fi2#2fmq_x i9#2fd2lat i9#2fi2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn12 i9#2fi1#2fmq_x i9#2fd2lat i9#2fi1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fn11 i9#2fi1#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn10 i9#2fd2lat i9#2fi1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fn7 i9#2fi1#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn6 i9#2fi1#2fmq_x i9#2fd1lat i9#2fi1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn12 i9#2fi0#2fmq_x i9#2fd1lat i9#2fi0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fn11 i9#2fi0#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn10 i9#2fd1lat i9#2fi0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fn7 i9#2fi0#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn6 i9#2fi0#2fmq_x i9#2fdb i9#2fi0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xsrcdff#2fp1 srcdff#2fckbb srcdff#2fckb vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fp0 srcdff#2fckb cksrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp11 srcdff#2fibase#2fnet045 srcdff#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp10 srcdff#2fmq srcdff#2fckb srcdff#2fibase#2fnet047 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp9 srcdff#2fibase#2fnet047 srcdff#2fmq_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp8 srcdff#2fmq_x srcdff#2fmq vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp7 srcdff#2fqf_x srcdff#2fckbb srcdff#2fibase#2fnet045 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp6 srcdff#2fqf srcdff#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp4 srcdff#2fmq srcdff#2fckbb srcdff#2fibase#2fnet027 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp3 srcdff#2fqf_x srcdff#2fckb srcdff#2fmq_x vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp1 srcdff#2fibase#2fnet027 srcdff#2fnet050 vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi3#2fp1 ddst srcdff#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi2#2fp1 srcdff_qb srcdff#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi0#2fp15 srcdff#2fi0#2fseb sensrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp3 srcdff#2fnet050 sensrc srcdff#2fi0#2fnet21 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp2 srcdff#2fi0#2fnet21 dsrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp1 srcdff#2fnet050 srcdff#2fi0#2fseb srcdff#2fi0#2fnet20 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp0 srcdff#2fi0#2fnet20 sdisrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xp18 qsrc srcdff_qb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xi9#2fsdi_latch#2fp23 i9#2fsdi_latch#2fdb sdidst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fp17 i9#2fsdi_latch#2fckbb i9#2fsdi_latch#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fsdi_latch#2fp16 i9#2fsdi_latch#2fckb ckdst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fsdi_latch#2fp11 i9#2fsdil_q i9#2fsdi_latch#2fqf_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fsdi_latch#2fi31#2fp21 i9#2fsdi_latch#2fqf_x i9#2fsdi_latch#2fckb i9#2fsdi_latch#2fi31#2fnet98 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fi31#2fp18 i9#2fsdi_latch#2fqf_x i9#2fsdi_latch#2fckbb i9#2fsdi_latch#2fdb vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fi31#2fp9 i9#2fsdi_latch#2fi31#2fnet98 i9#2fsdi_latch#2fqf vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fsdi_latch#2fi31#2fp8 i9#2fsdi_latch#2fqf i9#2fsdi_latch#2fqf_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fp18 q i9#2fd7lat vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fp17 i9#2fckbb i9#2fckb vdd vbp p08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi9#2fp16 i9#2fckb ckdst vdd vbp p08_rev3 l=0.014u nf=3 m=1 nfin=4   
xi9#2fi6#2fp10 i9#2fi6#2fmq_x i9#2fd7lat i9#2fi6#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fp9 i9#2fi6#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fp8 i9#2fd7lat i9#2fi6#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi6#2fp5 i9#2fi6#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fp4 i9#2fi6#2fmq_x i9#2fd6lat i9#2fi6#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp10 i9#2fi5#2fmq_x i9#2fd6lat i9#2fi5#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp9 i9#2fi5#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp8 i9#2fd6lat i9#2fi5#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi5#2fp5 i9#2fi5#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp4 i9#2fi5#2fmq_x i9#2fd5lat i9#2fi5#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp10 i9#2fi4#2fmq_x i9#2fd5lat i9#2fi4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp9 i9#2fi4#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp8 i9#2fd5lat i9#2fi4#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fp5 i9#2fi4#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp4 i9#2fi4#2fmq_x i9#2fd4lat i9#2fi4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi32#2fp15 i9#2fi32#2fseb sendst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi32#2fmp3 i9#2fdb sendst i9#2fi32#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi32#2fmp2 i9#2fi32#2fnet21 ddst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi32#2fmp1 i9#2fdb i9#2fi32#2fseb i9#2fi32#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi32#2fmp0 i9#2fi32#2fnet20 i9#2fsdil_q vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi3#2fp10 i9#2fi3#2fmq_x i9#2fd4lat i9#2fi3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp9 i9#2fi3#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp8 i9#2fd4lat i9#2fi3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fp5 i9#2fi3#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp4 i9#2fi3#2fmq_x i9#2fd3lat i9#2fi3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp10 i9#2fi2#2fmq_x i9#2fd3lat i9#2fi2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp9 i9#2fi2#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp8 i9#2fd3lat i9#2fi2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fp5 i9#2fi2#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp4 i9#2fi2#2fmq_x i9#2fd2lat i9#2fi2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp10 i9#2fi1#2fmq_x i9#2fd2lat i9#2fi1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp9 i9#2fi1#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp8 i9#2fd2lat i9#2fi1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fp5 i9#2fi1#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp4 i9#2fi1#2fmq_x i9#2fd1lat i9#2fi1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp10 i9#2fi0#2fmq_x i9#2fd1lat i9#2fi0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp9 i9#2fi0#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp8 i9#2fd1lat i9#2fi0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fp5 i9#2fi0#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp4 i9#2fi0#2fmq_x i9#2fdb i9#2fi0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC3P5CDCMSFQ_1




.subckt SAEDRVT14_SYNC3P5FLSHMSFQ_1 vdd vss vbp vbn q ck d flsh sdi sen
xsdi_latch#2fn24 sdi_latch#2fdb sdi vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn19 sdi_latch#2fckbb sdi_latch#2fckb vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn18 sdi_latch#2fckb ck vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn14 sdil_q sdi_latch#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fi31#2fn23 sdi_latch#2fi31#2fnet61 sdi_latch#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn20 sdi_latch#2fdb sdi_latch#2fckb sdi_latch#2fqf_x vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn12 sdi_latch#2fqf_x sdi_latch#2fckbb sdi_latch#2fi31#2fnet61 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn10 sdi_latch#2fqf sdi_latch#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xn16 sebb seb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn15 seb flshb net58 vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn14 net58 sen vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=3
xn4 q d7lat vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 flshb flsh vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xi6#2fn12 i6#2fmq_x d7lat i6#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi6#2fn11 i6#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fn10 d7lat i6#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi6#2fn7 i6#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fn6 i6#2fmq_x d6lat i6#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn12 i5#2fmq_x d6lat i5#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fn11 i5#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn10 d6lat i5#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fn7 i5#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn6 i5#2fmq_x d5lat i5#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi44#2fn4 i44#2fnet20 sebb db vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi44#2fn3 i44#2fnet18 seb db vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi44#2fn2 i44#2fnet20 sdil_q vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi44#2fn0 i44#2fnet18 d vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi43#2fn2 ckbb ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi43#2fn1 i43#2fmidn_a_b flshb vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi43#2fn0 ckb ck i43#2fmidn_a_b vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi42#2fmn2 cka ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmn1 ckab flsh vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmn0 ckab ck vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=2   
xi4#2fn12 i4#2fmq_x d5lat i4#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn11 i4#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn10 d5lat i4#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn7 i4#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn6 i4#2fmq_x d4lat i4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn11 i3#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn11 i2#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn11 i1#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn11 i0#2fnet048 ckab vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 cka vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn6 i0#2fmq_x db i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fp23 sdi_latch#2fdb sdi vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fp17 sdi_latch#2fckbb sdi_latch#2fckb vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fp16 sdi_latch#2fckb ck vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fp11 sdil_q sdi_latch#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fi31#2fp21 sdi_latch#2fqf_x sdi_latch#2fckb sdi_latch#2fi31#2fnet98 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp18 sdi_latch#2fqf_x sdi_latch#2fckbb sdi_latch#2fdb vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp9 sdi_latch#2fi31#2fnet98 sdi_latch#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp8 sdi_latch#2fqf sdi_latch#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xp14 seb sen vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp13 seb flshb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp12 sebb seb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=3
xp2 q d7lat vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp0 flshb flsh vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xi6#2fp10 i6#2fmq_x d7lat i6#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fp9 i6#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fp8 d7lat i6#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi6#2fp5 i6#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fp4 i6#2fmq_x d6lat i6#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp10 i5#2fmq_x d6lat i5#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp9 i5#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp8 d6lat i5#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fp5 i5#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp4 i5#2fmq_x d5lat i5#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi44#2fp4 i44#2fnet21 seb db vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi44#2fp3 i44#2fnet19 sebb db vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi44#2fp2 i44#2fnet21 sdil_q vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi44#2fp0 i44#2fnet19 d vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi43#2fp2 ckbb ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi43#2fp1 ckb ck vdd vbp p08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi43#2fp0 ckb flshb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp12 i42#2fmidp_a_b2 flsh vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp11 i42#2fmidp_a_b1 flsh vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp02 ckab ck i42#2fmidp_a_b2 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp01 ckab ck i42#2fmidp_a_b1 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp2 cka ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp1 i42#2fmidp_a_b flsh vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi42#2fmp0 ckab ck i42#2fmidp_a_b vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fp10 i4#2fmq_x d5lat i4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp9 i4#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp8 d5lat i4#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fp5 i4#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp4 i4#2fmq_x d4lat i4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 cka vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckab vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp4 i0#2fmq_x db i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC3P5FLSHMSFQ_1




.subckt SAEDRVT14_SYNC3P5MSFQ_1 vdd vss vbp vbn q ck d sdi sen
xsdi_latch#2fn24 sdi_latch#2fdb sdi vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn19 sdi_latch#2fckbb sdi_latch#2fckb vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn18 sdi_latch#2fckb ck vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fn14 sdil_q sdi_latch#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fi31#2fn23 sdi_latch#2fi31#2fnet61 sdi_latch#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn20 sdi_latch#2fdb sdi_latch#2fckb sdi_latch#2fqf_x vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn12 sdi_latch#2fqf_x sdi_latch#2fckbb sdi_latch#2fi31#2fnet61 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fn10 sdi_latch#2fqf sdi_latch#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xn20 q d7lat vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn19 ckbb ckb vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn18 ckb ck vss vbn n08_rev2 l=0.014u nf=3 m=1 nfin=4
xi6#2fn12 i6#2fmq_x d7lat i6#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi6#2fn11 i6#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fn10 d7lat i6#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi6#2fn7 i6#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fn6 i6#2fmq_x d6lat i6#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn12 i5#2fmq_x d6lat i5#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fn11 i5#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn10 d6lat i5#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fn7 i5#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn6 i5#2fmq_x d5lat i5#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn12 i4#2fmq_x d5lat i4#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn11 i4#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn10 d5lat i4#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn7 i4#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn6 i4#2fmq_x d4lat i4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi32#2fn17 i32#2fseb sen vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fmn3 db i32#2fseb i32#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fmn2 i32#2fnet22 d vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fmn1 db sen i32#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fmn0 i32#2fnet19 sdil_q vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn11 i3#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn11 i2#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn11 i1#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn11 i0#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn6 i0#2fmq_x db i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fp23 sdi_latch#2fdb sdi vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fp17 sdi_latch#2fckbb sdi_latch#2fckb vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fp16 sdi_latch#2fckb ck vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fp11 sdil_q sdi_latch#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=3   
xsdi_latch#2fi31#2fp21 sdi_latch#2fqf_x sdi_latch#2fckb sdi_latch#2fi31#2fnet98 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp18 sdi_latch#2fqf_x sdi_latch#2fckbb sdi_latch#2fdb vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp9 sdi_latch#2fi31#2fnet98 sdi_latch#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsdi_latch#2fi31#2fp8 sdi_latch#2fqf sdi_latch#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xp18 q d7lat vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp17 ckbb ckb vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp16 ckb ck vdd vbp p08_rev2 l=0.014u nf=3 m=1 nfin=4
xi6#2fp10 i6#2fmq_x d7lat i6#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fp9 i6#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fp8 d7lat i6#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi6#2fp5 i6#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fp4 i6#2fmq_x d6lat i6#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp10 i5#2fmq_x d6lat i5#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp9 i5#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp8 d6lat i5#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fp5 i5#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp4 i5#2fmq_x d5lat i5#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp10 i4#2fmq_x d5lat i4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp9 i4#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp8 d5lat i4#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fp5 i4#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp4 i4#2fmq_x d4lat i4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi32#2fp15 i32#2fseb sen vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fmp3 db sen i32#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fmp2 i32#2fnet21 d vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fmp1 db i32#2fseb i32#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi32#2fmp0 i32#2fnet20 sdil_q vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp4 i0#2fmq_x db i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC3P5MSFQ_1




.subckt SAEDRVT14_SYNC4CDCMSFQ_1 vdd vss vbp vbn q qsrc ckdst cksrc dsrc sdidst sdisrc sendst sensrc
xsrcdff#2fn1 srcdff#2fckbb srcdff#2fckb vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fn0 srcdff#2fckb cksrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn13 srcdff#2fibase#2fnet046 srcdff#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn12 srcdff#2fmq srcdff#2fckbb srcdff#2fibase#2fnet048 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn11 srcdff#2fibase#2fnet048 srcdff#2fmq_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn10 srcdff#2fmq_x srcdff#2fmq vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn9 srcdff#2fqf_x srcdff#2fckb srcdff#2fibase#2fnet046 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn8 srcdff#2fqf srcdff#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn6 srcdff#2fmq srcdff#2fckb srcdff#2fibase#2fnet028 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn5 srcdff#2fmq_x srcdff#2fckbb srcdff#2fqf_x vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn0 srcdff#2fibase#2fnet028 srcdff#2fnet050 vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi3#2fn0 ddst srcdff#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi2#2fn0 srcdff_qb srcdff#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi0#2fn17 srcdff#2fi0#2fseb sensrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn3 srcdff#2fnet050 srcdff#2fi0#2fseb srcdff#2fi0#2fnet22 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn2 srcdff#2fi0#2fnet22 dsrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn1 srcdff#2fnet050 sensrc srcdff#2fi0#2fnet19 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn0 srcdff#2fi0#2fnet19 sdisrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xn20 qsrc srcdff_qb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xi9#2fn20 q i9#2fd8lat vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fn19 i9#2fckbb i9#2fckb vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi9#2fn18 i9#2fckb ckdst vss vbn n08_rev3 l=0.014u nf=3 m=1 nfin=4   
xi9#2fi7#2fn12 i9#2fi7#2fmq_x i9#2fd8lat i9#2fi7#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi7#2fn11 i9#2fi7#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi7#2fn10 i9#2fd8lat i9#2fi7#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi7#2fn7 i9#2fi7#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi7#2fn6 i9#2fi7#2fmq_x i9#2fd7lat i9#2fi7#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fn12 i9#2fi6#2fmq_x i9#2fd7lat i9#2fi6#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi6#2fn11 i9#2fi6#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fn10 i9#2fd7lat i9#2fi6#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi6#2fn7 i9#2fi6#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fn6 i9#2fi6#2fmq_x i9#2fd6lat i9#2fi6#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fn12 i9#2fi5#2fmq_x i9#2fd6lat i9#2fi5#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi5#2fn11 i9#2fi5#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fn10 i9#2fd6lat i9#2fi5#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi5#2fn7 i9#2fi5#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fn6 i9#2fi5#2fmq_x i9#2fd5lat i9#2fi5#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fn12 i9#2fi4#2fmq_x i9#2fd5lat i9#2fi4#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fn11 i9#2fi4#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fn10 i9#2fd5lat i9#2fi4#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fn7 i9#2fi4#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fn6 i9#2fi4#2fmq_x i9#2fd4lat i9#2fi4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi31#2fn17 i9#2fi31#2fseb sendst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn3 i9#2fdb i9#2fi31#2fseb i9#2fi31#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn2 i9#2fi31#2fnet22 ddst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn1 i9#2fdb sendst i9#2fi31#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn0 i9#2fi31#2fnet19 sdidst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi3#2fn12 i9#2fi3#2fmq_x i9#2fd4lat i9#2fi3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fn11 i9#2fi3#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fn10 i9#2fd4lat i9#2fi3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fn7 i9#2fi3#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fn6 i9#2fi3#2fmq_x i9#2fd3lat i9#2fi3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn12 i9#2fi2#2fmq_x i9#2fd3lat i9#2fi2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fn11 i9#2fi2#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn10 i9#2fd3lat i9#2fi2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fn7 i9#2fi2#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn6 i9#2fi2#2fmq_x i9#2fd2lat i9#2fi2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn12 i9#2fi1#2fmq_x i9#2fd2lat i9#2fi1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fn11 i9#2fi1#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn10 i9#2fd2lat i9#2fi1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fn7 i9#2fi1#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn6 i9#2fi1#2fmq_x i9#2fd1lat i9#2fi1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn12 i9#2fi0#2fmq_x i9#2fd1lat i9#2fi0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fn11 i9#2fi0#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn10 i9#2fd1lat i9#2fi0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fn7 i9#2fi0#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn6 i9#2fi0#2fmq_x i9#2fdb i9#2fi0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xsrcdff#2fp1 srcdff#2fckbb srcdff#2fckb vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fp0 srcdff#2fckb cksrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp11 srcdff#2fibase#2fnet045 srcdff#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp10 srcdff#2fmq srcdff#2fckb srcdff#2fibase#2fnet047 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp9 srcdff#2fibase#2fnet047 srcdff#2fmq_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp8 srcdff#2fmq_x srcdff#2fmq vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp7 srcdff#2fqf_x srcdff#2fckbb srcdff#2fibase#2fnet045 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp6 srcdff#2fqf srcdff#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp4 srcdff#2fmq srcdff#2fckbb srcdff#2fibase#2fnet027 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp3 srcdff#2fqf_x srcdff#2fckb srcdff#2fmq_x vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp1 srcdff#2fibase#2fnet027 srcdff#2fnet050 vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi3#2fp1 ddst srcdff#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi2#2fp1 srcdff_qb srcdff#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi0#2fp15 srcdff#2fi0#2fseb sensrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp3 srcdff#2fnet050 sensrc srcdff#2fi0#2fnet21 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp2 srcdff#2fi0#2fnet21 dsrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp1 srcdff#2fnet050 srcdff#2fi0#2fseb srcdff#2fi0#2fnet20 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp0 srcdff#2fi0#2fnet20 sdisrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xp18 qsrc srcdff_qb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xi9#2fp18 q i9#2fd8lat vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fp17 i9#2fckbb i9#2fckb vdd vbp p08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi9#2fp16 i9#2fckb ckdst vdd vbp p08_rev3 l=0.014u nf=3 m=1 nfin=4   
xi9#2fi7#2fp10 i9#2fi7#2fmq_x i9#2fd8lat i9#2fi7#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi7#2fp9 i9#2fi7#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi7#2fp8 i9#2fd8lat i9#2fi7#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi7#2fp5 i9#2fi7#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi7#2fp4 i9#2fi7#2fmq_x i9#2fd7lat i9#2fi7#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fp10 i9#2fi6#2fmq_x i9#2fd7lat i9#2fi6#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fp9 i9#2fi6#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fp8 i9#2fd7lat i9#2fi6#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi6#2fp5 i9#2fi6#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fp4 i9#2fi6#2fmq_x i9#2fd6lat i9#2fi6#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp10 i9#2fi5#2fmq_x i9#2fd6lat i9#2fi5#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp9 i9#2fi5#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp8 i9#2fd6lat i9#2fi5#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi5#2fp5 i9#2fi5#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp4 i9#2fi5#2fmq_x i9#2fd5lat i9#2fi5#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp10 i9#2fi4#2fmq_x i9#2fd5lat i9#2fi4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp9 i9#2fi4#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp8 i9#2fd5lat i9#2fi4#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fp5 i9#2fi4#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp4 i9#2fi4#2fmq_x i9#2fd4lat i9#2fi4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi31#2fp15 i9#2fi31#2fseb sendst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp3 i9#2fdb sendst i9#2fi31#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp2 i9#2fi31#2fnet21 ddst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp1 i9#2fdb i9#2fi31#2fseb i9#2fi31#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp0 i9#2fi31#2fnet20 sdidst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi3#2fp10 i9#2fi3#2fmq_x i9#2fd4lat i9#2fi3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp9 i9#2fi3#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp8 i9#2fd4lat i9#2fi3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fp5 i9#2fi3#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp4 i9#2fi3#2fmq_x i9#2fd3lat i9#2fi3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp10 i9#2fi2#2fmq_x i9#2fd3lat i9#2fi2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp9 i9#2fi2#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp8 i9#2fd3lat i9#2fi2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fp5 i9#2fi2#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp4 i9#2fi2#2fmq_x i9#2fd2lat i9#2fi2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp10 i9#2fi1#2fmq_x i9#2fd2lat i9#2fi1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp9 i9#2fi1#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp8 i9#2fd2lat i9#2fi1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fp5 i9#2fi1#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp4 i9#2fi1#2fmq_x i9#2fd1lat i9#2fi1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp10 i9#2fi0#2fmq_x i9#2fd1lat i9#2fi0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp9 i9#2fi0#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp8 i9#2fd1lat i9#2fi0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fp5 i9#2fi0#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp4 i9#2fi0#2fmq_x i9#2fdb i9#2fi0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC4CDCMSFQ_1




.subckt SAEDRVT14_SYNC4MSFQ_1 vdd vss vbp vbn q ck d sdi sen
xn20 q d8lat vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn19 ckbb ckb vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=4
xn18 ckb ck vss vbn n08_rev2 l=0.014u nf=3 m=1 nfin=4
xi7#2fn12 i7#2fmq_x d8lat i7#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi7#2fn11 i7#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi7#2fn10 d8lat i7#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi7#2fn7 i7#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi7#2fn6 i7#2fmq_x d7lat i7#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fn12 i6#2fmq_x d7lat i6#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi6#2fn11 i6#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fn10 d7lat i6#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi6#2fn7 i6#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fn6 i6#2fmq_x d6lat i6#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn12 i5#2fmq_x d6lat i5#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fn11 i5#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn10 d6lat i5#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fn7 i5#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn6 i5#2fmq_x d5lat i5#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn12 i4#2fmq_x d5lat i4#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn11 i4#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn10 d5lat i4#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn7 i4#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn6 i4#2fmq_x d4lat i4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi31#2fn17 i31#2fseb sen vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmn3 db i31#2fseb i31#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmn2 i31#2fnet22 d vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmn1 db sen i31#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmn0 i31#2fnet19 sdi vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn11 i3#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn11 i2#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn11 i1#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn11 i0#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn6 i0#2fmq_x db i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xp18 q d8lat vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp17 ckbb ckb vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=4
xp16 ckb ck vdd vbp p08_rev2 l=0.014u nf=3 m=1 nfin=4
xi7#2fp10 i7#2fmq_x d8lat i7#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi7#2fp9 i7#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi7#2fp8 d8lat i7#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi7#2fp5 i7#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi7#2fp4 i7#2fmq_x d7lat i7#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fp10 i6#2fmq_x d7lat i6#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fp9 i6#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fp8 d7lat i6#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi6#2fp5 i6#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fp4 i6#2fmq_x d6lat i6#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp10 i5#2fmq_x d6lat i5#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp9 i5#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp8 d6lat i5#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fp5 i5#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp4 i5#2fmq_x d5lat i5#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp10 i4#2fmq_x d5lat i4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp9 i4#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp8 d5lat i4#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fp5 i4#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp4 i4#2fmq_x d4lat i4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi31#2fp15 i31#2fseb sen vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmp3 db sen i31#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmp2 i31#2fnet21 d vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmp1 db i31#2fseb i31#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi31#2fmp0 i31#2fnet20 sdi vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp4 i0#2fmq_x db i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC4MSFQ_1




.subckt SAEDRVT14_SYNC4ORMSFQNS_1 vdd vss vbp vbn q ck d en setb te
xn19 ckb ckbb vss vbn n08_rev2 l=0.014u nf=2 m=1 nfin=3
xn3 db d vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
xmn1 q d8lat net031 vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmn0 net031 setb vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xi7#2fn12 i7#2fmq_x d8lat i7#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi7#2fn11 i7#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi7#2fn10 d8lat i7#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi7#2fn7 i7#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi7#2fn6 i7#2fmq_x d7lat i7#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fn12 i6#2fmq_x d7lat i6#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi6#2fn11 i6#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fn10 d7lat i6#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi6#2fn7 i6#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fn6 i6#2fmq_x d6lat i6#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn12 i5#2fmq_x d6lat i5#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fn11 i5#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn10 d6lat i5#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fn7 i5#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fn6 i5#2fmq_x d5lat i5#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn12 i4#2fmq_x d5lat i4#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn11 i4#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn10 d5lat i4#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fn7 i4#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fn6 i4#2fmq_x d4lat i4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn12 i3#2fmq_x d4lat i3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn11 i3#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn10 d4lat i3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fn7 i3#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fn6 i3#2fmq_x d3lat i3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn12 i2#2fmq_x d3lat i2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn11 i2#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn10 d3lat i2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fn7 i2#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fn6 i2#2fmq_x d2lat i2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn12 i1#2fmq_x d2lat i1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn11 i1#2fnet048 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn10 d2lat i1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fn7 i1#2fnet050 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fn6 i1#2fmq_x d1lat i1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn12 i0#2fmq_x d1lat i0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn11 i0#2fnet048 ckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn10 d1lat i0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fn7 i0#2fnet050 ckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fn6 i0#2fmq_x db i0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xck_gater#2fn24 ck_gater#2fe_nr_te te vss vbn n08 l=0.014u nf=1 m=1 nfin=3
xck_gater#2fn10 ck_gater#2fe_nr_te en vss vbn n08 l=0.014u nf=1 m=1 nfin=3
xck_gater#2fn1 ck_gater#2fckbb ck_gater#2fckb vss vbn n08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fn0 ck_gater#2fckb ck vss vbn n08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi31#2fn11 ck_gater#2fi31#2fmidn_en_ck1 ck_gater#2fqf vss vbn n08 l=0.014u nf=1 m=1 nfin=3
xck_gater#2fi31#2fn01 ck_gater#2fzn ck ck_gater#2fi31#2fmidn_en_ck1 vbn n08 l=0.014u nf=1 m=1 nfin=3
xck_gater#2fi31#2fn2 ckbb ck_gater#2fzn vss vbn n08 l=0.014u nf=4 m=1 nfin=4
xck_gater#2fi31#2fn1 ck_gater#2fi31#2fmidn_en_ck ck_gater#2fqf vss vbn n08 l=0.014u nf=1 m=1 nfin=3
xck_gater#2fi31#2fn0 ck_gater#2fzn ck ck_gater#2fi31#2fmidn_en_ck vbn n08 l=0.014u nf=1 m=1 nfin=3
xck_gater#2fi1#2fn23 ck_gater#2fi1#2fnet61 ck_gater#2fqf vss vbn n08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi1#2fn20 ck_gater#2fe_nr_te ck_gater#2fckb ck_gater#2fqf_x vbn n08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi1#2fn12 ck_gater#2fqf_x ck_gater#2fckbb ck_gater#2fi1#2fnet61 vbn n08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi1#2fn10 ck_gater#2fqf ck_gater#2fqf_x vss vbn n08 l=0.014u nf=1 m=1 nfin=2
xp17 ckb ckbb vdd vbp p08_rev2 l=0.014u nf=2 m=1 nfin=3
xp1 db d vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xmp1 q setb vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmp0 q d8lat vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xi7#2fp10 i7#2fmq_x d8lat i7#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi7#2fp9 i7#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi7#2fp8 d8lat i7#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi7#2fp5 i7#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi7#2fp4 i7#2fmq_x d7lat i7#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fp10 i6#2fmq_x d7lat i6#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fp9 i6#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fp8 d7lat i6#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi6#2fp5 i6#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi6#2fp4 i6#2fmq_x d6lat i6#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp10 i5#2fmq_x d6lat i5#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp9 i5#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp8 d6lat i5#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi5#2fp5 i5#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi5#2fp4 i5#2fmq_x d5lat i5#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp10 i4#2fmq_x d5lat i4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp9 i4#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp8 d5lat i4#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi4#2fp5 i4#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi4#2fp4 i4#2fmq_x d4lat i4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp10 i3#2fmq_x d4lat i3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp9 i3#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp8 d4lat i3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi3#2fp5 i3#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi3#2fp4 i3#2fmq_x d3lat i3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp10 i2#2fmq_x d3lat i2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp9 i2#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp8 d3lat i2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi2#2fp5 i2#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi2#2fp4 i2#2fmq_x d2lat i2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp10 i1#2fmq_x d2lat i1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp9 i1#2fnet047 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp8 d2lat i1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi1#2fp5 i1#2fnet049 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi1#2fp4 i1#2fmq_x d1lat i1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp10 i0#2fmq_x d1lat i0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp9 i0#2fnet047 ckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp8 d1lat i0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi0#2fp5 i0#2fnet049 ckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi0#2fp4 i0#2fmq_x db i0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xck_gater#2fp23 ck_gater#2fe_nr_te te ck_gater#2fnet42 vbp p08 l=0.014u nf=1 m=1 nfin=3
xck_gater#2fp22 ck_gater#2fnet42 en vdd vbp p08 l=0.014u nf=1 m=1 nfin=3
xck_gater#2fp1 ck_gater#2fckbb ck_gater#2fckb vdd vbp p08 l=0.014u nf=1 m=1 nfin=3
xck_gater#2fp0 ck_gater#2fckb ck vdd vbp p08 l=0.014u nf=1 m=1 nfin=3
xck_gater#2fi31#2fp2 ckbb ck_gater#2fzn vdd vbp p08 l=0.014u nf=4 m=1 nfin=4
xck_gater#2fi31#2fp1 ck_gater#2fzn ck vdd vbp p08 l=0.014u nf=1 m=1 nfin=4
xck_gater#2fi31#2fp0 ck_gater#2fzn ck_gater#2fqf vdd vbp p08 l=0.014u nf=2 m=1 nfin=4
xck_gater#2fi31#2fmp2 vdd ck vdd vbp p08 l=0.014u nf=1 m=1 nfin=4
xck_gater#2fi1#2fp21 ck_gater#2fqf_x ck_gater#2fckb ck_gater#2fi1#2fnet98 vbp p08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi1#2fp18 ck_gater#2fqf_x ck_gater#2fckbb ck_gater#2fe_nr_te vbp p08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi1#2fp9 ck_gater#2fi1#2fnet98 ck_gater#2fqf vdd vbp p08 l=0.014u nf=1 m=1 nfin=2
xck_gater#2fi1#2fp8 ck_gater#2fqf ck_gater#2fqf_x vdd vbp p08 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_SYNC4ORMSFQNS_1




.subckt SAEDRVT14_SYNC5CDCMSFQ_1 ckdst cksrc dsrc q qsrc sdidst sdisrc sendst sensrc vbn vbp vdd vss
xi9#2fi9#2fn7 i9#2fi9#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi9#2fn6 i9#2fi9#2fmq_x i9#2fd9lat i9#2fi9#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi8#2fn12 i9#2fi8#2fmq_x i9#2fd9lat i9#2fi8#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi8#2fn11 i9#2fi8#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi8#2fn10 i9#2fd9lat i9#2fi8#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi8#2fn7 i9#2fi8#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi8#2fn6 i9#2fi8#2fmq_x i9#2fd8lat i9#2fi8#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi7#2fn12 i9#2fi7#2fmq_x i9#2fd8lat i9#2fi7#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi7#2fn11 i9#2fi7#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi7#2fn10 i9#2fd8lat i9#2fi7#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi7#2fn7 i9#2fi7#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi7#2fn6 i9#2fi7#2fmq_x i9#2fd7lat i9#2fi7#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fn12 i9#2fi6#2fmq_x i9#2fd7lat i9#2fi6#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi6#2fn11 i9#2fi6#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fn10 i9#2fd7lat i9#2fi6#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi6#2fn7 i9#2fi6#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fn6 i9#2fi6#2fmq_x i9#2fd6lat i9#2fi6#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fn12 i9#2fi5#2fmq_x i9#2fd6lat i9#2fi5#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi5#2fn11 i9#2fi5#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fn10 i9#2fd6lat i9#2fi5#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi5#2fn7 i9#2fi5#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fn6 i9#2fi5#2fmq_x i9#2fd5lat i9#2fi5#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fn12 i9#2fi4#2fmq_x i9#2fd5lat i9#2fi4#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fn11 i9#2fi4#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fn10 i9#2fd5lat i9#2fi4#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fn7 i9#2fi4#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fn6 i9#2fi4#2fmq_x i9#2fd4lat i9#2fi4#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi31#2fn17 i9#2fi31#2fseb sendst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn3 i9#2fdb i9#2fi31#2fseb i9#2fi31#2fnet22 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn2 i9#2fi31#2fnet22 ddst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn1 i9#2fdb sendst i9#2fi31#2fnet19 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmn0 i9#2fi31#2fnet19 sdidst vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi3#2fn12 i9#2fi3#2fmq_x i9#2fd4lat i9#2fi3#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fn11 i9#2fi3#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fn10 i9#2fd4lat i9#2fi3#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fn7 i9#2fi3#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fn6 i9#2fi3#2fmq_x i9#2fd3lat i9#2fi3#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn12 i9#2fi2#2fmq_x i9#2fd3lat i9#2fi2#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fn11 i9#2fi2#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn10 i9#2fd3lat i9#2fi2#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fn7 i9#2fi2#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fn6 i9#2fi2#2fmq_x i9#2fd2lat i9#2fi2#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn12 i9#2fi1#2fmq_x i9#2fd2lat i9#2fi1#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fn11 i9#2fi1#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn10 i9#2fd2lat i9#2fi1#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fn7 i9#2fi1#2fnet050 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fn6 i9#2fi1#2fmq_x i9#2fd1lat i9#2fi1#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn12 i9#2fi0#2fmq_x i9#2fd1lat i9#2fi0#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fn11 i9#2fi0#2fnet048 i9#2fckbb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn10 i9#2fd1lat i9#2fi0#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fn7 i9#2fi0#2fnet050 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fn6 i9#2fi0#2fmq_x i9#2fdb i9#2fi0#2fnet050 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xsrcdff#2fn1 srcdff#2fckbb srcdff#2fckb vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fn0 srcdff#2fckb cksrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn13 srcdff#2fibase#2fnet046 srcdff#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn12 srcdff#2fmq srcdff#2fckbb srcdff#2fibase#2fnet048 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn11 srcdff#2fibase#2fnet048 srcdff#2fmq_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn10 srcdff#2fmq_x srcdff#2fmq vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn9 srcdff#2fqf_x srcdff#2fckb srcdff#2fibase#2fnet046 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn8 srcdff#2fqf srcdff#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn6 srcdff#2fmq srcdff#2fckb srcdff#2fibase#2fnet028 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn5 srcdff#2fmq_x srcdff#2fckbb srcdff#2fqf_x vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fn0 srcdff#2fibase#2fnet028 srcdff#2fnet050 vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi3#2fn0 ddst srcdff#2fqf_x vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi2#2fn0 srcdff_qb srcdff#2fqf vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi0#2fn17 srcdff#2fi0#2fseb sensrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn3 srcdff#2fnet050 srcdff#2fi0#2fseb srcdff#2fi0#2fnet22 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn2 srcdff#2fi0#2fnet22 dsrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn1 srcdff#2fnet050 sensrc srcdff#2fi0#2fnet19 vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmn0 srcdff#2fi0#2fnet19 sdisrc vss vbn n08_rev4 l=0.014u nf=1 m=1 nfin=2   
xn20 qsrc srcdff_qb vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xi9#2fn20 q i9#2fd10lat vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fn19 i9#2fckbb i9#2fckb vss vbn n08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi9#2fn18 i9#2fckb ckdst vss vbn n08_rev3 l=0.014u nf=3 m=1 nfin=4   
xi9#2fi9#2fn12 i9#2fi9#2fmq_x i9#2fd10lat i9#2fi9#2fnet048 vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi9#2fn11 i9#2fi9#2fnet048 i9#2fckb vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi9#2fn10 i9#2fd10lat i9#2fi9#2fmq_x vss vbn n08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi8#2fp10 i9#2fi8#2fmq_x i9#2fd9lat i9#2fi8#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi8#2fp9 i9#2fi8#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi8#2fp8 i9#2fd9lat i9#2fi8#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi8#2fp5 i9#2fi8#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi8#2fp4 i9#2fi8#2fmq_x i9#2fd8lat i9#2fi8#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi7#2fp10 i9#2fi7#2fmq_x i9#2fd8lat i9#2fi7#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi7#2fp9 i9#2fi7#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi7#2fp8 i9#2fd8lat i9#2fi7#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi7#2fp5 i9#2fi7#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi7#2fp4 i9#2fi7#2fmq_x i9#2fd7lat i9#2fi7#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fp10 i9#2fi6#2fmq_x i9#2fd7lat i9#2fi6#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fp9 i9#2fi6#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fp8 i9#2fd7lat i9#2fi6#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi6#2fp5 i9#2fi6#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi6#2fp4 i9#2fi6#2fmq_x i9#2fd6lat i9#2fi6#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp10 i9#2fi5#2fmq_x i9#2fd6lat i9#2fi5#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp9 i9#2fi5#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp8 i9#2fd6lat i9#2fi5#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi5#2fp5 i9#2fi5#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi5#2fp4 i9#2fi5#2fmq_x i9#2fd5lat i9#2fi5#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp10 i9#2fi4#2fmq_x i9#2fd5lat i9#2fi4#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp9 i9#2fi4#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp8 i9#2fd5lat i9#2fi4#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi4#2fp5 i9#2fi4#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi4#2fp4 i9#2fi4#2fmq_x i9#2fd4lat i9#2fi4#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi31#2fp15 i9#2fi31#2fseb sendst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp3 i9#2fdb sendst i9#2fi31#2fnet21 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp2 i9#2fi31#2fnet21 ddst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp1 i9#2fdb i9#2fi31#2fseb i9#2fi31#2fnet20 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi31#2fmp0 i9#2fi31#2fnet20 sdidst vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=2   
xi9#2fi3#2fp10 i9#2fi3#2fmq_x i9#2fd4lat i9#2fi3#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp9 i9#2fi3#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp8 i9#2fd4lat i9#2fi3#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi3#2fp5 i9#2fi3#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi3#2fp4 i9#2fi3#2fmq_x i9#2fd3lat i9#2fi3#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp10 i9#2fi2#2fmq_x i9#2fd3lat i9#2fi2#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp9 i9#2fi2#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp8 i9#2fd3lat i9#2fi2#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi2#2fp5 i9#2fi2#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi2#2fp4 i9#2fi2#2fmq_x i9#2fd2lat i9#2fi2#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp10 i9#2fi1#2fmq_x i9#2fd2lat i9#2fi1#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp9 i9#2fi1#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp8 i9#2fd2lat i9#2fi1#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi1#2fp5 i9#2fi1#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi1#2fp4 i9#2fi1#2fmq_x i9#2fd1lat i9#2fi1#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp10 i9#2fi0#2fmq_x i9#2fd1lat i9#2fi0#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp9 i9#2fi0#2fnet047 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp8 i9#2fd1lat i9#2fi0#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi0#2fp5 i9#2fi0#2fnet049 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi0#2fp4 i9#2fi0#2fmq_x i9#2fdb i9#2fi0#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xsrcdff#2fp1 srcdff#2fckbb srcdff#2fckb vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fp0 srcdff#2fckb cksrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp11 srcdff#2fibase#2fnet045 srcdff#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp10 srcdff#2fmq srcdff#2fckb srcdff#2fibase#2fnet047 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp9 srcdff#2fibase#2fnet047 srcdff#2fmq_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp8 srcdff#2fmq_x srcdff#2fmq vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp7 srcdff#2fqf_x srcdff#2fckbb srcdff#2fibase#2fnet045 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp6 srcdff#2fqf srcdff#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp4 srcdff#2fmq srcdff#2fckbb srcdff#2fibase#2fnet027 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp3 srcdff#2fqf_x srcdff#2fckb srcdff#2fmq_x vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fibase#2fp1 srcdff#2fibase#2fnet027 srcdff#2fnet050 vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi3#2fp1 ddst srcdff#2fqf_x vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi2#2fp1 srcdff_qb srcdff#2fqf vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=4   
xsrcdff#2fi0#2fp15 srcdff#2fi0#2fseb sensrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp3 srcdff#2fnet050 sensrc srcdff#2fi0#2fnet21 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp2 srcdff#2fi0#2fnet21 dsrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp1 srcdff#2fnet050 srcdff#2fi0#2fseb srcdff#2fi0#2fnet20 vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xsrcdff#2fi0#2fmp0 srcdff#2fi0#2fnet20 sdisrc vdd vbp p08_rev4 l=0.014u nf=1 m=1 nfin=2   
xp18 qsrc srcdff_qb vdd vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xi9#2fp18 q i9#2fd10lat vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fp17 i9#2fckbb i9#2fckb vdd vbp p08_rev3 l=0.014u nf=2 m=1 nfin=4   
xi9#2fp16 i9#2fckb ckdst vdd vbp p08_rev3 l=0.014u nf=3 m=1 nfin=4   
xi9#2fi9#2fp10 i9#2fi9#2fmq_x i9#2fd10lat i9#2fi9#2fnet047 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi9#2fp9 i9#2fi9#2fnet047 i9#2fckbb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi9#2fp8 i9#2fd10lat i9#2fi9#2fmq_x vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=4   
xi9#2fi9#2fp5 i9#2fi9#2fnet049 i9#2fckb vdd vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
xi9#2fi9#2fp4 i9#2fi9#2fmq_x i9#2fd9lat i9#2fi9#2fnet049 vbp p08_rev3 l=0.014u nf=1 m=1 nfin=3   
.ends SAEDRVT14_SYNC5CDCMSFQ_1




.subckt SAEDRVT14_TAPDS vdd vss
.ends SAEDRVT14_TAPDS




.subckt SAEDRVT14_TAPPN vdd vss
.ends SAEDRVT14_TAPPN




.subckt SAEDRVT14_TAPPP10 vdd vss vddr
.ends SAEDRVT14_TAPPP10




.subckt SAEDRVT14_TIE0_4 vdd vss vbp vbn x
xmn0 net19 net19 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn0 x net015 vss vbn n08_rev l=0.014u nf=6 m=1 nfin=3
xmp0 net015 net19 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 x net015 vdd vbp p08_rev l=0.014u nf=6 m=1 nfin=3
.ends SAEDRVT14_TIE0_4




.subckt SAEDRVT14_TIE0_PV1ECO_1 vdd vss vddr vbp vbn x
xp0 net16 net16 vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=2
xn0 x net16 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=2
.ends SAEDRVT14_TIE0_PV1ECO_1




.subckt SAEDRVT14_TIE0_V1_2 vdd vss vbp vbn x
xmn0 x net16 vss vbn n08_rev l=0.014u nf=8 m=1 nfin=4
xmp0 net16 net16 vdd vbp p08_rev l=0.014u nf=8 m=1 nfin=4
.ends SAEDRVT14_TIE0_V1_2




.subckt SAEDRVT14_TIE0_V1ECO_1 vdd vss vbp vbn x
xmn0 x net16 vss vbn n08_rev l=0.014u nf=1 m=4 nfin=4
xmp0 net16 net16 vdd vbp p08_rev l=0.014u nf=1 m=4 nfin=4
.ends SAEDRVT14_TIE0_V1ECO_1




.subckt SAEDRVT14_TIE1_4 vdd vss vbp vbn x
xmn0 net014 net16 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=4
xmmn0 x net014 vss vbn n08_rev l=0.014u nf=3 m=1 nfin=3
xmp0 net16 net16 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=4
xmmp0 x net014 vdd vbp p08_rev l=0.014u nf=3 m=1 nfin=3
.ends SAEDRVT14_TIE1_4




.subckt SAEDRVT14_TIE1_PV1ECO_1 vdd vss vddr vbp vbn x
xp0 x net19 vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 net19 net19 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_TIE1_PV1ECO_1




.subckt SAEDRVT14_TIE1_V1_2 vdd vss vbp vbn x
xmn0 net19 net19 vss vbn n08_rev l=0.014u nf=2 m=1 nfin=3
xmp0 x net19 vdd vbp p08_rev l=0.014u nf=2 m=1 nfin=3
.ends SAEDRVT14_TIE1_V1_2




.subckt SAEDRVT14_TIE1_V1ECO_1 vdd vss vbp vbn x
xmn0 net19 net19 vss vbn n08_rev l=0.014u nf=1 m=1 nfin=3
xmp0 x net19 vdd vbp p08_rev l=0.014u nf=1 m=1 nfin=3
.ends SAEDRVT14_TIE1_V1ECO_1




.subckt SAEDRVT14_TIEDIN_4 vdd vss vbp vbn x
xmn1 x int_zn vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn0 int_zn net8 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 net8 int_zn vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp0 net8 net8 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_TIEDIN_4




.subckt SAEDRVT14_TIEDIN_PV1ECO_6 vdd vss vddr vbp vbn x
xp1 net5 net9 vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xp0 net5 net5 vddr vbp p08_rev2 l=0.014u nf=1 m=1 nfin=4
xn1 x net9 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
xn0 net9 net5 vss vbn n08_rev2 l=0.014u nf=1 m=1 nfin=4
.ends SAEDRVT14_TIEDIN_PV1ECO_6




.subckt SAEDRVT14_TIEDIN_V1ECO_6 vdd vss vbp vbn x
xmn1 x net9 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmn0 net9 net5 vss vbn n08_rev l=0.014u nf=4 m=1 nfin=4
xmp1 net5 net9 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
xmp0 net5 net5 vdd vbp p08_rev l=0.014u nf=4 m=1 nfin=4
.ends SAEDRVT14_TIEDIN_V1ECO_6


