
//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  localparam stallOff = 0; 
  wire                  stall_ctrl;
  assign stall_ctrl = stallOff;

  assign idat = dat;
  assign rdy = irdy && !stall_ctrl;
  assign ivld = vld && !stall_ctrl;

endmodule


//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  localparam stallOff = 0; 
  wire stall_ctrl;
  assign stall_ctrl = stallOff;

  assign dat = idat;
  assign irdy = rdy && !stall_ctrl;
  assign vld = ivld && !stall_ctrl;

endmodule



//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ../td_ccore_solutions/leading_sign_53_0_fab32403c768e182f2743a5a858355d3a89f_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Sun Oct  6 01:34:12 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_53_0
// ------------------------------------------------------------------


module leading_sign_53_0 (
  mantissa, rtn
);
  input [52:0] mantissa;
  output [5:0] rtn;


  // Interconnect Declarations
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_18_3_sdt_3;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_42_4_sdt_4;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_62_3_sdt_3;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_90_5_sdt_5;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_110_3_sdt_3;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_134_4_sdt_4;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_14_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_34_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_58_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_78_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_106_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_126_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_23;
  wire c_h_1_24;
  wire c_h_1_25;

  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_205_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_216_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_3_nl;

  // Interconnect Declarations for Component Instantiations 
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_2
      = ~((mantissa[50:49]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_1
      = ~((mantissa[52:51]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_14_2_sdt_1
      = ~((mantissa[48:47]!=2'b00));
  assign c_h_1_2 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_2;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_18_3_sdt_3
      = (mantissa[46:45]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_14_2_sdt_1;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_2
      = ~((mantissa[42:41]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_1
      = ~((mantissa[44:43]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_34_2_sdt_1
      = ~((mantissa[40:39]!=2'b00));
  assign c_h_1_5 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_18_3_sdt_3;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_42_4_sdt_4
      = (mantissa[38:37]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_34_2_sdt_1
      & c_h_1_5;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_2
      = ~((mantissa[34:33]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_1
      = ~((mantissa[36:35]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_58_2_sdt_1
      = ~((mantissa[32:31]!=2'b00));
  assign c_h_1_9 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_2;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_62_3_sdt_3
      = (mantissa[30:29]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_58_2_sdt_1;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_2
      = ~((mantissa[26:25]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_1
      = ~((mantissa[28:27]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_78_2_sdt_1
      = ~((mantissa[24:23]!=2'b00));
  assign c_h_1_12 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_42_4_sdt_4;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_90_5_sdt_5
      = (mantissa[22:21]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_78_2_sdt_1
      & c_h_1_12 & c_h_1_13;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_2
      = ~((mantissa[18:17]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_1
      = ~((mantissa[20:19]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_106_2_sdt_1
      = ~((mantissa[16:15]!=2'b00));
  assign c_h_1_17 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_2;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_110_3_sdt_3
      = (mantissa[14:13]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_106_2_sdt_1;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_2
      = ~((mantissa[10:9]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_1
      = ~((mantissa[12:11]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_126_2_sdt_1
      = ~((mantissa[8:7]!=2'b00));
  assign c_h_1_20 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_110_3_sdt_3;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_134_4_sdt_4
      = (mantissa[6:5]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_126_2_sdt_1
      & c_h_1_20;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_2
      = ~((mantissa[2:1]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_1
      = ~((mantissa[4:3]!=2'b00));
  assign c_h_1_23 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_2;
  assign c_h_1_24 = c_h_1_21 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_25 = c_h_1_14 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_90_5_sdt_5;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_205_nl
      = c_h_1_14 & (c_h_1_24 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_90_5_sdt_5));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_nl
      = c_h_1_6 & (c_h_1_13 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_42_4_sdt_4))
      & (~((~(c_h_1_21 & (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_134_4_sdt_4)))
      & c_h_1_25));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_216_nl
      = c_h_1_2 & (c_h_1_5 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_18_3_sdt_3))
      & (~((~(c_h_1_9 & (c_h_1_12 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~((~(c_h_1_17 & (c_h_1_20 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_110_3_sdt_3))
      & (c_h_1_23 | (~ c_h_1_24)))) & c_h_1_25));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_1_nl
      = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_14_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_34_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_58_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_2))
      & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_78_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_106_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_2))
      & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_126_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_2))))
      & c_h_1_21)) & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_1
      & (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_2)))
      & c_h_1_24)))) & c_h_1_25));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_3_nl
      = ((~((mantissa[52]) | (~((mantissa[51:50]!=2'b01))))) & (~(((mantissa[48])
      | (~((mantissa[47:46]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[44]) | (~((mantissa[43:42]!=2'b01)))))
      & (~(((mantissa[40]) | (~((mantissa[39:38]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[36]) | (~((mantissa[35:34]!=2'b01))))) & (~(((mantissa[32])
      | (~((mantissa[31:30]!=2'b01)))) & c_h_1_9)) & (~((~((~((mantissa[28]) | (~((mantissa[27:26]!=2'b01)))))
      & (~(((mantissa[24]) | (~((mantissa[23:22]!=2'b01)))) & c_h_1_12)))) & c_h_1_13))))
      & c_h_1_14)) & (~((~((~((mantissa[20]) | (~((mantissa[19:18]!=2'b01))))) &
      (~(((mantissa[16]) | (~((mantissa[15:14]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[12])
      | (~((mantissa[11:10]!=2'b01))))) & (~(((mantissa[8]) | (~((mantissa[7:6]!=2'b01))))
      & c_h_1_20)))) & c_h_1_21)) & (~(((mantissa[4]) | (~((mantissa[3:2]!=2'b01)))
      | c_h_1_23) & c_h_1_24)))) & c_h_1_25))) | ((~ (mantissa[0])) & c_h_1_23 &
      c_h_1_24 & c_h_1_25);
  assign rtn = {c_h_1_25 , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_205_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_216_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_1_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_3_nl};
endmodule




//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ../td_ccore_solutions/leading_sign_57_0_1_0_8314b0004a517a8de2b01928bce9c178b0a9_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Sun Oct  6 01:34:25 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_57_0_1_0
// ------------------------------------------------------------------


module leading_sign_57_0_1_0 (
  mantissa, all_same, rtn
);
  input [56:0] mantissa;
  output all_same;
  output [5:0] rtn;


  // Interconnect Declarations
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_18_3_sdt_3;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_42_4_sdt_4;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_62_3_sdt_3;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_90_5_sdt_5;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_110_3_sdt_3;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_134_4_sdt_4;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_154_3_sdt_3;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_168_6_sdt_6;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_14_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_34_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_58_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_78_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_106_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_126_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_150_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_24;
  wire c_h_1_25;
  wire c_h_1_26;
  wire c_h_1_27;

  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_and_221_nl;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_and_219_nl;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_nl;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_or_4_nl;

  // Interconnect Declarations for Component Instantiations 
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_2 = ~((mantissa[54:53]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_1 = ~((mantissa[56:55]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_14_2_sdt_1 = ~((mantissa[52:51]!=2'b00));
  assign c_h_1_2 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_2;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_18_3_sdt_3 = (mantissa[50:49]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_14_2_sdt_1;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_2 = ~((mantissa[46:45]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_1 = ~((mantissa[48:47]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_34_2_sdt_1 = ~((mantissa[44:43]!=2'b00));
  assign c_h_1_5 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_18_3_sdt_3;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_42_4_sdt_4 = (mantissa[42:41]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_34_2_sdt_1 & c_h_1_5;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_2 = ~((mantissa[38:37]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_1 = ~((mantissa[40:39]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_58_2_sdt_1 = ~((mantissa[36:35]!=2'b00));
  assign c_h_1_9 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_2;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_62_3_sdt_3 = (mantissa[34:33]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_58_2_sdt_1;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_2 = ~((mantissa[30:29]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_1 = ~((mantissa[32:31]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_78_2_sdt_1 = ~((mantissa[28:27]!=2'b00));
  assign c_h_1_12 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_42_4_sdt_4;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_90_5_sdt_5 = (mantissa[26:25]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_78_2_sdt_1 & c_h_1_12
      & c_h_1_13;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_2 = ~((mantissa[22:21]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_1 = ~((mantissa[24:23]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_106_2_sdt_1 = ~((mantissa[20:19]!=2'b00));
  assign c_h_1_17 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_2;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_110_3_sdt_3 = (mantissa[18:17]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_106_2_sdt_1;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_2 = ~((mantissa[14:13]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_1 = ~((mantissa[16:15]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_126_2_sdt_1 = ~((mantissa[12:11]!=2'b00));
  assign c_h_1_20 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_110_3_sdt_3;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_134_4_sdt_4 = (mantissa[10:9]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_126_2_sdt_1 & c_h_1_20;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_2 = ~((mantissa[6:5]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_1 = ~((mantissa[8:7]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_150_2_sdt_1 = ~((mantissa[4:3]!=2'b00));
  assign c_h_1_24 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_2;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_154_3_sdt_3 = (mantissa[2:1]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_150_2_sdt_1;
  assign c_h_1_25 = c_h_1_24 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_154_3_sdt_3;
  assign c_h_1_26 = c_h_1_21 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_134_4_sdt_4;
  assign c_h_1_27 = c_h_1_14 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_90_5_sdt_5;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_168_6_sdt_6 = (~
      (mantissa[0])) & c_h_1_25 & c_h_1_26 & c_h_1_27;
  assign all_same = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_168_6_sdt_6;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_and_221_nl = c_h_1_14 &
      (c_h_1_26 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_90_5_sdt_5));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_and_219_nl = c_h_1_6 &
      (c_h_1_13 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_42_4_sdt_4))
      & (~((~(c_h_1_21 & (c_h_1_25 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_134_4_sdt_4))))
      & c_h_1_27));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_nl
      = c_h_1_2 & (c_h_1_5 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_18_3_sdt_3))
      & (~((~(c_h_1_9 & (c_h_1_12 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~((~(c_h_1_17 & (c_h_1_20 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_110_3_sdt_3))
      & (~((~(c_h_1_24 & (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_154_3_sdt_3)))
      & c_h_1_26)))) & c_h_1_27));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_1_nl
      = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_1 & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_14_2_sdt_1
      | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_2)) & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_34_2_sdt_1 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_58_2_sdt_1 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_2))
      & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_1 &
      (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_78_2_sdt_1 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_106_2_sdt_1 | (~
      return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_2)) & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_126_2_sdt_1 | (~
      return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_2)))) & c_h_1_21))
      & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_150_2_sdt_1 | (~
      return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_2)) & (~ c_h_1_25)))
      & c_h_1_26)))) & c_h_1_27));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_or_4_nl
      = ((~((mantissa[56]) | (~((mantissa[55:54]!=2'b01))))) & (~(((mantissa[52])
      | (~((mantissa[51:50]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[48]) | (~((mantissa[47:46]!=2'b01)))))
      & (~(((mantissa[44]) | (~((mantissa[43:42]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[40]) | (~((mantissa[39:38]!=2'b01))))) & (~(((mantissa[36])
      | (~((mantissa[35:34]!=2'b01)))) & c_h_1_9)) & (~((~((~((mantissa[32]) | (~((mantissa[31:30]!=2'b01)))))
      & (~(((mantissa[28]) | (~((mantissa[27:26]!=2'b01)))) & c_h_1_12)))) & c_h_1_13))))
      & c_h_1_14)) & (~((~((~((mantissa[24]) | (~((mantissa[23:22]!=2'b01))))) &
      (~(((mantissa[20]) | (~((mantissa[19:18]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[16])
      | (~((mantissa[15:14]!=2'b01))))) & (~(((mantissa[12]) | (~((mantissa[11:10]!=2'b01))))
      & c_h_1_20)))) & c_h_1_21)) & (~(((mantissa[8]) | (~((mantissa[7:6]!=2'b01)))
      | (((mantissa[4]) | (~((mantissa[3:2]!=2'b01)))) & c_h_1_24) | c_h_1_25) &
      c_h_1_26)))) & c_h_1_27))) | return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_168_6_sdt_6;
  assign rtn = {c_h_1_27 , return_add_generic_AC_RND_CONV_false_ls_all_sign_and_221_nl
      , return_add_generic_AC_RND_CONV_false_ls_all_sign_and_219_nl , return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_nl
      , return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_1_nl
      , return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_or_4_nl};
endmodule




//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/mgc_shift_r_beh_v5.v 
module mgc_shift_r_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

endmodule

//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_generic_reg_beh.v 

module mgc_generic_reg (d, clk, en, a_rst, s_rst, q);
   parameter width = 8;
   parameter ph_clk = 1;    //clock polarity, 1=rising_edge
   parameter ph_en = 1;
   parameter ph_a_rst = 1;  // 0 to 1 
   parameter ph_s_rst = 1;  // 0 to 1
   parameter a_rst_used = 1;
   parameter s_rst_used = 0;
   parameter en_used = 0;

   input [width-1:0]      d;
   input                  clk;
   input                  en;
   input                  a_rst;
   input                  s_rst;
   output reg [width-1:0] q;

   generate
      if (ph_clk==1 && ph_a_rst==1)
      begin: GEN_CLK1_ARST1
         always@(posedge a_rst or posedge clk)
           if (a_rst == 1'b1)
             q <= {width{1'b0}};
           else if (s_rst == $unsigned(ph_s_rst))
             q <= {width{1'b0}};
           else if (en == $unsigned(ph_en))
             q <= d;
      end //GEN_CLK1_ARST1

      else if (ph_clk==1 && ph_a_rst==0)
      begin: GEN_CLK1_ARST0
         always@(negedge a_rst or posedge clk)
           if (a_rst == 1'b0)
             q <= {width{1'b0}};
           else if (s_rst == $unsigned(ph_s_rst))
             q <= {width{1'b0}};
           else if (en == $unsigned(ph_en))
             q <= d;
      end //GEN_CLK1_ARST0

      else if (ph_clk==0 && ph_a_rst==1)
      begin: GEN_CLK0_ARST1
         always@(posedge a_rst or negedge clk)
           if (a_rst == 1'b1)
             q <= {width{1'b0}};
           else if (s_rst == $unsigned(ph_s_rst))
             q <= {width{1'b0}};
           else if (en == $unsigned(ph_en))
             q <= d;
      end //GEN_CLK0_ARST1

      else if (ph_clk==0 && ph_a_rst==0)
      begin: GEN_CLK0_ARST0
         always@(negedge a_rst or negedge clk)
           if (a_rst == 1'b0)
             q <= {width{1'b0}};
           else if (s_rst == $unsigned(ph_s_rst))
             q <= {width{1'b0}};
           else if (en == $unsigned(ph_en))
             q <= d;
      end //GEN_CLK0_ARST0

   endgenerate

endmodule

//------> ./rtl_stagemgc_rom_sync_regout_14_1024_14_1_0_0_1_0_1_0_0_0_1_60.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Sun Oct  6 01:48:34 2024
// ----------------------------------------------------------------------

// 
module stagemgc_rom_sync_regout_14_1024_14_1_0_0_1_0_1_0_0_0_1_60 (addr, data_out,
    clk, s_rst, a_rst, en
);
  input [9:0]addr ;
  output [13:0]data_out ;
  input clk ;
  input s_rst ;
  input a_rst ;
  input en ;


  // Constants for ROM dimensions
  parameter n_width    = 14;
  parameter n_size     = 1024;
  parameter n_numports = 1;
  parameter n_addr_w   = 10;
  parameter n_inreg    = 0;
  parameter n_outreg   = 1;
  wire [9:0] addr_f;

  // Build input address registers
  wire [9:0] addr_reg [n_inreg:0];
  genvar i;
  generate if (n_inreg > 0)
  begin
    for( i=n_inreg-1; i >= 1; i=i-1)
    begin: addr_reg_stage
      mgc_generic_reg #(
        .width(10), 
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_addr_reg (
        .d(addr_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(addr_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(10), 
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_addr_reg_init (
      .d(addr),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(addr_reg[0])
    );
    assign addr_f = addr_reg[n_inreg-1];
  end
  else
  begin
    assign addr_f = addr;
  end
  endgenerate

  // Declare storage for memory elements
  wire [13:0] mem [1023:0];

  // Declare output registers
  reg [13:0] data_out_t;

  // Initialize ROM contents
  assign mem[0] = 14'b00111111111011;
  assign mem[1] = 14'b01111011010000;
  assign mem[2] = 14'b10101100110100;
  assign mem[3] = 14'b10101111001000;
  assign mem[4] = 14'b01101100110000;
  assign mem[5] = 14'b01000011110110;
  assign mem[6] = 14'b01100010000011;
  assign mem[7] = 14'b10011000011111;
  assign mem[8] = 14'b00011000110111;
  assign mem[9] = 14'b01100011111111;
  assign mem[10] = 14'b10010100000101;
  assign mem[11] = 14'b01010010010010;
  assign mem[12] = 14'b00001001001010;
  assign mem[13] = 14'b01011011000001;
  assign mem[14] = 14'b01110101110010;
  assign mem[15] = 14'b10010111101110;
  assign mem[16] = 14'b00010001101110;
  assign mem[17] = 14'b01100100000111;
  assign mem[18] = 14'b00011010101111;
  assign mem[19] = 14'b00001111000101;
  assign mem[20] = 14'b01101110111011;
  assign mem[21] = 14'b01110111111010;
  assign mem[22] = 14'b00111010011111;
  assign mem[23] = 14'b01100100101010;
  assign mem[24] = 14'b10100010101110;
  assign mem[25] = 14'b01111110100100;
  assign mem[26] = 14'b00011101011101;
  assign mem[27] = 14'b00011010011000;
  assign mem[28] = 14'b00010101010100;
  assign mem[29] = 14'b10100001011001;
  assign mem[30] = 14'b10011110110100;
  assign mem[31] = 14'b10001111011100;
  assign mem[32] = 14'b10111110110010;
  assign mem[33] = 14'b01100001100000;
  assign mem[34] = 14'b00001111100101;
  assign mem[35] = 14'b00000001110101;
  assign mem[36] = 14'b01001010101111;
  assign mem[37] = 14'b01000100110111;
  assign mem[38] = 14'b00011000001101;
  assign mem[39] = 14'b01101110100000;
  assign mem[40] = 14'b00101100001101;
  assign mem[41] = 14'b01100100111010;
  assign mem[42] = 14'b01000101001111;
  assign mem[43] = 14'b10001010101101;
  assign mem[44] = 14'b01101111101000;
  assign mem[45] = 14'b00101000000100;
  assign mem[46] = 14'b01011000100000;
  assign mem[47] = 14'b00111111001010;
  assign mem[48] = 14'b10111110011101;
  assign mem[49] = 14'b00000110110000;
  assign mem[50] = 14'b10100111111111;
  assign mem[51] = 14'b00010011010101;
  assign mem[52] = 14'b01110110111010;
  assign mem[53] = 14'b00010111111110;
  assign mem[54] = 14'b00111110001111;
  assign mem[55] = 14'b01111010110111;
  assign mem[56] = 14'b00100010000101;
  assign mem[57] = 14'b01100010100100;
  assign mem[58] = 14'b10001000010000;
  assign mem[59] = 14'b01100110101010;
  assign mem[60] = 14'b01001011101011;
  assign mem[61] = 14'b00011010011010;
  assign mem[62] = 14'b00000000001110;
  assign mem[63] = 14'b00111100100000;
  assign mem[64] = 14'b01010111000001;
  assign mem[65] = 14'b10010010011000;
  assign mem[66] = 14'b10111110000011;
  assign mem[67] = 14'b00011111100011;
  assign mem[68] = 14'b01110101110111;
  assign mem[69] = 14'b00100100001011;
  assign mem[70] = 14'b01001001000001;
  assign mem[71] = 14'b01110010101100;
  assign mem[72] = 14'b00011000010001;
  assign mem[73] = 14'b00010010000100;
  assign mem[74] = 14'b10000011010001;
  assign mem[75] = 14'b10110001111101;
  assign mem[76] = 14'b00001111111100;
  assign mem[77] = 14'b00101110010111;
  assign mem[78] = 14'b10101000010100;
  assign mem[79] = 14'b01101110000101;
  assign mem[80] = 14'b00110011110100;
  assign mem[81] = 14'b10101111100100;
  assign mem[82] = 14'b01010010100101;
  assign mem[83] = 14'b10110100111010;
  assign mem[84] = 14'b10100110001101;
  assign mem[85] = 14'b10011101100110;
  assign mem[86] = 14'b10010100010101;
  assign mem[87] = 14'b01100000100100;
  assign mem[88] = 14'b10010000111101;
  assign mem[89] = 14'b01011111110010;
  assign mem[90] = 14'b00110011111011;
  assign mem[91] = 14'b00001101110011;
  assign mem[92] = 14'b10100011100101;
  assign mem[93] = 14'b00000111101001;
  assign mem[94] = 14'b00010111011110;
  assign mem[95] = 14'b00101100100011;
  assign mem[96] = 14'b10101100110101;
  assign mem[97] = 14'b10011000000001;
  assign mem[98] = 14'b00101010110110;
  assign mem[99] = 14'b10111111010001;
  assign mem[100] = 14'b01001101101010;
  assign mem[101] = 14'b10100011110001;
  assign mem[102] = 14'b10011101011110;
  assign mem[103] = 14'b00010010101011;
  assign mem[104] = 14'b00001011011010;
  assign mem[105] = 14'b00011011100010;
  assign mem[106] = 14'b00111100001110;
  assign mem[107] = 14'b00011111101110;
  assign mem[108] = 14'b01011100000100;
  assign mem[109] = 14'b10101010101010;
  assign mem[110] = 14'b10001100111100;
  assign mem[111] = 14'b01010010011010;
  assign mem[112] = 14'b10001111011011;
  assign mem[113] = 14'b00111000010100;
  assign mem[114] = 14'b00111011000110;
  assign mem[115] = 14'b10011111011110;
  assign mem[116] = 14'b00110001101100;
  assign mem[117] = 14'b00110110001011;
  assign mem[118] = 14'b01001000111100;
  assign mem[119] = 14'b00100110001110;
  assign mem[120] = 14'b01110110111101;
  assign mem[121] = 14'b10010010101010;
  assign mem[122] = 14'b00001101000010;
  assign mem[123] = 14'b01111000010111;
  assign mem[124] = 14'b01101010110100;
  assign mem[125] = 14'b00110101001011;
  assign mem[126] = 14'b01010011100111;
  assign mem[127] = 14'b10111111110100;
  assign mem[128] = 14'b00110111111100;
  assign mem[129] = 14'b00011011001011;
  assign mem[130] = 14'b10101001000100;
  assign mem[131] = 14'b10011000111011;
  assign mem[132] = 14'b10011111100001;
  assign mem[133] = 14'b00111111100110;
  assign mem[134] = 14'b10111111011010;
  assign mem[135] = 14'b10000101001101;
  assign mem[136] = 14'b10100010100001;
  assign mem[137] = 14'b00101010111101;
  assign mem[138] = 14'b01110010101010;
  assign mem[139] = 14'b10100101001110;
  assign mem[140] = 14'b01011110011000;
  assign mem[141] = 14'b00001110101111;
  assign mem[142] = 14'b10010001110010;
  assign mem[143] = 14'b00010111000101;
  assign mem[144] = 14'b01101011010001;
  assign mem[145] = 14'b10010111000100;
  assign mem[146] = 14'b00111000000001;
  assign mem[147] = 14'b01100111101001;
  assign mem[148] = 14'b10111101110001;
  assign mem[149] = 14'b00111111011111;
  assign mem[150] = 14'b00111001100100;
  assign mem[151] = 14'b01111000000000;
  assign mem[152] = 14'b01111111111100;
  assign mem[153] = 14'b01101011110110;
  assign mem[154] = 14'b00110111001101;
  assign mem[155] = 14'b10011001001111;
  assign mem[156] = 14'b01011111001010;
  assign mem[157] = 14'b00001011010111;
  assign mem[158] = 14'b10011101110011;
  assign mem[159] = 14'b01101101011011;
  assign mem[160] = 14'b01101100100001;
  assign mem[161] = 14'b00011110011101;
  assign mem[162] = 14'b10011000000011;
  assign mem[163] = 14'b10100100111111;
  assign mem[164] = 14'b01011110101001;
  assign mem[165] = 14'b00000101111010;
  assign mem[166] = 14'b01111010111111;
  assign mem[167] = 14'b10001000111011;
  assign mem[168] = 14'b10001011000101;
  assign mem[169] = 14'b10010000001101;
  assign mem[170] = 14'b10001010001110;
  assign mem[171] = 14'b01000111000111;
  assign mem[172] = 14'b10010101110101;
  assign mem[173] = 14'b10110110010000;
  assign mem[174] = 14'b01110111001110;
  assign mem[175] = 14'b10001001110101;
  assign mem[176] = 14'b01011000110000;
  assign mem[177] = 14'b01001101011100;
  assign mem[178] = 14'b01100001101011;
  assign mem[179] = 14'b10000011000100;
  assign mem[180] = 14'b10011110101100;
  assign mem[181] = 14'b10001000010011;
  assign mem[182] = 14'b00100100100101;
  assign mem[183] = 14'b00110001010111;
  assign mem[184] = 14'b00010110111011;
  assign mem[185] = 14'b01010101010100;
  assign mem[186] = 14'b10000101101001;
  assign mem[187] = 14'b01111001100111;
  assign mem[188] = 14'b00101001011001;
  assign mem[189] = 14'b00100100010000;
  assign mem[190] = 14'b10001101001100;
  assign mem[191] = 14'b01100000101100;
  assign mem[192] = 14'b00001011100001;
  assign mem[193] = 14'b00111001110010;
  assign mem[194] = 14'b01001001011011;
  assign mem[195] = 14'b01011001111001;
  assign mem[196] = 14'b10001101010110;
  assign mem[197] = 14'b00111001100111;
  assign mem[198] = 14'b00000000010000;
  assign mem[199] = 14'b00001110010010;
  assign mem[200] = 14'b01010001000010;
  assign mem[201] = 14'b10100100100011;
  assign mem[202] = 14'b01000111001000;
  assign mem[203] = 14'b00011110101100;
  assign mem[204] = 14'b00110110110101;
  assign mem[205] = 14'b10000011110100;
  assign mem[206] = 14'b01110101011100;
  assign mem[207] = 14'b01010100000101;
  assign mem[208] = 14'b10100111101101;
  assign mem[209] = 14'b00110011010001;
  assign mem[210] = 14'b01101101111101;
  assign mem[211] = 14'b00010000100100;
  assign mem[212] = 14'b00101101001111;
  assign mem[213] = 14'b01101111110100;
  assign mem[214] = 14'b10001010110111;
  assign mem[215] = 14'b01010011101101;
  assign mem[216] = 14'b01100100001001;
  assign mem[217] = 14'b10000000000101;
  assign mem[218] = 14'b00101110010010;
  assign mem[219] = 14'b01100011100111;
  assign mem[220] = 14'b01001111001000;
  assign mem[221] = 14'b01100111101010;
  assign mem[222] = 14'b01010111111001;
  assign mem[223] = 14'b00000100010110;
  assign mem[224] = 14'b00001110100100;
  assign mem[225] = 14'b10011111110101;
  assign mem[226] = 14'b10001011011111;
  assign mem[227] = 14'b01110111011010;
  assign mem[228] = 14'b00000101011111;
  assign mem[229] = 14'b10010001010010;
  assign mem[230] = 14'b00000011101101;
  assign mem[231] = 14'b01011011100010;
  assign mem[232] = 14'b01111000001100;
  assign mem[233] = 14'b00110001001010;
  assign mem[234] = 14'b10111101011110;
  assign mem[235] = 14'b01110110100010;
  assign mem[236] = 14'b00100000000101;
  assign mem[237] = 14'b10110000010101;
  assign mem[238] = 14'b00111011011010;
  assign mem[239] = 14'b01010001010100;
  assign mem[240] = 14'b01000111111010;
  assign mem[241] = 14'b00011011010100;
  assign mem[242] = 14'b10110000100100;
  assign mem[243] = 14'b00000101010100;
  assign mem[244] = 14'b00111001111111;
  assign mem[245] = 14'b01001000000110;
  assign mem[246] = 14'b00000100101100;
  assign mem[247] = 14'b10101011110001;
  assign mem[248] = 14'b01001111001110;
  assign mem[249] = 14'b10011101000001;
  assign mem[250] = 14'b10110101100000;
  assign mem[251] = 14'b10111111010111;
  assign mem[252] = 14'b01110011111101;
  assign mem[253] = 14'b10100111010011;
  assign mem[254] = 14'b01011001110010;
  assign mem[255] = 14'b01011000010110;
  assign mem[256] = 14'b00111011111011;
  assign mem[257] = 14'b01010110110001;
  assign mem[258] = 14'b00010011001000;
  assign mem[259] = 14'b10000100011100;
  assign mem[260] = 14'b10010000010101;
  assign mem[261] = 14'b00111100000101;
  assign mem[262] = 14'b00000011111010;
  assign mem[263] = 14'b10101111001001;
  assign mem[264] = 14'b01000010000001;
  assign mem[265] = 14'b01100010110110;
  assign mem[266] = 14'b10010111010000;
  assign mem[267] = 14'b10111111011110;
  assign mem[268] = 14'b01000000101000;
  assign mem[269] = 14'b00101011011010;
  assign mem[270] = 14'b00001010110100;
  assign mem[271] = 14'b10001001101000;
  assign mem[272] = 14'b01100100001010;
  assign mem[273] = 14'b01101000111110;
  assign mem[274] = 14'b10011101111001;
  assign mem[275] = 14'b10100010110010;
  assign mem[276] = 14'b00111010101111;
  assign mem[277] = 14'b01110010111100;
  assign mem[278] = 14'b10110001100001;
  assign mem[279] = 14'b10000011110001;
  assign mem[280] = 14'b01100100100101;
  assign mem[281] = 14'b00111001000100;
  assign mem[282] = 14'b01100011000110;
  assign mem[283] = 14'b10001100010010;
  assign mem[284] = 14'b01010100001111;
  assign mem[285] = 14'b00100011100000;
  assign mem[286] = 14'b01100101001100;
  assign mem[287] = 14'b01110011111000;
  assign mem[288] = 14'b10000011100010;
  assign mem[289] = 14'b10101001001000;
  assign mem[290] = 14'b10111011010010;
  assign mem[291] = 14'b01011001100101;
  assign mem[292] = 14'b00001101101100;
  assign mem[293] = 14'b01101101110110;
  assign mem[294] = 14'b00100001110111;
  assign mem[295] = 14'b00100110000100;
  assign mem[296] = 14'b00110101110010;
  assign mem[297] = 14'b10010000000001;
  assign mem[298] = 14'b10000000001110;
  assign mem[299] = 14'b01001011111010;
  assign mem[300] = 14'b01011101001100;
  assign mem[301] = 14'b00101010111010;
  assign mem[302] = 14'b01110000001010;
  assign mem[303] = 14'b00010110011010;
  assign mem[304] = 14'b01110011011101;
  assign mem[305] = 14'b10001010101111;
  assign mem[306] = 14'b10100110100101;
  assign mem[307] = 14'b10110011000001;
  assign mem[308] = 14'b01000001111100;
  assign mem[309] = 14'b00010110011000;
  assign mem[310] = 14'b10101001010000;
  assign mem[311] = 14'b01000011101000;
  assign mem[312] = 14'b10000101101101;
  assign mem[313] = 14'b00011101001011;
  assign mem[314] = 14'b10010011101110;
  assign mem[315] = 14'b00100101110000;
  assign mem[316] = 14'b00111011101000;
  assign mem[317] = 14'b10001101110100;
  assign mem[318] = 14'b00001010101110;
  assign mem[319] = 14'b01010100010001;
  assign mem[320] = 14'b00100111011011;
  assign mem[321] = 14'b01000011110011;
  assign mem[322] = 14'b01011111100011;
  assign mem[323] = 14'b00001001101011;
  assign mem[324] = 14'b00001110101001;
  assign mem[325] = 14'b00101100010010;
  assign mem[326] = 14'b01111001011111;
  assign mem[327] = 14'b00110011001111;
  assign mem[328] = 14'b00100100111011;
  assign mem[329] = 14'b01110101000000;
  assign mem[330] = 14'b01011111100000;
  assign mem[331] = 14'b01001111000000;
  assign mem[332] = 14'b00001100111000;
  assign mem[333] = 14'b10011111011100;
  assign mem[334] = 14'b10110110101010;
  assign mem[335] = 14'b00010001011001;
  assign mem[336] = 14'b00101010100111;
  assign mem[337] = 14'b10011001111000;
  assign mem[338] = 14'b00001110000000;
  assign mem[339] = 14'b00011111101100;
  assign mem[340] = 14'b01001111010011;
  assign mem[341] = 14'b00101001011110;
  assign mem[342] = 14'b10100011100000;
  assign mem[343] = 14'b01111011001100;
  assign mem[344] = 14'b10111110001001;
  assign mem[345] = 14'b01010100111010;
  assign mem[346] = 14'b00101111111110;
  assign mem[347] = 14'b01100100000000;
  assign mem[348] = 14'b10001110101100;
  assign mem[349] = 14'b10110110011000;
  assign mem[350] = 14'b10111101111001;
  assign mem[351] = 14'b01000110101000;
  assign mem[352] = 14'b00010011111001;
  assign mem[353] = 14'b10011000001011;
  assign mem[354] = 14'b10110011001100;
  assign mem[355] = 14'b10011011010001;
  assign mem[356] = 14'b10011100110111;
  assign mem[357] = 14'b10010111111000;
  assign mem[358] = 14'b00100011010110;
  assign mem[359] = 14'b10010010110111;
  assign mem[360] = 14'b10101110111000;
  assign mem[361] = 14'b00000100111011;
  assign mem[362] = 14'b01000110011111;
  assign mem[363] = 14'b00010010000110;
  assign mem[364] = 14'b01011110101101;
  assign mem[365] = 14'b01101001011111;
  assign mem[366] = 14'b10111001011001;
  assign mem[367] = 14'b00000101100101;
  assign mem[368] = 14'b01110011000111;
  assign mem[369] = 14'b01000111000110;
  assign mem[370] = 14'b00001111010111;
  assign mem[371] = 14'b10000101010110;
  assign mem[372] = 14'b10000010100000;
  assign mem[373] = 14'b10011110001110;
  assign mem[374] = 14'b01110101101010;
  assign mem[375] = 14'b10010000100101;
  assign mem[376] = 14'b01000100001111;
  assign mem[377] = 14'b01010001100101;
  assign mem[378] = 14'b00111110011111;
  assign mem[379] = 14'b10001001001001;
  assign mem[380] = 14'b00110001011001;
  assign mem[381] = 14'b01101101001110;
  assign mem[382] = 14'b01000000100010;
  assign mem[383] = 14'b10110110000100;
  assign mem[384] = 14'b00110100101110;
  assign mem[385] = 14'b10110011010101;
  assign mem[386] = 14'b00011011011001;
  assign mem[387] = 14'b00000100100100;
  assign mem[388] = 14'b10000111101001;
  assign mem[389] = 14'b00101011110110;
  assign mem[390] = 14'b10100010001010;
  assign mem[391] = 14'b10111110011100;
  assign mem[392] = 14'b01011010101000;
  assign mem[393] = 14'b10111000100011;
  assign mem[394] = 14'b00110001101101;
  assign mem[395] = 14'b00011111000100;
  assign mem[396] = 14'b00010000000000;
  assign mem[397] = 14'b10010001111100;
  assign mem[398] = 14'b00100110101101;
  assign mem[399] = 14'b10101010110000;
  assign mem[400] = 14'b01000111100110;
  assign mem[401] = 14'b01101001011110;
  assign mem[402] = 14'b00111000100011;
  assign mem[403] = 14'b01010101111111;
  assign mem[404] = 14'b01010001110001;
  assign mem[405] = 14'b00100110011111;
  assign mem[406] = 14'b10000100010110;
  assign mem[407] = 14'b01110111100010;
  assign mem[408] = 14'b01111100011100;
  assign mem[409] = 14'b01100011111011;
  assign mem[410] = 14'b00010000101111;
  assign mem[411] = 14'b00010011111000;
  assign mem[412] = 14'b00110110010010;
  assign mem[413] = 14'b10101100100101;
  assign mem[414] = 14'b00110011011011;
  assign mem[415] = 14'b10110001010000;
  assign mem[416] = 14'b10000100110110;
  assign mem[417] = 14'b10010100000110;
  assign mem[418] = 14'b10011001101101;
  assign mem[419] = 14'b00010011100101;
  assign mem[420] = 14'b00011101000001;
  assign mem[421] = 14'b01100001011001;
  assign mem[422] = 14'b01001001110000;
  assign mem[423] = 14'b10110100101001;
  assign mem[424] = 14'b01011110010010;
  assign mem[425] = 14'b10011001011001;
  assign mem[426] = 14'b00110100001011;
  assign mem[427] = 14'b00011100000101;
  assign mem[428] = 14'b00101100111111;
  assign mem[429] = 14'b01100001100010;
  assign mem[430] = 14'b01010001010000;
  assign mem[431] = 14'b00100001000010;
  assign mem[432] = 14'b01111100011010;
  assign mem[433] = 14'b10010010001001;
  assign mem[434] = 14'b10110001100011;
  assign mem[435] = 14'b01010101100011;
  assign mem[436] = 14'b01011111000100;
  assign mem[437] = 14'b10010110000001;
  assign mem[438] = 14'b01000000001100;
  assign mem[439] = 14'b01110010011011;
  assign mem[440] = 14'b10100011000110;
  assign mem[441] = 14'b10010011111111;
  assign mem[442] = 14'b00010011110111;
  assign mem[443] = 14'b00000110011000;
  assign mem[444] = 14'b01101011111111;
  assign mem[445] = 14'b00110000000111;
  assign mem[446] = 14'b00000101101000;
  assign mem[447] = 14'b10000001010100;
  assign mem[448] = 14'b10110100001111;
  assign mem[449] = 14'b10001111000100;
  assign mem[450] = 14'b10001101011001;
  assign mem[451] = 14'b10110100010011;
  assign mem[452] = 14'b00001101010010;
  assign mem[453] = 14'b10000110101001;
  assign mem[454] = 14'b00001100010000;
  assign mem[455] = 14'b01111011101111;
  assign mem[456] = 14'b10000010001110;
  assign mem[457] = 14'b10111110001010;
  assign mem[458] = 14'b00011100110110;
  assign mem[459] = 14'b10011111100101;
  assign mem[460] = 14'b10111110011000;
  assign mem[461] = 14'b01111010010011;
  assign mem[462] = 14'b10111001111111;
  assign mem[463] = 14'b01010111100000;
  assign mem[464] = 14'b10011000110011;
  assign mem[465] = 14'b00001111110100;
  assign mem[466] = 14'b00001011010001;
  assign mem[467] = 14'b00101011100000;
  assign mem[468] = 14'b01101000010100;
  assign mem[469] = 14'b01100110011000;
  assign mem[470] = 14'b01010011100100;
  assign mem[471] = 14'b01000101001000;
  assign mem[472] = 14'b01101010100000;
  assign mem[473] = 14'b10000011010101;
  assign mem[474] = 14'b10011011100111;
  assign mem[475] = 14'b01010000011110;
  assign mem[476] = 14'b00100100110100;
  assign mem[477] = 14'b01010110110000;
  assign mem[478] = 14'b01010010010011;
  assign mem[479] = 14'b00010100110101;
  assign mem[480] = 14'b10001001100001;
  assign mem[481] = 14'b10010110111101;
  assign mem[482] = 14'b01110010001100;
  assign mem[483] = 14'b01011010011100;
  assign mem[484] = 14'b01001100101110;
  assign mem[485] = 14'b00001110001101;
  assign mem[486] = 14'b10110101011101;
  assign mem[487] = 14'b01000100101011;
  assign mem[488] = 14'b10000000101110;
  assign mem[489] = 14'b01101000011110;
  assign mem[490] = 14'b01000011001110;
  assign mem[491] = 14'b00101111100100;
  assign mem[492] = 14'b00100011101101;
  assign mem[493] = 14'b10111111011001;
  assign mem[494] = 14'b00011110101011;
  assign mem[495] = 14'b10010000000000;
  assign mem[496] = 14'b01000011001000;
  assign mem[497] = 14'b10111010001110;
  assign mem[498] = 14'b00001010110111;
  assign mem[499] = 14'b01000100010011;
  assign mem[500] = 14'b10011001000001;
  assign mem[501] = 14'b01001100010100;
  assign mem[502] = 14'b00100101101011;
  assign mem[503] = 14'b10011111110110;
  assign mem[504] = 14'b00101001011010;
  assign mem[505] = 14'b00001101001001;
  assign mem[506] = 14'b00111100110010;
  assign mem[507] = 14'b10011111110111;
  assign mem[508] = 14'b01110001010000;
  assign mem[509] = 14'b10000100111001;
  assign mem[510] = 14'b10101110111100;
  assign mem[511] = 14'b01101000100000;
  assign mem[512] = 14'b00111111011011;
  assign mem[513] = 14'b01011110101100;
  assign mem[514] = 14'b00111001100110;
  assign mem[515] = 14'b01001001110010;
  assign mem[516] = 14'b10111001001101;
  assign mem[517] = 14'b01011010111000;
  assign mem[518] = 14'b01101110010010;
  assign mem[519] = 14'b01101011010100;
  assign mem[520] = 14'b10101110000001;
  assign mem[521] = 14'b01111011110110;
  assign mem[522] = 14'b01001100011110;
  assign mem[523] = 14'b10111111111100;
  assign mem[524] = 14'b01000000000110;
  assign mem[525] = 14'b00111101000100;
  assign mem[526] = 14'b00111000011010;
  assign mem[527] = 14'b01100101111101;
  assign mem[528] = 14'b01111100000010;
  assign mem[529] = 14'b01111100101110;
  assign mem[530] = 14'b10111011001001;
  assign mem[531] = 14'b01101001100011;
  assign mem[532] = 14'b00001000011001;
  assign mem[533] = 14'b01000111010010;
  assign mem[534] = 14'b00011001010111;
  assign mem[535] = 14'b10000000100011;
  assign mem[536] = 14'b10110010111101;
  assign mem[537] = 14'b01110101111000;
  assign mem[538] = 14'b00001110001010;
  assign mem[539] = 14'b10111000101000;
  assign mem[540] = 14'b10010101001100;
  assign mem[541] = 14'b10101001101010;
  assign mem[542] = 14'b10010111100111;
  assign mem[543] = 14'b00101011111111;
  assign mem[544] = 14'b10110111011000;
  assign mem[545] = 14'b01101010011101;
  assign mem[546] = 14'b01101101000011;
  assign mem[547] = 14'b00001100110011;
  assign mem[548] = 14'b10001011000111;
  assign mem[549] = 14'b01100001111111;
  assign mem[550] = 14'b10101001011011;
  assign mem[551] = 14'b00000101011100;
  assign mem[552] = 14'b01110101011010;
  assign mem[553] = 14'b10000010010011;
  assign mem[554] = 14'b01100100100111;
  assign mem[555] = 14'b00001010110110;
  assign mem[556] = 14'b00001101010100;
  assign mem[557] = 14'b01011000011011;
  assign mem[558] = 14'b00101011011101;
  assign mem[559] = 14'b00111010000100;
  assign mem[560] = 14'b10110101000101;
  assign mem[561] = 14'b00101111010000;
  assign mem[562] = 14'b00010111110011;
  assign mem[563] = 14'b10000111010011;
  assign mem[564] = 14'b01000000010010;
  assign mem[565] = 14'b10100111110010;
  assign mem[566] = 14'b00110011100111;
  assign mem[567] = 14'b01011011111101;
  assign mem[568] = 14'b00101110100010;
  assign mem[569] = 14'b01110001111001;
  assign mem[570] = 14'b10111001101100;
  assign mem[571] = 14'b10001110100011;
  assign mem[572] = 14'b10010001101011;
  assign mem[573] = 14'b10111000110110;
  assign mem[574] = 14'b00000001100010;
  assign mem[575] = 14'b00100111011110;
  assign mem[576] = 14'b00100001000100;
  assign mem[577] = 14'b01000000100011;
  assign mem[578] = 14'b10110010001111;
  assign mem[579] = 14'b00011100110100;
  assign mem[580] = 14'b00111000111101;
  assign mem[581] = 14'b00111101001100;
  assign mem[582] = 14'b01111111000101;
  assign mem[583] = 14'b00100010110000;
  assign mem[584] = 14'b10101001110111;
  assign mem[585] = 14'b01111110011100;
  assign mem[586] = 14'b10010110110011;
  assign mem[587] = 14'b01011101100101;
  assign mem[588] = 14'b01101111100100;
  assign mem[589] = 14'b10000100100000;
  assign mem[590] = 14'b00011010000110;
  assign mem[591] = 14'b00000010011111;
  assign mem[592] = 14'b10101010101011;
  assign mem[593] = 14'b01001100110110;
  assign mem[594] = 14'b00000010000000;
  assign mem[595] = 14'b01110010010000;
  assign mem[596] = 14'b00001011010101;
  assign mem[597] = 14'b10001111000101;
  assign mem[598] = 14'b01001110001110;
  assign mem[599] = 14'b01100011111001;
  assign mem[600] = 14'b00110110100110;
  assign mem[601] = 14'b01011110011011;
  assign mem[602] = 14'b10101011011100;
  assign mem[603] = 14'b01100000100101;
  assign mem[604] = 14'b10111000111110;
  assign mem[605] = 14'b00110101011111;
  assign mem[606] = 14'b10100100010010;
  assign mem[607] = 14'b01110111110100;
  assign mem[608] = 14'b00111001101101;
  assign mem[609] = 14'b01101000000010;
  assign mem[610] = 14'b01101011111001;
  assign mem[611] = 14'b10111010110001;
  assign mem[612] = 14'b10011111100100;
  assign mem[613] = 14'b10111010010010;
  assign mem[614] = 14'b10001110001101;
  assign mem[615] = 14'b10000010101101;
  assign mem[616] = 14'b01001111110110;
  assign mem[617] = 14'b00000000101101;
  assign mem[618] = 14'b00100101100000;
  assign mem[619] = 14'b00011110000001;
  assign mem[620] = 14'b01000100011001;
  assign mem[621] = 14'b00101010100000;
  assign mem[622] = 14'b00011010011111;
  assign mem[623] = 14'b00000000110011;
  assign mem[624] = 14'b00101011111000;
  assign mem[625] = 14'b00001010001010;
  assign mem[626] = 14'b00011101101000;
  assign mem[627] = 14'b10011100001101;
  assign mem[628] = 14'b10011011110011;
  assign mem[629] = 14'b10111011001100;
  assign mem[630] = 14'b01111110100010;
  assign mem[631] = 14'b01001011100001;
  assign mem[632] = 14'b01000000100111;
  assign mem[633] = 14'b01000010100001;
  assign mem[634] = 14'b01011011001110;
  assign mem[635] = 14'b01001010011101;
  assign mem[636] = 14'b10101011101001;
  assign mem[637] = 14'b10110100001100;
  assign mem[638] = 14'b00001001001110;
  assign mem[639] = 14'b10111110100110;
  assign mem[640] = 14'b00000111100010;
  assign mem[641] = 14'b10111110001101;
  assign mem[642] = 14'b00011111010110;
  assign mem[643] = 14'b01101110011000;
  assign mem[644] = 14'b10011100100010;
  assign mem[645] = 14'b00111101001000;
  assign mem[646] = 14'b10111011110000;
  assign mem[647] = 14'b10100100010111;
  assign mem[648] = 14'b10110001100010;
  assign mem[649] = 14'b01101100101010;
  assign mem[650] = 14'b00100010100010;
  assign mem[651] = 14'b00000100011100;
  assign mem[652] = 14'b01010100100101;
  assign mem[653] = 14'b01100111001001;
  assign mem[654] = 14'b00111100011001;
  assign mem[655] = 14'b10100001100011;
  assign mem[656] = 14'b10101110110100;
  assign mem[657] = 14'b01100001010111;
  assign mem[658] = 14'b00001000000101;
  assign mem[659] = 14'b10010101011100;
  assign mem[660] = 14'b10110000010001;
  assign mem[661] = 14'b00111100010111;
  assign mem[662] = 14'b00010010111010;
  assign mem[663] = 14'b01000111111100;
  assign mem[664] = 14'b01111111100000;
  assign mem[665] = 14'b10110010110111;
  assign mem[666] = 14'b00000010011001;
  assign mem[667] = 14'b01110000100100;
  assign mem[668] = 14'b01011010000011;
  assign mem[669] = 14'b01001111100001;
  assign mem[670] = 14'b10010000100000;
  assign mem[671] = 14'b10111101111010;
  assign mem[672] = 14'b10110111100100;
  assign mem[673] = 14'b00010101001010;
  assign mem[674] = 14'b01101000010000;
  assign mem[675] = 14'b00000010110011;
  assign mem[676] = 14'b01010110011100;
  assign mem[677] = 14'b00101001010110;
  assign mem[678] = 14'b01011100110101;
  assign mem[679] = 14'b10111110011001;
  assign mem[680] = 14'b00001101011110;
  assign mem[681] = 14'b00110001010110;
  assign mem[682] = 14'b00000111011101;
  assign mem[683] = 14'b01110001101111;
  assign mem[684] = 14'b01011000101110;
  assign mem[685] = 14'b01111011101010;
  assign mem[686] = 14'b01000010011110;
  assign mem[687] = 14'b00000100101110;
  assign mem[688] = 14'b00101101001101;
  assign mem[689] = 14'b10011110000010;
  assign mem[690] = 14'b01101011101010;
  assign mem[691] = 14'b10010101011000;
  assign mem[692] = 14'b10010110101111;
  assign mem[693] = 14'b10111010000001;
  assign mem[694] = 14'b01000000000010;
  assign mem[695] = 14'b10011001100000;
  assign mem[696] = 14'b10100000011101;
  assign mem[697] = 14'b00010101001001;
  assign mem[698] = 14'b10100111011011;
  assign mem[699] = 14'b01010011001101;
  assign mem[700] = 14'b01100001101110;
  assign mem[701] = 14'b00111101101111;
  assign mem[702] = 14'b00011100001111;
  assign mem[703] = 14'b01100100110001;
  assign mem[704] = 14'b01010000100111;
  assign mem[705] = 14'b00010100011100;
  assign mem[706] = 14'b10000001111011;
  assign mem[707] = 14'b00110101001100;
  assign mem[708] = 14'b00011101010101;
  assign mem[709] = 14'b00010011001111;
  assign mem[710] = 14'b00000001110000;
  assign mem[711] = 14'b01100011111110;
  assign mem[712] = 14'b10110111001100;
  assign mem[713] = 14'b10111111110000;
  assign mem[714] = 14'b01110001110110;
  assign mem[715] = 14'b00010110110011;
  assign mem[716] = 14'b10111111110010;
  assign mem[717] = 14'b10011010101000;
  assign mem[718] = 14'b00110110000000;
  assign mem[719] = 14'b00001100100000;
  assign mem[720] = 14'b00010101110101;
  assign mem[721] = 14'b10100110110110;
  assign mem[722] = 14'b00000001100111;
  assign mem[723] = 14'b01110011111100;
  assign mem[724] = 14'b01111100101000;
  assign mem[725] = 14'b00001110101000;
  assign mem[726] = 14'b00001011111100;
  assign mem[727] = 14'b00001001111000;
  assign mem[728] = 14'b01111100111100;
  assign mem[729] = 14'b10000000011111;
  assign mem[730] = 14'b10000011111101;
  assign mem[731] = 14'b01111001001110;
  assign mem[732] = 14'b10101001110110;
  assign mem[733] = 14'b10010101100011;
  assign mem[734] = 14'b00100111001100;
  assign mem[735] = 14'b00011110011010;
  assign mem[736] = 14'b01100101111100;
  assign mem[737] = 14'b10011110101110;
  assign mem[738] = 14'b00010000010100;
  assign mem[739] = 14'b01000011110010;
  assign mem[740] = 14'b00100110011001;
  assign mem[741] = 14'b00111000111001;
  assign mem[742] = 14'b00011001111011;
  assign mem[743] = 14'b01000000101011;
  assign mem[744] = 14'b01001001010000;
  assign mem[745] = 14'b10011000000101;
  assign mem[746] = 14'b10101110001100;
  assign mem[747] = 14'b00111101101010;
  assign mem[748] = 14'b00100000100010;
  assign mem[749] = 14'b01010010001101;
  assign mem[750] = 14'b00011111110100;
  assign mem[751] = 14'b10111001001010;
  assign mem[752] = 14'b01110111010100;
  assign mem[753] = 14'b10111111001100;
  assign mem[754] = 14'b01010011110110;
  assign mem[755] = 14'b00100101001100;
  assign mem[756] = 14'b00010101110111;
  assign mem[757] = 14'b01111000101000;
  assign mem[758] = 14'b00100000110100;
  assign mem[759] = 14'b00110010010001;
  assign mem[760] = 14'b10101010100000;
  assign mem[761] = 14'b10001011000010;
  assign mem[762] = 14'b01110110011010;
  assign mem[763] = 14'b10111011011011;
  assign mem[764] = 14'b00101011100111;
  assign mem[765] = 14'b00010010111111;
  assign mem[766] = 14'b00110100011011;
  assign mem[767] = 14'b00101010010111;
  assign mem[768] = 14'b00100011011011;
  assign mem[769] = 14'b00011111010100;
  assign mem[770] = 14'b10000101111000;
  assign mem[771] = 14'b10011111000000;
  assign mem[772] = 14'b00110010001110;
  assign mem[773] = 14'b00100100100001;
  assign mem[774] = 14'b00011011010110;
  assign mem[775] = 14'b01001001111001;
  assign mem[776] = 14'b01001110000101;
  assign mem[777] = 14'b01110011110111;
  assign mem[778] = 14'b01100010101011;
  assign mem[779] = 14'b10111100001100;
  assign mem[780] = 14'b01000100010110;
  assign mem[781] = 14'b01101111110101;
  assign mem[782] = 14'b01001011101100;
  assign mem[783] = 14'b00000011010011;
  assign mem[784] = 14'b01111101000011;
  assign mem[785] = 14'b10011110101111;
  assign mem[786] = 14'b10010001001010;
  assign mem[787] = 14'b10110011011001;
  assign mem[788] = 14'b00011011000111;
  assign mem[789] = 14'b00100100100000;
  assign mem[790] = 14'b01011010100001;
  assign mem[791] = 14'b10011010010011;
  assign mem[792] = 14'b10000000000000;
  assign mem[793] = 14'b00001111011010;
  assign mem[794] = 14'b01110101100111;
  assign mem[795] = 14'b00010101111001;
  assign mem[796] = 14'b00001101100110;
  assign mem[797] = 14'b00111000011111;
  assign mem[798] = 14'b10000100010001;
  assign mem[799] = 14'b00101011000100;
  assign mem[800] = 14'b10011000101010;
  assign mem[801] = 14'b00011111110010;
  assign mem[802] = 14'b10011110111000;
  assign mem[803] = 14'b00110011000000;
  assign mem[804] = 14'b01011111110100;
  assign mem[805] = 14'b00000000110110;
  assign mem[806] = 14'b00101101000000;
  assign mem[807] = 14'b01001010011011;
  assign mem[808] = 14'b10111000011101;
  assign mem[809] = 14'b00110000000010;
  assign mem[810] = 14'b10000001011110;
  assign mem[811] = 14'b10010011010100;
  assign mem[812] = 14'b01001100010001;
  assign mem[813] = 14'b01101100010101;
  assign mem[814] = 14'b00010001000010;
  assign mem[815] = 14'b10011100110110;
  assign mem[816] = 14'b00101000000111;
  assign mem[817] = 14'b00001011000100;
  assign mem[818] = 14'b00001101111101;
  assign mem[819] = 14'b01100101000001;
  assign mem[820] = 14'b01001101100010;
  assign mem[821] = 14'b10011100101000;
  assign mem[822] = 14'b00100000101010;
  assign mem[823] = 14'b01011001010110;
  assign mem[824] = 14'b10100111110111;
  assign mem[825] = 14'b00001100001100;
  assign mem[826] = 14'b01001001111101;
  assign mem[827] = 14'b01001000001111;
  assign mem[828] = 14'b00100001010110;
  assign mem[829] = 14'b00100000100111;
  assign mem[830] = 14'b01001011000010;
  assign mem[831] = 14'b00001101110100;
  assign mem[832] = 14'b01010011111100;
  assign mem[833] = 14'b01011010100011;
  assign mem[834] = 14'b01011100110010;
  assign mem[835] = 14'b01000011101101;
  assign mem[836] = 14'b01100110011111;
  assign mem[837] = 14'b01110101111101;
  assign mem[838] = 14'b01010010010101;
  assign mem[839] = 14'b10100110101000;
  assign mem[840] = 14'b01000010011100;
  assign mem[841] = 14'b00110010111100;
  assign mem[842] = 14'b01011100011101;
  assign mem[843] = 14'b10101000111110;
  assign mem[844] = 14'b01011010001000;
  assign mem[845] = 14'b10011011111111;
  assign mem[846] = 14'b01111110100000;
  assign mem[847] = 14'b01111001101111;
  assign mem[848] = 14'b01101010010000;
  assign mem[849] = 14'b01110101000011;
  assign mem[850] = 14'b01100010000000;
  assign mem[851] = 14'b00011101110011;
  assign mem[852] = 14'b10101011000011;
  assign mem[853] = 14'b01100010010001;
  assign mem[854] = 14'b10111000011011;
  assign mem[855] = 14'b01011110010000;
  assign mem[856] = 14'b10110010111001;
  assign mem[857] = 14'b00010010010011;
  assign mem[858] = 14'b10001111110001;
  assign mem[859] = 14'b01111011111101;
  assign mem[860] = 14'b00100110101111;
  assign mem[861] = 14'b01111100100010;
  assign mem[862] = 14'b10110001001001;
  assign mem[863] = 14'b01101110010110;
  assign mem[864] = 14'b10001011001111;
  assign mem[865] = 14'b01101001001000;
  assign mem[866] = 14'b01100110001110;
  assign mem[867] = 14'b01111110110010;
  assign mem[868] = 14'b10001001111100;
  assign mem[869] = 14'b01100111000011;
  assign mem[870] = 14'b00110111011001;
  assign mem[871] = 14'b01000011111100;
  assign mem[872] = 14'b01001000000010;
  assign mem[873] = 14'b00100010011101;
  assign mem[874] = 14'b01101101010111;
  assign mem[875] = 14'b01111110101010;
  assign mem[876] = 14'b01010110111000;
  assign mem[877] = 14'b10100010010110;
  assign mem[878] = 14'b10010001101001;
  assign mem[879] = 14'b00100111000011;
  assign mem[880] = 14'b00100101101101;
  assign mem[881] = 14'b01110001101000;
  assign mem[882] = 14'b01101011100001;
  assign mem[883] = 14'b10100101010110;
  assign mem[884] = 14'b10010001011100;
  assign mem[885] = 14'b10010011011101;
  assign mem[886] = 14'b00110111100010;
  assign mem[887] = 14'b00110011111110;
  assign mem[888] = 14'b01011101100111;
  assign mem[889] = 14'b10111011000001;
  assign mem[890] = 14'b00110101010111;
  assign mem[891] = 14'b10111111111011;
  assign mem[892] = 14'b10011001101110;
  assign mem[893] = 14'b10111100011111;
  assign mem[894] = 14'b01000011101100;
  assign mem[895] = 14'b01111010010110;
  assign mem[896] = 14'b10110001000001;
  assign mem[897] = 14'b01100111001101;
  assign mem[898] = 14'b10111111101111;
  assign mem[899] = 14'b00011111111100;
  assign mem[900] = 14'b10110101011011;
  assign mem[901] = 14'b01110010111001;
  assign mem[902] = 14'b10101111000001;
  assign mem[903] = 14'b10110100111110;
  assign mem[904] = 14'b00111010010101;
  assign mem[905] = 14'b10001011101111;
  assign mem[906] = 14'b10011011111010;
  assign mem[907] = 14'b00011001011011;
  assign mem[908] = 14'b01110000000000;
  assign mem[909] = 14'b00111101011111;
  assign mem[910] = 14'b01001110111010;
  assign mem[911] = 14'b00101011001010;
  assign mem[912] = 14'b01110101001000;
  assign mem[913] = 14'b10100010001111;
  assign mem[914] = 14'b00001011110011;
  assign mem[915] = 14'b00011001110110;
  assign mem[916] = 14'b10111100010101;
  assign mem[917] = 14'b01001101011000;
  assign mem[918] = 14'b10011110010110;
  assign mem[919] = 14'b01000100101010;
  assign mem[920] = 14'b01100111000000;
  assign mem[921] = 14'b01111011011010;
  assign mem[922] = 14'b01110101001001;
  assign mem[923] = 14'b10001011001000;
  assign mem[924] = 14'b10111011111101;
  assign mem[925] = 14'b00110111111101;
  assign mem[926] = 14'b10100111111100;
  assign mem[927] = 14'b01011000101010;
  assign mem[928] = 14'b10100001110110;
  assign mem[929] = 14'b01001100100101;
  assign mem[930] = 14'b01110011110110;
  assign mem[931] = 14'b10001001000011;
  assign mem[932] = 14'b00001011000110;
  assign mem[933] = 14'b01101001101100;
  assign mem[934] = 14'b10000100001110;
  assign mem[935] = 14'b01110000011001;
  assign mem[936] = 14'b01010011111011;
  assign mem[937] = 14'b01110001101010;
  assign mem[938] = 14'b10101101001100;
  assign mem[939] = 14'b00000100100010;
  assign mem[940] = 14'b01111010111000;
  assign mem[941] = 14'b01101010101011;
  assign mem[942] = 14'b10111000101110;
  assign mem[943] = 14'b00100111001101;
  assign mem[944] = 14'b01100110110010;
  assign mem[945] = 14'b00111110111010;
  assign mem[946] = 14'b01011010101111;
  assign mem[947] = 14'b00010110110010;
  assign mem[948] = 14'b01011001011001;
  assign mem[949] = 14'b01011010000010;
  assign mem[950] = 14'b01000001010010;
  assign mem[951] = 14'b00100000111001;
  assign mem[952] = 14'b10110101100101;
  assign mem[953] = 14'b01001011110100;
  assign mem[954] = 14'b10001011000001;
  assign mem[955] = 14'b00101100101000;
  assign mem[956] = 14'b10110011110110;
  assign mem[957] = 14'b10010000110000;
  assign mem[958] = 14'b00100111011000;
  assign mem[959] = 14'b10001001001000;
  assign mem[960] = 14'b01101101100011;
  assign mem[961] = 14'b00101001010111;
  assign mem[962] = 14'b00011101101010;
  assign mem[963] = 14'b01101101111111;
  assign mem[964] = 14'b01011100111110;
  assign mem[965] = 14'b10101110011011;
  assign mem[966] = 14'b01010101110000;
  assign mem[967] = 14'b01100010000101;
  assign mem[968] = 14'b10001111011110;
  assign mem[969] = 14'b10110011000000;
  assign mem[970] = 14'b00001001111001;
  assign mem[971] = 14'b10011100111110;
  assign mem[972] = 14'b10110100100010;
  assign mem[973] = 14'b01011000000001;
  assign mem[974] = 14'b10010101110011;
  assign mem[975] = 14'b00100100011101;
  assign mem[976] = 14'b01101101100000;
  assign mem[977] = 14'b01101110101100;
  assign mem[978] = 14'b01001110110111;
  assign mem[979] = 14'b01110000011111;
  assign mem[980] = 14'b10011010001001;
  assign mem[981] = 14'b10001100100101;
  assign mem[982] = 14'b00001000111001;
  assign mem[983] = 14'b01100011110110;
  assign mem[984] = 14'b10101001011101;
  assign mem[985] = 14'b10010111001111;
  assign mem[986] = 14'b10000001001100;
  assign mem[987] = 14'b10110011010000;
  assign mem[988] = 14'b01000001101011;
  assign mem[989] = 14'b00011111001101;
  assign mem[990] = 14'b00000000000010;
  assign mem[991] = 14'b10010001110011;
  assign mem[992] = 14'b00000010100010;
  assign mem[993] = 14'b01100000100110;
  assign mem[994] = 14'b00011111010000;
  assign mem[995] = 14'b00111001000001;
  assign mem[996] = 14'b10011001000000;
  assign mem[997] = 14'b01100011011011;
  assign mem[998] = 14'b01110110000101;
  assign mem[999] = 14'b01100000101011;
  assign mem[1000] = 14'b10000100111110;
  assign mem[1001] = 14'b10011011001111;
  assign mem[1002] = 14'b01010110100000;
  assign mem[1003] = 14'b10001100111011;
  assign mem[1004] = 14'b00111001111010;
  assign mem[1005] = 14'b10111011101001;
  assign mem[1006] = 14'b00010110101100;
  assign mem[1007] = 14'b00101111111011;
  assign mem[1008] = 14'b01010101110110;
  assign mem[1009] = 14'b10010111011100;
  assign mem[1010] = 14'b01001100000001;
  assign mem[1011] = 14'b01011110000011;
  assign mem[1012] = 14'b01101111000010;
  assign mem[1013] = 14'b10010110001010;
  assign mem[1014] = 14'b01000111101100;
  assign mem[1015] = 14'b10011110110101;
  assign mem[1016] = 14'b01100001110101;
  assign mem[1017] = 14'b01011011111111;
  assign mem[1018] = 14'b00101001011100;
  assign mem[1019] = 14'b10011110111100;
  assign mem[1020] = 14'b00011000101100;
  assign mem[1021] = 14'b10100010001011;
  assign mem[1022] = 14'b01001000011110;
  assign mem[1023] = 14'b10011011011101;

  always@(*)
  begin
    data_out_t <= mem[addr_f];
  end

  // Build output registers
  wire [13:0] data_out_reg [n_outreg:0];
  generate if (n_outreg > 0)
  begin
    for( i=n_outreg-1; i >= 1; i=i-1)
    begin: data_out_reg_stage
      mgc_generic_reg #(
        .width(14), 
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_data_out_reg (
        .d(data_out_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(data_out_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(14), 
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_data_out_reg_init (
      .d(data_out_t),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(data_out_reg[0])
    );
    assign data_out = data_out_reg[n_outreg-1];
  end
  else
  begin
    assign data_out = data_out_t;
  end
  endgenerate

endmodule



//------> ./rtl_stagemgc_rom_sync_regout_13_1024_14_1_0_0_1_0_1_0_0_0_1_60.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Sun Oct  6 01:48:34 2024
// ----------------------------------------------------------------------

// 
module stagemgc_rom_sync_regout_13_1024_14_1_0_0_1_0_1_0_0_0_1_60 (addr, data_out,
    clk, s_rst, a_rst, en
);
  input [9:0]addr ;
  output [13:0]data_out ;
  input clk ;
  input s_rst ;
  input a_rst ;
  input en ;


  // Constants for ROM dimensions
  parameter n_width    = 14;
  parameter n_size     = 1024;
  parameter n_numports = 1;
  parameter n_addr_w   = 10;
  parameter n_inreg    = 0;
  parameter n_outreg   = 1;
  wire [9:0] addr_f;

  // Build input address registers
  wire [9:0] addr_reg [n_inreg:0];
  genvar i;
  generate if (n_inreg > 0)
  begin
    for( i=n_inreg-1; i >= 1; i=i-1)
    begin: addr_reg_stage
      mgc_generic_reg #(
        .width(10), 
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_addr_reg (
        .d(addr_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(addr_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(10), 
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_addr_reg_init (
      .d(addr),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(addr_reg[0])
    );
    assign addr_f = addr_reg[n_inreg-1];
  end
  else
  begin
    assign addr_f = addr;
  end
  endgenerate

  // Declare storage for memory elements
  wire [13:0] mem [1023:0];

  // Declare output registers
  reg [13:0] data_out_t;

  // Initialize ROM contents
  assign mem[0] = 14'b00111111111011;
  assign mem[1] = 14'b01000100110001;
  assign mem[2] = 14'b00010000111001;
  assign mem[3] = 14'b00010011001101;
  assign mem[4] = 14'b00100111100010;
  assign mem[5] = 14'b01011101111110;
  assign mem[6] = 14'b01111100001011;
  assign mem[7] = 14'b01010011010001;
  assign mem[8] = 14'b00101000010011;
  assign mem[9] = 14'b01001010001111;
  assign mem[10] = 14'b01100101000000;
  assign mem[11] = 14'b10110110110111;
  assign mem[12] = 14'b01101101101111;
  assign mem[13] = 14'b00101011111100;
  assign mem[14] = 14'b01011100000010;
  assign mem[15] = 14'b10100111001010;
  assign mem[16] = 14'b00110000100101;
  assign mem[17] = 14'b00100001001101;
  assign mem[18] = 14'b00011110101000;
  assign mem[19] = 14'b10101010101101;
  assign mem[20] = 14'b10100101101001;
  assign mem[21] = 14'b10100010100100;
  assign mem[22] = 14'b01000001011101;
  assign mem[23] = 14'b00011101010011;
  assign mem[24] = 14'b01011011010111;
  assign mem[25] = 14'b10000101100010;
  assign mem[26] = 14'b01001000000111;
  assign mem[27] = 14'b01010001000110;
  assign mem[28] = 14'b10110000111100;
  assign mem[29] = 14'b10100101010010;
  assign mem[30] = 14'b01011011111010;
  assign mem[31] = 14'b10101110010011;
  assign mem[32] = 14'b10000011100001;
  assign mem[33] = 14'b10111111110011;
  assign mem[34] = 14'b10100101100111;
  assign mem[35] = 14'b01110100010110;
  assign mem[36] = 14'b01011001010111;
  assign mem[37] = 14'b00110111110001;
  assign mem[38] = 14'b01011101011101;
  assign mem[39] = 14'b10011101111100;
  assign mem[40] = 14'b01000101001010;
  assign mem[41] = 14'b10000001110010;
  assign mem[42] = 14'b10101000000011;
  assign mem[43] = 14'b01001001000111;
  assign mem[44] = 14'b10101100101100;
  assign mem[45] = 14'b00011000000010;
  assign mem[46] = 14'b10111001010001;
  assign mem[47] = 14'b00000001100100;
  assign mem[48] = 14'b10000000110111;
  assign mem[49] = 14'b01100111100001;
  assign mem[50] = 14'b10010111111101;
  assign mem[51] = 14'b01010000011001;
  assign mem[52] = 14'b00110101010100;
  assign mem[53] = 14'b01111010110010;
  assign mem[54] = 14'b01011011000111;
  assign mem[55] = 14'b10010011110100;
  assign mem[56] = 14'b01010001100001;
  assign mem[57] = 14'b10100111110100;
  assign mem[58] = 14'b01111011001010;
  assign mem[59] = 14'b01110101010010;
  assign mem[60] = 14'b10111110001100;
  assign mem[61] = 14'b10110000011100;
  assign mem[62] = 14'b01011110100001;
  assign mem[63] = 14'b00000001001111;
  assign mem[64] = 14'b00000000001101;
  assign mem[65] = 14'b01101100011010;
  assign mem[66] = 14'b10001010110110;
  assign mem[67] = 14'b01010101001101;
  assign mem[68] = 14'b01000111101010;
  assign mem[69] = 14'b10110010111111;
  assign mem[70] = 14'b00101101010111;
  assign mem[71] = 14'b01001001000100;
  assign mem[72] = 14'b10011001110011;
  assign mem[73] = 14'b01110111000101;
  assign mem[74] = 14'b10001001110110;
  assign mem[75] = 14'b10001110010101;
  assign mem[76] = 14'b00100000100011;
  assign mem[77] = 14'b10000100111011;
  assign mem[78] = 14'b10000111101101;
  assign mem[79] = 14'b00110000100110;
  assign mem[80] = 14'b01101101100111;
  assign mem[81] = 14'b00110011000101;
  assign mem[82] = 14'b00010101010111;
  assign mem[83] = 14'b01100011111101;
  assign mem[84] = 14'b10100000010011;
  assign mem[85] = 14'b10000011110011;
  assign mem[86] = 14'b10100100011111;
  assign mem[87] = 14'b10110100100111;
  assign mem[88] = 14'b10101101010110;
  assign mem[89] = 14'b00100010100011;
  assign mem[90] = 14'b00011100010000;
  assign mem[91] = 14'b01110010010111;
  assign mem[92] = 14'b00000000110000;
  assign mem[93] = 14'b10010101001011;
  assign mem[94] = 14'b00101000000000;
  assign mem[95] = 14'b00010011001100;
  assign mem[96] = 14'b10010011011110;
  assign mem[97] = 14'b10101000100011;
  assign mem[98] = 14'b10111000011000;
  assign mem[99] = 14'b00011100011100;
  assign mem[100] = 14'b10110010001110;
  assign mem[101] = 14'b10001100000110;
  assign mem[102] = 14'b01100000001111;
  assign mem[103] = 14'b00101111000100;
  assign mem[104] = 14'b01011111011101;
  assign mem[105] = 14'b00101011101100;
  assign mem[106] = 14'b00100010011011;
  assign mem[107] = 14'b00011001110100;
  assign mem[108] = 14'b00001011000111;
  assign mem[109] = 14'b01101101011100;
  assign mem[110] = 14'b00010000011101;
  assign mem[111] = 14'b10001100001101;
  assign mem[112] = 14'b01010001111100;
  assign mem[113] = 14'b00010111101101;
  assign mem[114] = 14'b10010001101010;
  assign mem[115] = 14'b10110000000101;
  assign mem[116] = 14'b00001110000100;
  assign mem[117] = 14'b00111100110000;
  assign mem[118] = 14'b10101101111101;
  assign mem[119] = 14'b10100111110000;
  assign mem[120] = 14'b01001101010101;
  assign mem[121] = 14'b01110111000000;
  assign mem[122] = 14'b10011011110110;
  assign mem[123] = 14'b01001010001010;
  assign mem[124] = 14'b10100000011110;
  assign mem[125] = 14'b00000001111110;
  assign mem[126] = 14'b00101101101001;
  assign mem[127] = 14'b01101001000000;
  assign mem[128] = 14'b01100111101011;
  assign mem[129] = 14'b01100110001111;
  assign mem[130] = 14'b00011000101110;
  assign mem[131] = 14'b01001100000100;
  assign mem[132] = 14'b00000000101010;
  assign mem[133] = 14'b00001010100001;
  assign mem[134] = 14'b00100011000000;
  assign mem[135] = 14'b01110000110011;
  assign mem[136] = 14'b00010100010000;
  assign mem[137] = 14'b10111011010101;
  assign mem[138] = 14'b01110111111011;
  assign mem[139] = 14'b10000110000010;
  assign mem[140] = 14'b10111010101101;
  assign mem[141] = 14'b00001111011101;
  assign mem[142] = 14'b10100100101101;
  assign mem[143] = 14'b01111000000111;
  assign mem[144] = 14'b01101110101101;
  assign mem[145] = 14'b10000100100111;
  assign mem[146] = 14'b00001111101100;
  assign mem[147] = 14'b10011111111100;
  assign mem[148] = 14'b01001001011111;
  assign mem[149] = 14'b00000010100011;
  assign mem[150] = 14'b10001110110111;
  assign mem[151] = 14'b01000111110101;
  assign mem[152] = 14'b01100100011111;
  assign mem[153] = 14'b10111100010100;
  assign mem[154] = 14'b00101110101111;
  assign mem[155] = 14'b10111010100010;
  assign mem[156] = 14'b01001000100111;
  assign mem[157] = 14'b00110100100010;
  assign mem[158] = 14'b00100000001100;
  assign mem[159] = 14'b10110001011101;
  assign mem[160] = 14'b10111011101011;
  assign mem[161] = 14'b01101000001000;
  assign mem[162] = 14'b01011000010111;
  assign mem[163] = 14'b01110000111001;
  assign mem[164] = 14'b01011100011010;
  assign mem[165] = 14'b10010001101111;
  assign mem[166] = 14'b00111111111100;
  assign mem[167] = 14'b01011011111000;
  assign mem[168] = 14'b01101100010100;
  assign mem[169] = 14'b00110101001010;
  assign mem[170] = 14'b01010000001101;
  assign mem[171] = 14'b10010010110010;
  assign mem[172] = 14'b10101111011101;
  assign mem[173] = 14'b01010010000100;
  assign mem[174] = 14'b10001100110000;
  assign mem[175] = 14'b00011000010100;
  assign mem[176] = 14'b01101011111100;
  assign mem[177] = 14'b01001010100101;
  assign mem[178] = 14'b00111100001101;
  assign mem[179] = 14'b10001001001100;
  assign mem[180] = 14'b10100001010101;
  assign mem[181] = 14'b01111000111001;
  assign mem[182] = 14'b00011011011110;
  assign mem[183] = 14'b01101110111111;
  assign mem[184] = 14'b10110001101111;
  assign mem[185] = 14'b10111111110001;
  assign mem[186] = 14'b10000110011010;
  assign mem[187] = 14'b00110010101011;
  assign mem[188] = 14'b01100110001000;
  assign mem[189] = 14'b01110110100110;
  assign mem[190] = 14'b10000110001111;
  assign mem[191] = 14'b10110100100000;
  assign mem[192] = 14'b01011111010101;
  assign mem[193] = 14'b00110010110101;
  assign mem[194] = 14'b10011011110001;
  assign mem[195] = 14'b10010110101000;
  assign mem[196] = 14'b01000110011010;
  assign mem[197] = 14'b00111010011000;
  assign mem[198] = 14'b01101010101101;
  assign mem[199] = 14'b10101001000110;
  assign mem[200] = 14'b10001110101010;
  assign mem[201] = 14'b10011011011100;
  assign mem[202] = 14'b00110111101110;
  assign mem[203] = 14'b00100001010101;
  assign mem[204] = 14'b00111100111101;
  assign mem[205] = 14'b01011110010110;
  assign mem[206] = 14'b01110010100101;
  assign mem[207] = 14'b01100111010001;
  assign mem[208] = 14'b00110110001100;
  assign mem[209] = 14'b01001000110011;
  assign mem[210] = 14'b00001001110001;
  assign mem[211] = 14'b00101010001100;
  assign mem[212] = 14'b01111000111010;
  assign mem[213] = 14'b00110101110011;
  assign mem[214] = 14'b00101111110100;
  assign mem[215] = 14'b00110100111100;
  assign mem[216] = 14'b00110111000110;
  assign mem[217] = 14'b01000101000010;
  assign mem[218] = 14'b10111010000111;
  assign mem[219] = 14'b01100001011000;
  assign mem[220] = 14'b00011011000010;
  assign mem[221] = 14'b00100111111110;
  assign mem[222] = 14'b10100001100100;
  assign mem[223] = 14'b01010011100000;
  assign mem[224] = 14'b01010010100110;
  assign mem[225] = 14'b00100010001110;
  assign mem[226] = 14'b10110100101010;
  assign mem[227] = 14'b01100000110111;
  assign mem[228] = 14'b00100110110010;
  assign mem[229] = 14'b10001000110100;
  assign mem[230] = 14'b01010100001011;
  assign mem[231] = 14'b01000000000101;
  assign mem[232] = 14'b01001000000001;
  assign mem[233] = 14'b10000110011101;
  assign mem[234] = 14'b10000000100010;
  assign mem[235] = 14'b00000010010000;
  assign mem[236] = 14'b01011000011000;
  assign mem[237] = 14'b10001000000000;
  assign mem[238] = 14'b00101000111101;
  assign mem[239] = 14'b01010100110000;
  assign mem[240] = 14'b10101000111100;
  assign mem[241] = 14'b00101110001111;
  assign mem[242] = 14'b10110001010010;
  assign mem[243] = 14'b01100001101001;
  assign mem[244] = 14'b00011010110011;
  assign mem[245] = 14'b01001101010111;
  assign mem[246] = 14'b10010101000100;
  assign mem[247] = 14'b00011101100000;
  assign mem[248] = 14'b00111010110100;
  assign mem[249] = 14'b00000000100111;
  assign mem[250] = 14'b10000000011011;
  assign mem[251] = 14'b00100000100000;
  assign mem[252] = 14'b00100111000110;
  assign mem[253] = 14'b00010110111101;
  assign mem[254] = 14'b10100100110110;
  assign mem[255] = 14'b10001000000101;
  assign mem[256] = 14'b01010111100001;
  assign mem[257] = 14'b00010001000101;
  assign mem[258] = 14'b00111011001000;
  assign mem[259] = 14'b01001110110001;
  assign mem[260] = 14'b00100000001010;
  assign mem[261] = 14'b10000011001111;
  assign mem[262] = 14'b10110010111000;
  assign mem[263] = 14'b10010110100111;
  assign mem[264] = 14'b00100000001011;
  assign mem[265] = 14'b10011010010110;
  assign mem[266] = 14'b01110011101101;
  assign mem[267] = 14'b00100111000000;
  assign mem[268] = 14'b01111011101110;
  assign mem[269] = 14'b10110101001010;
  assign mem[270] = 14'b00000101110011;
  assign mem[271] = 14'b01111100111001;
  assign mem[272] = 14'b00110000000001;
  assign mem[273] = 14'b10100001010110;
  assign mem[274] = 14'b00000000101000;
  assign mem[275] = 14'b10011100010100;
  assign mem[276] = 14'b10010000011101;
  assign mem[277] = 14'b01111100110011;
  assign mem[278] = 14'b01010111100011;
  assign mem[279] = 14'b00111111010011;
  assign mem[280] = 14'b01111011010110;
  assign mem[281] = 14'b00001010100100;
  assign mem[282] = 14'b10110001110100;
  assign mem[283] = 14'b01110011010011;
  assign mem[284] = 14'b01100101100101;
  assign mem[285] = 14'b01001101110101;
  assign mem[286] = 14'b00101001000100;
  assign mem[287] = 14'b00110110100000;
  assign mem[288] = 14'b10101011001100;
  assign mem[289] = 14'b01101101101110;
  assign mem[290] = 14'b01101001010001;
  assign mem[291] = 14'b10011011001101;
  assign mem[292] = 14'b01101111100011;
  assign mem[293] = 14'b00100100011010;
  assign mem[294] = 14'b00111100101100;
  assign mem[295] = 14'b01010101100001;
  assign mem[296] = 14'b01111010111001;
  assign mem[297] = 14'b01101100011101;
  assign mem[298] = 14'b01011001101001;
  assign mem[299] = 14'b01010111101101;
  assign mem[300] = 14'b10010100100001;
  assign mem[301] = 14'b10110100110000;
  assign mem[302] = 14'b10110000001101;
  assign mem[303] = 14'b00100111001110;
  assign mem[304] = 14'b01101000100001;
  assign mem[305] = 14'b00000110000010;
  assign mem[306] = 14'b01000101101110;
  assign mem[307] = 14'b00000001101001;
  assign mem[308] = 14'b00100000011100;
  assign mem[309] = 14'b10100011001011;
  assign mem[310] = 14'b00000001110111;
  assign mem[311] = 14'b00111101110011;
  assign mem[312] = 14'b01000100010010;
  assign mem[313] = 14'b10110011110001;
  assign mem[314] = 14'b00111001011000;
  assign mem[315] = 14'b10110010101111;
  assign mem[316] = 14'b00001011101110;
  assign mem[317] = 14'b00110010101000;
  assign mem[318] = 14'b00110000111101;
  assign mem[319] = 14'b00001011110010;
  assign mem[320] = 14'b00111110101101;
  assign mem[321] = 14'b10111010011001;
  assign mem[322] = 14'b10001111111010;
  assign mem[323] = 14'b01010100000010;
  assign mem[324] = 14'b10111001101001;
  assign mem[325] = 14'b10101100001010;
  assign mem[326] = 14'b00101100000010;
  assign mem[327] = 14'b00011100111011;
  assign mem[328] = 14'b01001101100110;
  assign mem[329] = 14'b01111111110101;
  assign mem[330] = 14'b00101010000000;
  assign mem[331] = 14'b01100000111101;
  assign mem[332] = 14'b01101010011110;
  assign mem[333] = 14'b00001110011110;
  assign mem[334] = 14'b00101101111000;
  assign mem[335] = 14'b01000011100111;
  assign mem[336] = 14'b10011110111111;
  assign mem[337] = 14'b01101110110001;
  assign mem[338] = 14'b01011110011111;
  assign mem[339] = 14'b10010011000010;
  assign mem[340] = 14'b10100011111100;
  assign mem[341] = 14'b10001011110110;
  assign mem[342] = 14'b00100110101000;
  assign mem[343] = 14'b01100001101111;
  assign mem[344] = 14'b00001011011000;
  assign mem[345] = 14'b01110110010001;
  assign mem[346] = 14'b01011110101000;
  assign mem[347] = 14'b10100011000000;
  assign mem[348] = 14'b10101100011100;
  assign mem[349] = 14'b00100110010100;
  assign mem[350] = 14'b00101011111011;
  assign mem[351] = 14'b00111011001011;
  assign mem[352] = 14'b00001110110001;
  assign mem[353] = 14'b10001100100110;
  assign mem[354] = 14'b00010011011100;
  assign mem[355] = 14'b10001001101111;
  assign mem[356] = 14'b10101100001001;
  assign mem[357] = 14'b10101111010010;
  assign mem[358] = 14'b01011100000110;
  assign mem[359] = 14'b01000011100101;
  assign mem[360] = 14'b01001000011111;
  assign mem[361] = 14'b00111011101011;
  assign mem[362] = 14'b10011001100010;
  assign mem[363] = 14'b01101110010000;
  assign mem[364] = 14'b01101010000010;
  assign mem[365] = 14'b10000111011110;
  assign mem[366] = 14'b01010110100011;
  assign mem[367] = 14'b01111000011011;
  assign mem[368] = 14'b00010101010001;
  assign mem[369] = 14'b10011001010100;
  assign mem[370] = 14'b00101110000101;
  assign mem[371] = 14'b10110000000001;
  assign mem[372] = 14'b10100000111101;
  assign mem[373] = 14'b10001110010100;
  assign mem[374] = 14'b00000111011110;
  assign mem[375] = 14'b01100101011001;
  assign mem[376] = 14'b00000001100101;
  assign mem[377] = 14'b00011101110111;
  assign mem[378] = 14'b10010100001011;
  assign mem[379] = 14'b00111000011000;
  assign mem[380] = 14'b10111011011101;
  assign mem[381] = 14'b10100100101000;
  assign mem[382] = 14'b00001100101100;
  assign mem[383] = 14'b10001011010011;
  assign mem[384] = 14'b00001001111101;
  assign mem[385] = 14'b01111111011111;
  assign mem[386] = 14'b01010010110011;
  assign mem[387] = 14'b10001110101000;
  assign mem[388] = 14'b00110110111000;
  assign mem[389] = 14'b10000001100010;
  assign mem[390] = 14'b01101110011100;
  assign mem[391] = 14'b01111011110010;
  assign mem[392] = 14'b00101111011100;
  assign mem[393] = 14'b01001010010111;
  assign mem[394] = 14'b00100001110011;
  assign mem[395] = 14'b00111101100001;
  assign mem[396] = 14'b00111010101011;
  assign mem[397] = 14'b10110000101010;
  assign mem[398] = 14'b01111000111011;
  assign mem[399] = 14'b01001100111010;
  assign mem[400] = 14'b10111010011100;
  assign mem[401] = 14'b00000110101000;
  assign mem[402] = 14'b01010110100010;
  assign mem[403] = 14'b01100001010100;
  assign mem[404] = 14'b10101101111011;
  assign mem[405] = 14'b01111001100010;
  assign mem[406] = 14'b10111011000110;
  assign mem[407] = 14'b00010001001001;
  assign mem[408] = 14'b00101101001010;
  assign mem[409] = 14'b10011100101011;
  assign mem[410] = 14'b00101000001001;
  assign mem[411] = 14'b00100011001010;
  assign mem[412] = 14'b00100100110000;
  assign mem[413] = 14'b00001100110101;
  assign mem[414] = 14'b00100111110110;
  assign mem[415] = 14'b10101100001000;
  assign mem[416] = 14'b01111001011001;
  assign mem[417] = 14'b00000010001000;
  assign mem[418] = 14'b00001001101001;
  assign mem[419] = 14'b00110001010101;
  assign mem[420] = 14'b01011100000001;
  assign mem[421] = 14'b10010000000011;
  assign mem[422] = 14'b01101011000111;
  assign mem[423] = 14'b00000001111000;
  assign mem[424] = 14'b01000100110101;
  assign mem[425] = 14'b00011100100001;
  assign mem[426] = 14'b10010110100011;
  assign mem[427] = 14'b01110000101110;
  assign mem[428] = 14'b10100000010101;
  assign mem[429] = 14'b10110010000001;
  assign mem[430] = 14'b00100110001001;
  assign mem[431] = 14'b10010101011010;
  assign mem[432] = 14'b10101110101000;
  assign mem[433] = 14'b00001001010111;
  assign mem[434] = 14'b00100000100101;
  assign mem[435] = 14'b10110011001001;
  assign mem[436] = 14'b01110001000001;
  assign mem[437] = 14'b01100000100001;
  assign mem[438] = 14'b01001011000001;
  assign mem[439] = 14'b10011011000110;
  assign mem[440] = 14'b10001100110010;
  assign mem[441] = 14'b01000110100010;
  assign mem[442] = 14'b10010011101111;
  assign mem[443] = 14'b10110001011000;
  assign mem[444] = 14'b10110110010110;
  assign mem[445] = 14'b01100000011110;
  assign mem[446] = 14'b01111100001110;
  assign mem[447] = 14'b10011000100110;
  assign mem[448] = 14'b01101011110000;
  assign mem[449] = 14'b10110101010011;
  assign mem[450] = 14'b00110010001101;
  assign mem[451] = 14'b10000100011001;
  assign mem[452] = 14'b10011010010001;
  assign mem[453] = 14'b00101100010011;
  assign mem[454] = 14'b10100010110110;
  assign mem[455] = 14'b00111010010100;
  assign mem[456] = 14'b01111100011001;
  assign mem[457] = 14'b00010110110001;
  assign mem[458] = 14'b10101001101001;
  assign mem[459] = 14'b01111110000101;
  assign mem[460] = 14'b00001101000000;
  assign mem[461] = 14'b00011001011100;
  assign mem[462] = 14'b00110101010010;
  assign mem[463] = 14'b01001100100100;
  assign mem[464] = 14'b10101001100111;
  assign mem[465] = 14'b01001111110111;
  assign mem[466] = 14'b10010101000111;
  assign mem[467] = 14'b01100010110101;
  assign mem[468] = 14'b01110100000111;
  assign mem[469] = 14'b00111111110011;
  assign mem[470] = 14'b00110000000000;
  assign mem[471] = 14'b10001010001111;
  assign mem[472] = 14'b10011001111101;
  assign mem[473] = 14'b10011110001010;
  assign mem[474] = 14'b01010010001011;
  assign mem[475] = 14'b10110010010101;
  assign mem[476] = 14'b01100110011100;
  assign mem[477] = 14'b00000100101111;
  assign mem[478] = 14'b00010110111001;
  assign mem[479] = 14'b00111100011111;
  assign mem[480] = 14'b01001100001001;
  assign mem[481] = 14'b01011010110101;
  assign mem[482] = 14'b10011100100001;
  assign mem[483] = 14'b01101011110010;
  assign mem[484] = 14'b00110011101111;
  assign mem[485] = 14'b01011100111011;
  assign mem[486] = 14'b10000110111101;
  assign mem[487] = 14'b01011011011100;
  assign mem[488] = 14'b00111100010000;
  assign mem[489] = 14'b00001110100000;
  assign mem[490] = 14'b01001101000101;
  assign mem[491] = 14'b10000101010010;
  assign mem[492] = 14'b00011101001111;
  assign mem[493] = 14'b00100010001000;
  assign mem[494] = 14'b01010111000011;
  assign mem[495] = 14'b01011011110111;
  assign mem[496] = 14'b00110110011001;
  assign mem[497] = 14'b10110101001101;
  assign mem[498] = 14'b10010100100111;
  assign mem[499] = 14'b01111111011001;
  assign mem[500] = 14'b00000000100011;
  assign mem[501] = 14'b00101000110001;
  assign mem[502] = 14'b01011101001011;
  assign mem[503] = 14'b01111110000000;
  assign mem[504] = 14'b00010000111000;
  assign mem[505] = 14'b10111100000111;
  assign mem[506] = 14'b10000011111100;
  assign mem[507] = 14'b00101111101100;
  assign mem[508] = 14'b00111011100101;
  assign mem[509] = 14'b10101100111001;
  assign mem[510] = 14'b01101001010000;
  assign mem[511] = 14'b10000100000110;
  assign mem[512] = 14'b00100100100100;
  assign mem[513] = 14'b01110111100011;
  assign mem[514] = 14'b00011101110110;
  assign mem[515] = 14'b10100111010101;
  assign mem[516] = 14'b00100001000101;
  assign mem[517] = 14'b10010110100101;
  assign mem[518] = 14'b01100100000010;
  assign mem[519] = 14'b01011110001100;
  assign mem[520] = 14'b00100001001100;
  assign mem[521] = 14'b01111000010101;
  assign mem[522] = 14'b00101001110111;
  assign mem[523] = 14'b01010000111111;
  assign mem[524] = 14'b01100001111110;
  assign mem[525] = 14'b01110100000000;
  assign mem[526] = 14'b00101000100101;
  assign mem[527] = 14'b01101010001011;
  assign mem[528] = 14'b10010000000110;
  assign mem[529] = 14'b10101001010101;
  assign mem[530] = 14'b00000100011000;
  assign mem[531] = 14'b10000110000111;
  assign mem[532] = 14'b00110011000110;
  assign mem[533] = 14'b01101001100001;
  assign mem[534] = 14'b00100100110010;
  assign mem[535] = 14'b00111011000011;
  assign mem[536] = 14'b01011111010110;
  assign mem[537] = 14'b01001001111100;
  assign mem[538] = 14'b01011100100110;
  assign mem[539] = 14'b00100111000001;
  assign mem[540] = 14'b10000111000000;
  assign mem[541] = 14'b10100000110001;
  assign mem[542] = 14'b01011111011011;
  assign mem[543] = 14'b10111101011111;
  assign mem[544] = 14'b00101110001110;
  assign mem[545] = 14'b10111111111111;
  assign mem[546] = 14'b10100000110100;
  assign mem[547] = 14'b01111110010110;
  assign mem[548] = 14'b00001100110001;
  assign mem[549] = 14'b00111110110101;
  assign mem[550] = 14'b00101000110010;
  assign mem[551] = 14'b00010110100100;
  assign mem[552] = 14'b01011100001011;
  assign mem[553] = 14'b10110111001000;
  assign mem[554] = 14'b00110011011100;
  assign mem[555] = 14'b00100101111000;
  assign mem[556] = 14'b01001111100010;
  assign mem[557] = 14'b01110001001010;
  assign mem[558] = 14'b01010001010101;
  assign mem[559] = 14'b01010010100001;
  assign mem[560] = 14'b10011011100100;
  assign mem[561] = 14'b00101010001110;
  assign mem[562] = 14'b01101000000000;
  assign mem[563] = 14'b00001011011111;
  assign mem[564] = 14'b00100011000011;
  assign mem[565] = 14'b10110110001000;
  assign mem[566] = 14'b00001101000001;
  assign mem[567] = 14'b00110000100011;
  assign mem[568] = 14'b01011101111100;
  assign mem[569] = 14'b01101010010001;
  assign mem[570] = 14'b00010001100110;
  assign mem[571] = 14'b01100011000011;
  assign mem[572] = 14'b01010010000010;
  assign mem[573] = 14'b10100010010111;
  assign mem[574] = 14'b10010110101010;
  assign mem[575] = 14'b01010010011110;
  assign mem[576] = 14'b00110110111001;
  assign mem[577] = 14'b10011000101001;
  assign mem[578] = 14'b00101111010001;
  assign mem[579] = 14'b00001100001011;
  assign mem[580] = 14'b10010011011001;
  assign mem[581] = 14'b00110101000000;
  assign mem[582] = 14'b01110100001101;
  assign mem[583] = 14'b00001010011100;
  assign mem[584] = 14'b10011111001000;
  assign mem[585] = 14'b01111110101111;
  assign mem[586] = 14'b01100101111111;
  assign mem[587] = 14'b01100110101000;
  assign mem[588] = 14'b10101001001111;
  assign mem[589] = 14'b01100101010010;
  assign mem[590] = 14'b10000001000111;
  assign mem[591] = 14'b01011001001111;
  assign mem[592] = 14'b10011000110100;
  assign mem[593] = 14'b00000111010011;
  assign mem[594] = 14'b01010101010110;
  assign mem[595] = 14'b01000101001001;
  assign mem[596] = 14'b10111011011111;
  assign mem[597] = 14'b00010010110101;
  assign mem[598] = 14'b01001110010111;
  assign mem[599] = 14'b01101100000110;
  assign mem[600] = 14'b01001111101000;
  assign mem[601] = 14'b00111011110011;
  assign mem[602] = 14'b01010110010101;
  assign mem[603] = 14'b10110100111011;
  assign mem[604] = 14'b00110110111110;
  assign mem[605] = 14'b01001100001011;
  assign mem[606] = 14'b01110011011100;
  assign mem[607] = 14'b00011110001011;
  assign mem[608] = 14'b01100111010111;
  assign mem[609] = 14'b00011000000101;
  assign mem[610] = 14'b10001000000100;
  assign mem[611] = 14'b00000100000100;
  assign mem[612] = 14'b00110100111001;
  assign mem[613] = 14'b01001010111000;
  assign mem[614] = 14'b01000100100111;
  assign mem[615] = 14'b01011001000001;
  assign mem[616] = 14'b01111011010111;
  assign mem[617] = 14'b00100001101011;
  assign mem[618] = 14'b01110010101001;
  assign mem[619] = 14'b00000011101100;
  assign mem[620] = 14'b10100110001011;
  assign mem[621] = 14'b10110100001110;
  assign mem[622] = 14'b00011101110010;
  assign mem[623] = 14'b01001010111001;
  assign mem[624] = 14'b10010100110111;
  assign mem[625] = 14'b01110001000111;
  assign mem[626] = 14'b10000010100010;
  assign mem[627] = 14'b01010000000001;
  assign mem[628] = 14'b10100110100110;
  assign mem[629] = 14'b00100100000111;
  assign mem[630] = 14'b00110100010010;
  assign mem[631] = 14'b10000101101100;
  assign mem[632] = 14'b00001011000011;
  assign mem[633] = 14'b00010001000000;
  assign mem[634] = 14'b01001101001000;
  assign mem[635] = 14'b00001010100110;
  assign mem[636] = 14'b10100000000101;
  assign mem[637] = 14'b00000000010010;
  assign mem[638] = 14'b01011000110100;
  assign mem[639] = 14'b00001111000000;
  assign mem[640] = 14'b01000101101011;
  assign mem[641] = 14'b01111100010101;
  assign mem[642] = 14'b00000011100010;
  assign mem[643] = 14'b00100110010011;
  assign mem[644] = 14'b00000000000110;
  assign mem[645] = 14'b10001010101010;
  assign mem[646] = 14'b00000101000000;
  assign mem[647] = 14'b01100010011010;
  assign mem[648] = 14'b10001100000011;
  assign mem[649] = 14'b10001000011111;
  assign mem[650] = 14'b00101100100100;
  assign mem[651] = 14'b00101110100101;
  assign mem[652] = 14'b00011010101011;
  assign mem[653] = 14'b01010100100000;
  assign mem[654] = 14'b01001110011001;
  assign mem[655] = 14'b10011010010100;
  assign mem[656] = 14'b10011000111110;
  assign mem[657] = 14'b00101110011000;
  assign mem[658] = 14'b00011101101011;
  assign mem[659] = 14'b01101001001001;
  assign mem[660] = 14'b01000001010111;
  assign mem[661] = 14'b01010010101010;
  assign mem[662] = 14'b10011101100100;
  assign mem[663] = 14'b01110111111111;
  assign mem[664] = 14'b01111100000101;
  assign mem[665] = 14'b10001000101000;
  assign mem[666] = 14'b01011000111110;
  assign mem[667] = 14'b00110110000101;
  assign mem[668] = 14'b01000001001111;
  assign mem[669] = 14'b01011001110011;
  assign mem[670] = 14'b01010110111001;
  assign mem[671] = 14'b00110100110010;
  assign mem[672] = 14'b01010001101011;
  assign mem[673] = 14'b00001110111000;
  assign mem[674] = 14'b01000011011111;
  assign mem[675] = 14'b10011001010010;
  assign mem[676] = 14'b01000100000100;
  assign mem[677] = 14'b00110000010000;
  assign mem[678] = 14'b10101101101110;
  assign mem[679] = 14'b00001101001000;
  assign mem[680] = 14'b01100001110001;
  assign mem[681] = 14'b00000111100110;
  assign mem[682] = 14'b01011101110000;
  assign mem[683] = 14'b00010100111110;
  assign mem[684] = 14'b10100010001110;
  assign mem[685] = 14'b01011110000001;
  assign mem[686] = 14'b01001010111110;
  assign mem[687] = 14'b01010101110001;
  assign mem[688] = 14'b01000110010010;
  assign mem[689] = 14'b01000001100001;
  assign mem[690] = 14'b00100100000010;
  assign mem[691] = 14'b01100101111001;
  assign mem[692] = 14'b00010111000011;
  assign mem[693] = 14'b01100011100100;
  assign mem[694] = 14'b10001101000101;
  assign mem[695] = 14'b01111101100101;
  assign mem[696] = 14'b00011001011001;
  assign mem[697] = 14'b01101101101100;
  assign mem[698] = 14'b01001010000100;
  assign mem[699] = 14'b01011001100010;
  assign mem[700] = 14'b01111100010100;
  assign mem[701] = 14'b01100011001111;
  assign mem[702] = 14'b01100101011110;
  assign mem[703] = 14'b01101100000101;
  assign mem[704] = 14'b10110010001101;
  assign mem[705] = 14'b01110100111111;
  assign mem[706] = 14'b10011111011010;
  assign mem[707] = 14'b10011110101011;
  assign mem[708] = 14'b01110111110010;
  assign mem[709] = 14'b01110110000100;
  assign mem[710] = 14'b10110011110101;
  assign mem[711] = 14'b00011000001010;
  assign mem[712] = 14'b01100110101011;
  assign mem[713] = 14'b10011111010111;
  assign mem[714] = 14'b00100011011001;
  assign mem[715] = 14'b01110010011111;
  assign mem[716] = 14'b01011011000000;
  assign mem[717] = 14'b10110010000100;
  assign mem[718] = 14'b10110100111101;
  assign mem[719] = 14'b10010111111010;
  assign mem[720] = 14'b00100011001011;
  assign mem[721] = 14'b10101110111111;
  assign mem[722] = 14'b01010011101100;
  assign mem[723] = 14'b01110011110000;
  assign mem[724] = 14'b00101100101101;
  assign mem[725] = 14'b00111110100011;
  assign mem[726] = 14'b10001111111111;
  assign mem[727] = 14'b00000111100100;
  assign mem[728] = 14'b01110101100110;
  assign mem[729] = 14'b10010011000001;
  assign mem[730] = 14'b10111111001011;
  assign mem[731] = 14'b01100000001101;
  assign mem[732] = 14'b10001101000001;
  assign mem[733] = 14'b00100001001001;
  assign mem[734] = 14'b10100000001111;
  assign mem[735] = 14'b00100111010111;
  assign mem[736] = 14'b10010100111101;
  assign mem[737] = 14'b00111011110000;
  assign mem[738] = 14'b10000111100010;
  assign mem[739] = 14'b10110010011011;
  assign mem[740] = 14'b10101010001000;
  assign mem[741] = 14'b01001010011010;
  assign mem[742] = 14'b10110000100111;
  assign mem[743] = 14'b01000000000001;
  assign mem[744] = 14'b00100101101110;
  assign mem[745] = 14'b01100101100000;
  assign mem[746] = 14'b10011011100001;
  assign mem[747] = 14'b10100100111010;
  assign mem[748] = 14'b00001100101000;
  assign mem[749] = 14'b00101110110111;
  assign mem[750] = 14'b00100001010010;
  assign mem[751] = 14'b01000010111110;
  assign mem[752] = 14'b10111100101110;
  assign mem[753] = 14'b01110100010101;
  assign mem[754] = 14'b01010000001100;
  assign mem[755] = 14'b01111011101011;
  assign mem[756] = 14'b00000011110101;
  assign mem[757] = 14'b01011101010110;
  assign mem[758] = 14'b01001100001010;
  assign mem[759] = 14'b01110001111100;
  assign mem[760] = 14'b01110110001000;
  assign mem[761] = 14'b10100100101011;
  assign mem[762] = 14'b10011011100000;
  assign mem[763] = 14'b10001101110011;
  assign mem[764] = 14'b00100001000001;
  assign mem[765] = 14'b00111010001001;
  assign mem[766] = 14'b10100000101101;
  assign mem[767] = 14'b10011100100110;
  assign mem[768] = 14'b10010101101010;
  assign mem[769] = 14'b10001011100110;
  assign mem[770] = 14'b10101101000010;
  assign mem[771] = 14'b10010100011010;
  assign mem[772] = 14'b00000100100110;
  assign mem[773] = 14'b01001001100111;
  assign mem[774] = 14'b00110100111111;
  assign mem[775] = 14'b00010101100001;
  assign mem[776] = 14'b10001101110000;
  assign mem[777] = 14'b10011111001101;
  assign mem[778] = 14'b01000111011001;
  assign mem[779] = 14'b10101010001010;
  assign mem[780] = 14'b10011010110101;
  assign mem[781] = 14'b01101100001011;
  assign mem[782] = 14'b00000000110101;
  assign mem[783] = 14'b01001000101101;
  assign mem[784] = 14'b00000110110111;
  assign mem[785] = 14'b10100000001101;
  assign mem[786] = 14'b01101101110100;
  assign mem[787] = 14'b10011111011111;
  assign mem[788] = 14'b10000010010111;
  assign mem[789] = 14'b00010001110101;
  assign mem[790] = 14'b00100111111100;
  assign mem[791] = 14'b01110110110001;
  assign mem[792] = 14'b01111111010110;
  assign mem[793] = 14'b10100110000110;
  assign mem[794] = 14'b10000111001000;
  assign mem[795] = 14'b10011001101000;
  assign mem[796] = 14'b01111100001111;
  assign mem[797] = 14'b10101111101101;
  assign mem[798] = 14'b00100001010011;
  assign mem[799] = 14'b01011010000101;
  assign mem[800] = 14'b10100001100111;
  assign mem[801] = 14'b10011000110101;
  assign mem[802] = 14'b00101010011110;
  assign mem[803] = 14'b00010110001011;
  assign mem[804] = 14'b01000110110011;
  assign mem[805] = 14'b00111100000100;
  assign mem[806] = 14'b00111111100010;
  assign mem[807] = 14'b01000011000101;
  assign mem[808] = 14'b10110110001001;
  assign mem[809] = 14'b10110100000101;
  assign mem[810] = 14'b10110001011001;
  assign mem[811] = 14'b01000011011001;
  assign mem[812] = 14'b01001100000101;
  assign mem[813] = 14'b10111110011010;
  assign mem[814] = 14'b00011001001011;
  assign mem[815] = 14'b10101010001100;
  assign mem[816] = 14'b10110011100001;
  assign mem[817] = 14'b10001010000001;
  assign mem[818] = 14'b00100101011001;
  assign mem[819] = 14'b00000000001111;
  assign mem[820] = 14'b10101001001110;
  assign mem[821] = 14'b01001110001011;
  assign mem[822] = 14'b00000000010001;
  assign mem[823] = 14'b00001000110101;
  assign mem[824] = 14'b01011100000011;
  assign mem[825] = 14'b10111110010001;
  assign mem[826] = 14'b10101100110010;
  assign mem[827] = 14'b10100010101100;
  assign mem[828] = 14'b10001010110101;
  assign mem[829] = 14'b00111110000110;
  assign mem[830] = 14'b10101011100101;
  assign mem[831] = 14'b01101111011010;
  assign mem[832] = 14'b01011011010000;
  assign mem[833] = 14'b10100011110010;
  assign mem[834] = 14'b10000010010010;
  assign mem[835] = 14'b01011110010011;
  assign mem[836] = 14'b01101100110100;
  assign mem[837] = 14'b00011000100110;
  assign mem[838] = 14'b10101010111000;
  assign mem[839] = 14'b00011111100100;
  assign mem[840] = 14'b00100110100001;
  assign mem[841] = 14'b01111111111111;
  assign mem[842] = 14'b00000110000000;
  assign mem[843] = 14'b00101001010010;
  assign mem[844] = 14'b00101010101001;
  assign mem[845] = 14'b01010100010111;
  assign mem[846] = 14'b00100001111111;
  assign mem[847] = 14'b10010010110100;
  assign mem[848] = 14'b10111011010011;
  assign mem[849] = 14'b01111101100011;
  assign mem[850] = 14'b01000100010111;
  assign mem[851] = 14'b01100111010011;
  assign mem[852] = 14'b01001110010010;
  assign mem[853] = 14'b10111000100100;
  assign mem[854] = 14'b10001110101011;
  assign mem[855] = 14'b10110010100011;
  assign mem[856] = 14'b00000001101000;
  assign mem[857] = 14'b01100011001100;
  assign mem[858] = 14'b10010110101011;
  assign mem[859] = 14'b01101001100101;
  assign mem[860] = 14'b10111101001110;
  assign mem[861] = 14'b01010111110001;
  assign mem[862] = 14'b10101010110111;
  assign mem[863] = 14'b00001000011101;
  assign mem[864] = 14'b00000010000111;
  assign mem[865] = 14'b00101111100001;
  assign mem[866] = 14'b01110000100000;
  assign mem[867] = 14'b01100101111110;
  assign mem[868] = 14'b01001111011101;
  assign mem[869] = 14'b10111101101000;
  assign mem[870] = 14'b00001101001010;
  assign mem[871] = 14'b01000000100001;
  assign mem[872] = 14'b01111000000101;
  assign mem[873] = 14'b10101101000111;
  assign mem[874] = 14'b10000011101010;
  assign mem[875] = 14'b00001111110000;
  assign mem[876] = 14'b00101010100101;
  assign mem[877] = 14'b10110111111100;
  assign mem[878] = 14'b01011110101010;
  assign mem[879] = 14'b00010001001101;
  assign mem[880] = 14'b00011110011110;
  assign mem[881] = 14'b10000011101000;
  assign mem[882] = 14'b01011000111000;
  assign mem[883] = 14'b01101011011100;
  assign mem[884] = 14'b10111011100101;
  assign mem[885] = 14'b10011101011111;
  assign mem[886] = 14'b01010011010111;
  assign mem[887] = 14'b00001110011111;
  assign mem[888] = 14'b00011011101010;
  assign mem[889] = 14'b00000100010001;
  assign mem[890] = 14'b10000010111001;
  assign mem[891] = 14'b00100011011111;
  assign mem[892] = 14'b01010001101001;
  assign mem[893] = 14'b10100000101011;
  assign mem[894] = 14'b00000001110100;
  assign mem[895] = 14'b10111000011111;
  assign mem[896] = 14'b00000001011011;
  assign mem[897] = 14'b10110110110011;
  assign mem[898] = 14'b00001011110101;
  assign mem[899] = 14'b00010100011000;
  assign mem[900] = 14'b01110101100100;
  assign mem[901] = 14'b01100100110011;
  assign mem[902] = 14'b01111101100000;
  assign mem[903] = 14'b01111111011010;
  assign mem[904] = 14'b01110100100000;
  assign mem[905] = 14'b01000001011111;
  assign mem[906] = 14'b00000100110101;
  assign mem[907] = 14'b00100100001110;
  assign mem[908] = 14'b00100011110100;
  assign mem[909] = 14'b10100010011001;
  assign mem[910] = 14'b10110101110111;
  assign mem[911] = 14'b10010100001001;
  assign mem[912] = 14'b10111111001110;
  assign mem[913] = 14'b10100101100010;
  assign mem[914] = 14'b10010101100001;
  assign mem[915] = 14'b01111011101000;
  assign mem[916] = 14'b10100010000000;
  assign mem[917] = 14'b10011010100001;
  assign mem[918] = 14'b10111111010100;
  assign mem[919] = 14'b01110000001011;
  assign mem[920] = 14'b00111101010100;
  assign mem[921] = 14'b00110001110100;
  assign mem[922] = 14'b00000101101111;
  assign mem[923] = 14'b00100000011101;
  assign mem[924] = 14'b00000101010000;
  assign mem[925] = 14'b01010100001000;
  assign mem[926] = 14'b01010111111111;
  assign mem[927] = 14'b10000110010100;
  assign mem[928] = 14'b01001000001101;
  assign mem[929] = 14'b00011011101111;
  assign mem[930] = 14'b10001010100010;
  assign mem[931] = 14'b00000111000011;
  assign mem[932] = 14'b01011111011100;
  assign mem[933] = 14'b00010100100101;
  assign mem[934] = 14'b01100001100110;
  assign mem[935] = 14'b10001001011011;
  assign mem[936] = 14'b01011100001000;
  assign mem[937] = 14'b01110001110011;
  assign mem[938] = 14'b00110000111100;
  assign mem[939] = 14'b10110100101100;
  assign mem[940] = 14'b01001101110001;
  assign mem[941] = 14'b10111110000001;
  assign mem[942] = 14'b01110011001011;
  assign mem[943] = 14'b00010101010110;
  assign mem[944] = 14'b10111101100010;
  assign mem[945] = 14'b10100101111011;
  assign mem[946] = 14'b00111011100001;
  assign mem[947] = 14'b01010000011101;
  assign mem[948] = 14'b01100010011100;
  assign mem[949] = 14'b00101001001110;
  assign mem[950] = 14'b01000001100101;
  assign mem[951] = 14'b00010110001010;
  assign mem[952] = 14'b10011101010001;
  assign mem[953] = 14'b01000000111100;
  assign mem[954] = 14'b10000010110101;
  assign mem[955] = 14'b10000111000100;
  assign mem[956] = 14'b10100011001101;
  assign mem[957] = 14'b00001101110010;
  assign mem[958] = 14'b01111111011110;
  assign mem[959] = 14'b10011110111101;
  assign mem[960] = 14'b10011000100011;
  assign mem[961] = 14'b10111110011111;
  assign mem[962] = 14'b00000111001011;
  assign mem[963] = 14'b00101110010110;
  assign mem[964] = 14'b00110001011110;
  assign mem[965] = 14'b00000110010101;
  assign mem[966] = 14'b01001110001000;
  assign mem[967] = 14'b10010001011111;
  assign mem[968] = 14'b01100100000100;
  assign mem[969] = 14'b10001100011010;
  assign mem[970] = 14'b00011000001111;
  assign mem[971] = 14'b01111111101111;
  assign mem[972] = 14'b00111000101110;
  assign mem[973] = 14'b10101000001110;
  assign mem[974] = 14'b10010000110001;
  assign mem[975] = 14'b00001010111100;
  assign mem[976] = 14'b10000101111101;
  assign mem[977] = 14'b10010100100100;
  assign mem[978] = 14'b01100111100110;
  assign mem[979] = 14'b10110010101101;
  assign mem[980] = 14'b10110101001011;
  assign mem[981] = 14'b01011011011010;
  assign mem[982] = 14'b00111101101110;
  assign mem[983] = 14'b01001010100111;
  assign mem[984] = 14'b10111010100101;
  assign mem[985] = 14'b00010110100110;
  assign mem[986] = 14'b01011110000010;
  assign mem[987] = 14'b00110100111010;
  assign mem[988] = 14'b10110011001110;
  assign mem[989] = 14'b01010010111110;
  assign mem[990] = 14'b01010101100100;
  assign mem[991] = 14'b00001000101001;
  assign mem[992] = 14'b10010100000010;
  assign mem[993] = 14'b00101000011010;
  assign mem[994] = 14'b00010110010111;
  assign mem[995] = 14'b00101010110101;
  assign mem[996] = 14'b00000111011001;
  assign mem[997] = 14'b10110001110111;
  assign mem[998] = 14'b01001010001001;
  assign mem[999] = 14'b00001101000100;
  assign mem[1000] = 14'b00111111011110;
  assign mem[1001] = 14'b10100110101010;
  assign mem[1002] = 14'b01111000101111;
  assign mem[1003] = 14'b10110111101000;
  assign mem[1004] = 14'b01010110011110;
  assign mem[1005] = 14'b00000100111000;
  assign mem[1006] = 14'b01000011010011;
  assign mem[1007] = 14'b01000011111111;
  assign mem[1008] = 14'b01011010000100;
  assign mem[1009] = 14'b10000111100111;
  assign mem[1010] = 14'b10000010111101;
  assign mem[1011] = 14'b01111111111011;
  assign mem[1012] = 14'b00000000000101;
  assign mem[1013] = 14'b01110011100011;
  assign mem[1014] = 14'b01000100001011;
  assign mem[1015] = 14'b00010010000000;
  assign mem[1016] = 14'b01010100101101;
  assign mem[1017] = 14'b01010001101111;
  assign mem[1018] = 14'b01100101001001;
  assign mem[1019] = 14'b00000110110100;
  assign mem[1020] = 14'b01110110001111;
  assign mem[1021] = 14'b10000110011011;
  assign mem[1022] = 14'b01100001010101;
  assign mem[1023] = 14'b10000000100110;

  always@(*)
  begin
    data_out_t <= mem[addr_f];
  end

  // Build output registers
  wire [13:0] data_out_reg [n_outreg:0];
  generate if (n_outreg > 0)
  begin
    for( i=n_outreg-1; i >= 1; i=i-1)
    begin: data_out_reg_stage
      mgc_generic_reg #(
        .width(14), 
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_data_out_reg (
        .d(data_out_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(data_out_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(14), 
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_data_out_reg_init (
      .d(data_out_t),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(data_out_reg[0])
    );
    assign data_out = data_out_reg[n_outreg-1];
  end
  else
  begin
    assign data_out = data_out_t;
  end
  endgenerate

endmodule



//------> ./rtl_stagemgc_rom_sync_regout_12_1024_14_1_0_0_1_0_1_0_0_0_1_60.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Sun Oct  6 01:48:34 2024
// ----------------------------------------------------------------------

// 
module stagemgc_rom_sync_regout_12_1024_14_1_0_0_1_0_1_0_0_0_1_60 (addr, data_out,
    clk, s_rst, a_rst, en
);
  input [9:0]addr ;
  output [13:0]data_out ;
  input clk ;
  input s_rst ;
  input a_rst ;
  input en ;


  // Constants for ROM dimensions
  parameter n_width    = 14;
  parameter n_size     = 1024;
  parameter n_numports = 1;
  parameter n_addr_w   = 10;
  parameter n_inreg    = 0;
  parameter n_outreg   = 1;
  wire [9:0] addr_f;

  // Build input address registers
  wire [9:0] addr_reg [n_inreg:0];
  genvar i;
  generate if (n_inreg > 0)
  begin
    for( i=n_inreg-1; i >= 1; i=i-1)
    begin: addr_reg_stage
      mgc_generic_reg #(
        .width(10), 
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_addr_reg (
        .d(addr_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(addr_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(10), 
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_addr_reg_init (
      .d(addr),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(addr_reg[0])
    );
    assign addr_f = addr_reg[n_inreg-1];
  end
  else
  begin
    assign addr_f = addr;
  end
  endgenerate

  // Declare storage for memory elements
  wire [13:0] mem [1023:0];

  // Declare output registers
  reg [13:0] data_out_t;

  // Initialize ROM contents
  assign mem[0] = 14'b00111111111011;
  assign mem[1] = 14'b01111011010000;
  assign mem[2] = 14'b10101100110100;
  assign mem[3] = 14'b10101111001000;
  assign mem[4] = 14'b01101100110000;
  assign mem[5] = 14'b01000011110110;
  assign mem[6] = 14'b01100010000011;
  assign mem[7] = 14'b10011000011111;
  assign mem[8] = 14'b00011000110111;
  assign mem[9] = 14'b01100011111111;
  assign mem[10] = 14'b10010100000101;
  assign mem[11] = 14'b01010010010010;
  assign mem[12] = 14'b00001001001010;
  assign mem[13] = 14'b01011011000001;
  assign mem[14] = 14'b01110101110010;
  assign mem[15] = 14'b10010111101110;
  assign mem[16] = 14'b00010001101110;
  assign mem[17] = 14'b01100100000111;
  assign mem[18] = 14'b00011010101111;
  assign mem[19] = 14'b00001111000101;
  assign mem[20] = 14'b01101110111011;
  assign mem[21] = 14'b01110111111010;
  assign mem[22] = 14'b00111010011111;
  assign mem[23] = 14'b01100100101010;
  assign mem[24] = 14'b10100010101110;
  assign mem[25] = 14'b01111110100100;
  assign mem[26] = 14'b00011101011101;
  assign mem[27] = 14'b00011010011000;
  assign mem[28] = 14'b00010101010100;
  assign mem[29] = 14'b10100001011001;
  assign mem[30] = 14'b10011110110100;
  assign mem[31] = 14'b10001111011100;
  assign mem[32] = 14'b10111110110010;
  assign mem[33] = 14'b01100001100000;
  assign mem[34] = 14'b00001111100101;
  assign mem[35] = 14'b00000001110101;
  assign mem[36] = 14'b01001010101111;
  assign mem[37] = 14'b01000100110111;
  assign mem[38] = 14'b00011000001101;
  assign mem[39] = 14'b01101110100000;
  assign mem[40] = 14'b00101100001101;
  assign mem[41] = 14'b01100100111010;
  assign mem[42] = 14'b01000101001111;
  assign mem[43] = 14'b10001010101101;
  assign mem[44] = 14'b01101111101000;
  assign mem[45] = 14'b00101000000100;
  assign mem[46] = 14'b01011000100000;
  assign mem[47] = 14'b00111111001010;
  assign mem[48] = 14'b10111110011101;
  assign mem[49] = 14'b00000110110000;
  assign mem[50] = 14'b10100111111111;
  assign mem[51] = 14'b00010011010101;
  assign mem[52] = 14'b01110110111010;
  assign mem[53] = 14'b00010111111110;
  assign mem[54] = 14'b00111110001111;
  assign mem[55] = 14'b01111010110111;
  assign mem[56] = 14'b00100010000101;
  assign mem[57] = 14'b01100010100100;
  assign mem[58] = 14'b10001000010000;
  assign mem[59] = 14'b01100110101010;
  assign mem[60] = 14'b01001011101011;
  assign mem[61] = 14'b00011010011010;
  assign mem[62] = 14'b00000000001110;
  assign mem[63] = 14'b00111100100000;
  assign mem[64] = 14'b01010111000001;
  assign mem[65] = 14'b10010010011000;
  assign mem[66] = 14'b10111110000011;
  assign mem[67] = 14'b00011111100011;
  assign mem[68] = 14'b01110101110111;
  assign mem[69] = 14'b00100100001011;
  assign mem[70] = 14'b01001001000001;
  assign mem[71] = 14'b01110010101100;
  assign mem[72] = 14'b00011000010001;
  assign mem[73] = 14'b00010010000100;
  assign mem[74] = 14'b10000011010001;
  assign mem[75] = 14'b10110001111101;
  assign mem[76] = 14'b00001111111100;
  assign mem[77] = 14'b00101110010111;
  assign mem[78] = 14'b10101000010100;
  assign mem[79] = 14'b01101110000101;
  assign mem[80] = 14'b00110011110100;
  assign mem[81] = 14'b10101111100100;
  assign mem[82] = 14'b01010010100101;
  assign mem[83] = 14'b10110100111010;
  assign mem[84] = 14'b10100110001101;
  assign mem[85] = 14'b10011101100110;
  assign mem[86] = 14'b10010100010101;
  assign mem[87] = 14'b01100000100100;
  assign mem[88] = 14'b10010000111101;
  assign mem[89] = 14'b01011111110010;
  assign mem[90] = 14'b00110011111011;
  assign mem[91] = 14'b00001101110011;
  assign mem[92] = 14'b10100011100101;
  assign mem[93] = 14'b00000111101001;
  assign mem[94] = 14'b00010111011110;
  assign mem[95] = 14'b00101100100011;
  assign mem[96] = 14'b10101100110101;
  assign mem[97] = 14'b10011000000001;
  assign mem[98] = 14'b00101010110110;
  assign mem[99] = 14'b10111111010001;
  assign mem[100] = 14'b01001101101010;
  assign mem[101] = 14'b10100011110001;
  assign mem[102] = 14'b10011101011110;
  assign mem[103] = 14'b00010010101011;
  assign mem[104] = 14'b00001011011010;
  assign mem[105] = 14'b00011011100010;
  assign mem[106] = 14'b00111100001110;
  assign mem[107] = 14'b00011111101110;
  assign mem[108] = 14'b01011100000100;
  assign mem[109] = 14'b10101010101010;
  assign mem[110] = 14'b10001100111100;
  assign mem[111] = 14'b01010010011010;
  assign mem[112] = 14'b10001111011011;
  assign mem[113] = 14'b00111000010100;
  assign mem[114] = 14'b00111011000110;
  assign mem[115] = 14'b10011111011110;
  assign mem[116] = 14'b00110001101100;
  assign mem[117] = 14'b00110110001011;
  assign mem[118] = 14'b01001000111100;
  assign mem[119] = 14'b00100110001110;
  assign mem[120] = 14'b01110110111101;
  assign mem[121] = 14'b10010010101010;
  assign mem[122] = 14'b00001101000010;
  assign mem[123] = 14'b01111000010111;
  assign mem[124] = 14'b01101010110100;
  assign mem[125] = 14'b00110101001011;
  assign mem[126] = 14'b01010011100111;
  assign mem[127] = 14'b10111111110100;
  assign mem[128] = 14'b00110111111100;
  assign mem[129] = 14'b00011011001011;
  assign mem[130] = 14'b10101001000100;
  assign mem[131] = 14'b10011000111011;
  assign mem[132] = 14'b10011111100001;
  assign mem[133] = 14'b00111111100110;
  assign mem[134] = 14'b10111111011010;
  assign mem[135] = 14'b10000101001101;
  assign mem[136] = 14'b10100010100001;
  assign mem[137] = 14'b00101010111101;
  assign mem[138] = 14'b01110010101010;
  assign mem[139] = 14'b10100101001110;
  assign mem[140] = 14'b01011110011000;
  assign mem[141] = 14'b00001110101111;
  assign mem[142] = 14'b10010001110010;
  assign mem[143] = 14'b00010111000101;
  assign mem[144] = 14'b01101011010001;
  assign mem[145] = 14'b10010111000100;
  assign mem[146] = 14'b00111000000001;
  assign mem[147] = 14'b01100111101001;
  assign mem[148] = 14'b10111101110001;
  assign mem[149] = 14'b00111111011111;
  assign mem[150] = 14'b00111001100100;
  assign mem[151] = 14'b01111000000000;
  assign mem[152] = 14'b01111111111100;
  assign mem[153] = 14'b01101011110110;
  assign mem[154] = 14'b00110111001101;
  assign mem[155] = 14'b10011001001111;
  assign mem[156] = 14'b01011111001010;
  assign mem[157] = 14'b00001011010111;
  assign mem[158] = 14'b10011101110011;
  assign mem[159] = 14'b01101101011011;
  assign mem[160] = 14'b01101100100001;
  assign mem[161] = 14'b00011110011101;
  assign mem[162] = 14'b10011000000011;
  assign mem[163] = 14'b10100100111111;
  assign mem[164] = 14'b01011110101001;
  assign mem[165] = 14'b00000101111010;
  assign mem[166] = 14'b01111010111111;
  assign mem[167] = 14'b10001000111011;
  assign mem[168] = 14'b10001011000101;
  assign mem[169] = 14'b10010000001101;
  assign mem[170] = 14'b10001010001110;
  assign mem[171] = 14'b01000111000111;
  assign mem[172] = 14'b10010101110101;
  assign mem[173] = 14'b10110110010000;
  assign mem[174] = 14'b01110111001110;
  assign mem[175] = 14'b10001001110101;
  assign mem[176] = 14'b01011000110000;
  assign mem[177] = 14'b01001101011100;
  assign mem[178] = 14'b01100001101011;
  assign mem[179] = 14'b10000011000100;
  assign mem[180] = 14'b10011110101100;
  assign mem[181] = 14'b10001000010011;
  assign mem[182] = 14'b00100100100101;
  assign mem[183] = 14'b00110001010111;
  assign mem[184] = 14'b00010110111011;
  assign mem[185] = 14'b01010101010100;
  assign mem[186] = 14'b10000101101001;
  assign mem[187] = 14'b01111001100111;
  assign mem[188] = 14'b00101001011001;
  assign mem[189] = 14'b00100100010000;
  assign mem[190] = 14'b10001101001100;
  assign mem[191] = 14'b01100000101100;
  assign mem[192] = 14'b00001011100001;
  assign mem[193] = 14'b00111001110010;
  assign mem[194] = 14'b01001001011011;
  assign mem[195] = 14'b01011001111001;
  assign mem[196] = 14'b10001101010110;
  assign mem[197] = 14'b00111001100111;
  assign mem[198] = 14'b00000000010000;
  assign mem[199] = 14'b00001110010010;
  assign mem[200] = 14'b01010001000010;
  assign mem[201] = 14'b10100100100011;
  assign mem[202] = 14'b01000111001000;
  assign mem[203] = 14'b00011110101100;
  assign mem[204] = 14'b00110110110101;
  assign mem[205] = 14'b10000011110100;
  assign mem[206] = 14'b01110101011100;
  assign mem[207] = 14'b01010100000101;
  assign mem[208] = 14'b10100111101101;
  assign mem[209] = 14'b00110011010001;
  assign mem[210] = 14'b01101101111101;
  assign mem[211] = 14'b00010000100100;
  assign mem[212] = 14'b00101101001111;
  assign mem[213] = 14'b01101111110100;
  assign mem[214] = 14'b10001010110111;
  assign mem[215] = 14'b01010011101101;
  assign mem[216] = 14'b01100100001001;
  assign mem[217] = 14'b10000000000101;
  assign mem[218] = 14'b00101110010010;
  assign mem[219] = 14'b01100011100111;
  assign mem[220] = 14'b01001111001000;
  assign mem[221] = 14'b01100111101010;
  assign mem[222] = 14'b01010111111001;
  assign mem[223] = 14'b00000100010110;
  assign mem[224] = 14'b00001110100100;
  assign mem[225] = 14'b10011111110101;
  assign mem[226] = 14'b10001011011111;
  assign mem[227] = 14'b01110111011010;
  assign mem[228] = 14'b00000101011111;
  assign mem[229] = 14'b10010001010010;
  assign mem[230] = 14'b00000011101101;
  assign mem[231] = 14'b01011011100010;
  assign mem[232] = 14'b01111000001100;
  assign mem[233] = 14'b00110001001010;
  assign mem[234] = 14'b10111101011110;
  assign mem[235] = 14'b01110110100010;
  assign mem[236] = 14'b00100000000101;
  assign mem[237] = 14'b10110000010101;
  assign mem[238] = 14'b00111011011010;
  assign mem[239] = 14'b01010001010100;
  assign mem[240] = 14'b01000111111010;
  assign mem[241] = 14'b00011011010100;
  assign mem[242] = 14'b10110000100100;
  assign mem[243] = 14'b00000101010100;
  assign mem[244] = 14'b00111001111111;
  assign mem[245] = 14'b01001000000110;
  assign mem[246] = 14'b00000100101100;
  assign mem[247] = 14'b10101011110001;
  assign mem[248] = 14'b01001111001110;
  assign mem[249] = 14'b10011101000001;
  assign mem[250] = 14'b10110101100000;
  assign mem[251] = 14'b10111111010111;
  assign mem[252] = 14'b01110011111101;
  assign mem[253] = 14'b10100111010011;
  assign mem[254] = 14'b01011001110010;
  assign mem[255] = 14'b01011000010110;
  assign mem[256] = 14'b00111011111011;
  assign mem[257] = 14'b01010110110001;
  assign mem[258] = 14'b00010011001000;
  assign mem[259] = 14'b10000100011100;
  assign mem[260] = 14'b10010000010101;
  assign mem[261] = 14'b00111100000101;
  assign mem[262] = 14'b00000011111010;
  assign mem[263] = 14'b10101111001001;
  assign mem[264] = 14'b01000010000001;
  assign mem[265] = 14'b01100010110110;
  assign mem[266] = 14'b10010111010000;
  assign mem[267] = 14'b10111111011110;
  assign mem[268] = 14'b01000000101000;
  assign mem[269] = 14'b00101011011010;
  assign mem[270] = 14'b00001010110100;
  assign mem[271] = 14'b10001001101000;
  assign mem[272] = 14'b01100100001010;
  assign mem[273] = 14'b01101000111110;
  assign mem[274] = 14'b10011101111001;
  assign mem[275] = 14'b10100010110010;
  assign mem[276] = 14'b00111010101111;
  assign mem[277] = 14'b01110010111100;
  assign mem[278] = 14'b10110001100001;
  assign mem[279] = 14'b10000011110001;
  assign mem[280] = 14'b01100100100101;
  assign mem[281] = 14'b00111001000100;
  assign mem[282] = 14'b01100011000110;
  assign mem[283] = 14'b10001100010010;
  assign mem[284] = 14'b01010100001111;
  assign mem[285] = 14'b00100011100000;
  assign mem[286] = 14'b01100101001100;
  assign mem[287] = 14'b01110011111000;
  assign mem[288] = 14'b10000011100010;
  assign mem[289] = 14'b10101001001000;
  assign mem[290] = 14'b10111011010010;
  assign mem[291] = 14'b01011001100101;
  assign mem[292] = 14'b00001101101100;
  assign mem[293] = 14'b01101101110110;
  assign mem[294] = 14'b00100001110111;
  assign mem[295] = 14'b00100110000100;
  assign mem[296] = 14'b00110101110010;
  assign mem[297] = 14'b10010000000001;
  assign mem[298] = 14'b10000000001110;
  assign mem[299] = 14'b01001011111010;
  assign mem[300] = 14'b01011101001100;
  assign mem[301] = 14'b00101010111010;
  assign mem[302] = 14'b01110000001010;
  assign mem[303] = 14'b00010110011010;
  assign mem[304] = 14'b01110011011101;
  assign mem[305] = 14'b10001010101111;
  assign mem[306] = 14'b10100110100101;
  assign mem[307] = 14'b10110011000001;
  assign mem[308] = 14'b01000001111100;
  assign mem[309] = 14'b00010110011000;
  assign mem[310] = 14'b10101001010000;
  assign mem[311] = 14'b01000011101000;
  assign mem[312] = 14'b10000101101101;
  assign mem[313] = 14'b00011101001011;
  assign mem[314] = 14'b10010011101110;
  assign mem[315] = 14'b00100101110000;
  assign mem[316] = 14'b00111011101000;
  assign mem[317] = 14'b10001101110100;
  assign mem[318] = 14'b00001010101110;
  assign mem[319] = 14'b01010100010001;
  assign mem[320] = 14'b00100111011011;
  assign mem[321] = 14'b01000011110011;
  assign mem[322] = 14'b01011111100011;
  assign mem[323] = 14'b00001001101011;
  assign mem[324] = 14'b00001110101001;
  assign mem[325] = 14'b00101100010010;
  assign mem[326] = 14'b01111001011111;
  assign mem[327] = 14'b00110011001111;
  assign mem[328] = 14'b00100100111011;
  assign mem[329] = 14'b01110101000000;
  assign mem[330] = 14'b01011111100000;
  assign mem[331] = 14'b01001111000000;
  assign mem[332] = 14'b00001100111000;
  assign mem[333] = 14'b10011111011100;
  assign mem[334] = 14'b10110110101010;
  assign mem[335] = 14'b00010001011001;
  assign mem[336] = 14'b00101010100111;
  assign mem[337] = 14'b10011001111000;
  assign mem[338] = 14'b00001110000000;
  assign mem[339] = 14'b00011111101100;
  assign mem[340] = 14'b01001111010011;
  assign mem[341] = 14'b00101001011110;
  assign mem[342] = 14'b10100011100000;
  assign mem[343] = 14'b01111011001100;
  assign mem[344] = 14'b10111110001001;
  assign mem[345] = 14'b01010100111010;
  assign mem[346] = 14'b00101111111110;
  assign mem[347] = 14'b01100100000000;
  assign mem[348] = 14'b10001110101100;
  assign mem[349] = 14'b10110110011000;
  assign mem[350] = 14'b10111101111001;
  assign mem[351] = 14'b01000110101000;
  assign mem[352] = 14'b00010011111001;
  assign mem[353] = 14'b10011000001011;
  assign mem[354] = 14'b10110011001100;
  assign mem[355] = 14'b10011011010001;
  assign mem[356] = 14'b10011100110111;
  assign mem[357] = 14'b10010111111000;
  assign mem[358] = 14'b00100011010110;
  assign mem[359] = 14'b10010010110111;
  assign mem[360] = 14'b10101110111000;
  assign mem[361] = 14'b00000100111011;
  assign mem[362] = 14'b01000110011111;
  assign mem[363] = 14'b00010010000110;
  assign mem[364] = 14'b01011110101101;
  assign mem[365] = 14'b01101001011111;
  assign mem[366] = 14'b10111001011001;
  assign mem[367] = 14'b00000101100101;
  assign mem[368] = 14'b01110011000111;
  assign mem[369] = 14'b01000111000110;
  assign mem[370] = 14'b00001111010111;
  assign mem[371] = 14'b10000101010110;
  assign mem[372] = 14'b10000010100000;
  assign mem[373] = 14'b10011110001110;
  assign mem[374] = 14'b01110101101010;
  assign mem[375] = 14'b10010000100101;
  assign mem[376] = 14'b01000100001111;
  assign mem[377] = 14'b01010001100101;
  assign mem[378] = 14'b00111110011111;
  assign mem[379] = 14'b10001001001001;
  assign mem[380] = 14'b00110001011001;
  assign mem[381] = 14'b01101101001110;
  assign mem[382] = 14'b01000000100010;
  assign mem[383] = 14'b10110110000100;
  assign mem[384] = 14'b00110100101110;
  assign mem[385] = 14'b10110011010101;
  assign mem[386] = 14'b00011011011001;
  assign mem[387] = 14'b00000100100100;
  assign mem[388] = 14'b10000111101001;
  assign mem[389] = 14'b00101011110110;
  assign mem[390] = 14'b10100010001010;
  assign mem[391] = 14'b10111110011100;
  assign mem[392] = 14'b01011010101000;
  assign mem[393] = 14'b10111000100011;
  assign mem[394] = 14'b00110001101101;
  assign mem[395] = 14'b00011111000100;
  assign mem[396] = 14'b00010000000000;
  assign mem[397] = 14'b10010001111100;
  assign mem[398] = 14'b00100110101101;
  assign mem[399] = 14'b10101010110000;
  assign mem[400] = 14'b01000111100110;
  assign mem[401] = 14'b01101001011110;
  assign mem[402] = 14'b00111000100011;
  assign mem[403] = 14'b01010101111111;
  assign mem[404] = 14'b01010001110001;
  assign mem[405] = 14'b00100110011111;
  assign mem[406] = 14'b10000100010110;
  assign mem[407] = 14'b01110111100010;
  assign mem[408] = 14'b01111100011100;
  assign mem[409] = 14'b01100011111011;
  assign mem[410] = 14'b00010000101111;
  assign mem[411] = 14'b00010011111000;
  assign mem[412] = 14'b00110110010010;
  assign mem[413] = 14'b10101100100101;
  assign mem[414] = 14'b00110011011011;
  assign mem[415] = 14'b10110001010000;
  assign mem[416] = 14'b10000100110110;
  assign mem[417] = 14'b10010100000110;
  assign mem[418] = 14'b10011001101101;
  assign mem[419] = 14'b00010011100101;
  assign mem[420] = 14'b00011101000001;
  assign mem[421] = 14'b01100001011001;
  assign mem[422] = 14'b01001001110000;
  assign mem[423] = 14'b10110100101001;
  assign mem[424] = 14'b01011110010010;
  assign mem[425] = 14'b10011001011001;
  assign mem[426] = 14'b00110100001011;
  assign mem[427] = 14'b00011100000101;
  assign mem[428] = 14'b00101100111111;
  assign mem[429] = 14'b01100001100010;
  assign mem[430] = 14'b01010001010000;
  assign mem[431] = 14'b00100001000010;
  assign mem[432] = 14'b01111100011010;
  assign mem[433] = 14'b10010010001001;
  assign mem[434] = 14'b10110001100011;
  assign mem[435] = 14'b01010101100011;
  assign mem[436] = 14'b01011111000100;
  assign mem[437] = 14'b10010110000001;
  assign mem[438] = 14'b01000000001100;
  assign mem[439] = 14'b01110010011011;
  assign mem[440] = 14'b10100011000110;
  assign mem[441] = 14'b10010011111111;
  assign mem[442] = 14'b00010011110111;
  assign mem[443] = 14'b00000110011000;
  assign mem[444] = 14'b01101011111111;
  assign mem[445] = 14'b00110000000111;
  assign mem[446] = 14'b00000101101000;
  assign mem[447] = 14'b10000001010100;
  assign mem[448] = 14'b10110100001111;
  assign mem[449] = 14'b10001111000100;
  assign mem[450] = 14'b10001101011001;
  assign mem[451] = 14'b10110100010011;
  assign mem[452] = 14'b00001101010010;
  assign mem[453] = 14'b10000110101001;
  assign mem[454] = 14'b00001100010000;
  assign mem[455] = 14'b01111011101111;
  assign mem[456] = 14'b10000010001110;
  assign mem[457] = 14'b10111110001010;
  assign mem[458] = 14'b00011100110110;
  assign mem[459] = 14'b10011111100101;
  assign mem[460] = 14'b10111110011000;
  assign mem[461] = 14'b01111010010011;
  assign mem[462] = 14'b10111001111111;
  assign mem[463] = 14'b01010111100000;
  assign mem[464] = 14'b10011000110011;
  assign mem[465] = 14'b00001111110100;
  assign mem[466] = 14'b00001011010001;
  assign mem[467] = 14'b00101011100000;
  assign mem[468] = 14'b01101000010100;
  assign mem[469] = 14'b01100110011000;
  assign mem[470] = 14'b01010011100100;
  assign mem[471] = 14'b01000101001000;
  assign mem[472] = 14'b01101010100000;
  assign mem[473] = 14'b10000011010101;
  assign mem[474] = 14'b10011011100111;
  assign mem[475] = 14'b01010000011110;
  assign mem[476] = 14'b00100100110100;
  assign mem[477] = 14'b01010110110000;
  assign mem[478] = 14'b01010010010011;
  assign mem[479] = 14'b00010100110101;
  assign mem[480] = 14'b10001001100001;
  assign mem[481] = 14'b10010110111101;
  assign mem[482] = 14'b01110010001100;
  assign mem[483] = 14'b01011010011100;
  assign mem[484] = 14'b01001100101110;
  assign mem[485] = 14'b00001110001101;
  assign mem[486] = 14'b10110101011101;
  assign mem[487] = 14'b01000100101011;
  assign mem[488] = 14'b10000000101110;
  assign mem[489] = 14'b01101000011110;
  assign mem[490] = 14'b01000011001110;
  assign mem[491] = 14'b00101111100100;
  assign mem[492] = 14'b00100011101101;
  assign mem[493] = 14'b10111111011001;
  assign mem[494] = 14'b00011110101011;
  assign mem[495] = 14'b10010000000000;
  assign mem[496] = 14'b01000011001000;
  assign mem[497] = 14'b10111010001110;
  assign mem[498] = 14'b00001010110111;
  assign mem[499] = 14'b01000100010011;
  assign mem[500] = 14'b10011001000001;
  assign mem[501] = 14'b01001100010100;
  assign mem[502] = 14'b00100101101011;
  assign mem[503] = 14'b10011111110110;
  assign mem[504] = 14'b00101001011010;
  assign mem[505] = 14'b00001101001001;
  assign mem[506] = 14'b00111100110010;
  assign mem[507] = 14'b10011111110111;
  assign mem[508] = 14'b01110001010000;
  assign mem[509] = 14'b10000100111001;
  assign mem[510] = 14'b10101110111100;
  assign mem[511] = 14'b01101000100000;
  assign mem[512] = 14'b00111111011011;
  assign mem[513] = 14'b01011110101100;
  assign mem[514] = 14'b00111001100110;
  assign mem[515] = 14'b01001001110010;
  assign mem[516] = 14'b10111001001101;
  assign mem[517] = 14'b01011010111000;
  assign mem[518] = 14'b01101110010010;
  assign mem[519] = 14'b01101011010100;
  assign mem[520] = 14'b10101110000001;
  assign mem[521] = 14'b01111011110110;
  assign mem[522] = 14'b01001100011110;
  assign mem[523] = 14'b10111111111100;
  assign mem[524] = 14'b01000000000110;
  assign mem[525] = 14'b00111101000100;
  assign mem[526] = 14'b00111000011010;
  assign mem[527] = 14'b01100101111101;
  assign mem[528] = 14'b01111100000010;
  assign mem[529] = 14'b01111100101110;
  assign mem[530] = 14'b10111011001001;
  assign mem[531] = 14'b01101001100011;
  assign mem[532] = 14'b00001000011001;
  assign mem[533] = 14'b01000111010010;
  assign mem[534] = 14'b00011001010111;
  assign mem[535] = 14'b10000000100011;
  assign mem[536] = 14'b10110010111101;
  assign mem[537] = 14'b01110101111000;
  assign mem[538] = 14'b00001110001010;
  assign mem[539] = 14'b10111000101000;
  assign mem[540] = 14'b10010101001100;
  assign mem[541] = 14'b10101001101010;
  assign mem[542] = 14'b10010111100111;
  assign mem[543] = 14'b00101011111111;
  assign mem[544] = 14'b10110111011000;
  assign mem[545] = 14'b01101010011101;
  assign mem[546] = 14'b01101101000011;
  assign mem[547] = 14'b00001100110011;
  assign mem[548] = 14'b10001011000111;
  assign mem[549] = 14'b01100001111111;
  assign mem[550] = 14'b10101001011011;
  assign mem[551] = 14'b00000101011100;
  assign mem[552] = 14'b01110101011010;
  assign mem[553] = 14'b10000010010011;
  assign mem[554] = 14'b01100100100111;
  assign mem[555] = 14'b00001010110110;
  assign mem[556] = 14'b00001101010100;
  assign mem[557] = 14'b01011000011011;
  assign mem[558] = 14'b00101011011101;
  assign mem[559] = 14'b00111010000100;
  assign mem[560] = 14'b10110101000101;
  assign mem[561] = 14'b00101111010000;
  assign mem[562] = 14'b00010111110011;
  assign mem[563] = 14'b10000111010011;
  assign mem[564] = 14'b01000000010010;
  assign mem[565] = 14'b10100111110010;
  assign mem[566] = 14'b00110011100111;
  assign mem[567] = 14'b01011011111101;
  assign mem[568] = 14'b00101110100010;
  assign mem[569] = 14'b01110001111001;
  assign mem[570] = 14'b10111001101100;
  assign mem[571] = 14'b10001110100011;
  assign mem[572] = 14'b10010001101011;
  assign mem[573] = 14'b10111000110110;
  assign mem[574] = 14'b00000001100010;
  assign mem[575] = 14'b00100111011110;
  assign mem[576] = 14'b00100001000100;
  assign mem[577] = 14'b01000000100011;
  assign mem[578] = 14'b10110010001111;
  assign mem[579] = 14'b00011100110100;
  assign mem[580] = 14'b00111000111101;
  assign mem[581] = 14'b00111101001100;
  assign mem[582] = 14'b01111111000101;
  assign mem[583] = 14'b00100010110000;
  assign mem[584] = 14'b10101001110111;
  assign mem[585] = 14'b01111110011100;
  assign mem[586] = 14'b10010110110011;
  assign mem[587] = 14'b01011101100101;
  assign mem[588] = 14'b01101111100100;
  assign mem[589] = 14'b10000100100000;
  assign mem[590] = 14'b00011010000110;
  assign mem[591] = 14'b00000010011111;
  assign mem[592] = 14'b10101010101011;
  assign mem[593] = 14'b01001100110110;
  assign mem[594] = 14'b00000010000000;
  assign mem[595] = 14'b01110010010000;
  assign mem[596] = 14'b00001011010101;
  assign mem[597] = 14'b10001111000101;
  assign mem[598] = 14'b01001110001110;
  assign mem[599] = 14'b01100011111001;
  assign mem[600] = 14'b00110110100110;
  assign mem[601] = 14'b01011110011011;
  assign mem[602] = 14'b10101011011100;
  assign mem[603] = 14'b01100000100101;
  assign mem[604] = 14'b10111000111110;
  assign mem[605] = 14'b00110101011111;
  assign mem[606] = 14'b10100100010010;
  assign mem[607] = 14'b01110111110100;
  assign mem[608] = 14'b00111001101101;
  assign mem[609] = 14'b01101000000010;
  assign mem[610] = 14'b01101011111001;
  assign mem[611] = 14'b10111010110001;
  assign mem[612] = 14'b10011111100100;
  assign mem[613] = 14'b10111010010010;
  assign mem[614] = 14'b10001110001101;
  assign mem[615] = 14'b10000010101101;
  assign mem[616] = 14'b01001111110110;
  assign mem[617] = 14'b00000000101101;
  assign mem[618] = 14'b00100101100000;
  assign mem[619] = 14'b00011110000001;
  assign mem[620] = 14'b01000100011001;
  assign mem[621] = 14'b00101010100000;
  assign mem[622] = 14'b00011010011111;
  assign mem[623] = 14'b00000000110011;
  assign mem[624] = 14'b00101011111000;
  assign mem[625] = 14'b00001010001010;
  assign mem[626] = 14'b00011101101000;
  assign mem[627] = 14'b10011100001101;
  assign mem[628] = 14'b10011011110011;
  assign mem[629] = 14'b10111011001100;
  assign mem[630] = 14'b01111110100010;
  assign mem[631] = 14'b01001011100001;
  assign mem[632] = 14'b01000000100111;
  assign mem[633] = 14'b01000010100001;
  assign mem[634] = 14'b01011011001110;
  assign mem[635] = 14'b01001010011101;
  assign mem[636] = 14'b10101011101001;
  assign mem[637] = 14'b10110100001100;
  assign mem[638] = 14'b00001001001110;
  assign mem[639] = 14'b10111110100110;
  assign mem[640] = 14'b00000111100010;
  assign mem[641] = 14'b10111110001101;
  assign mem[642] = 14'b00011111010110;
  assign mem[643] = 14'b01101110011000;
  assign mem[644] = 14'b10011100100010;
  assign mem[645] = 14'b00111101001000;
  assign mem[646] = 14'b10111011110000;
  assign mem[647] = 14'b10100100010111;
  assign mem[648] = 14'b10110001100010;
  assign mem[649] = 14'b01101100101010;
  assign mem[650] = 14'b00100010100010;
  assign mem[651] = 14'b00000100011100;
  assign mem[652] = 14'b01010100100101;
  assign mem[653] = 14'b01100111001001;
  assign mem[654] = 14'b00111100011001;
  assign mem[655] = 14'b10100001100011;
  assign mem[656] = 14'b10101110110100;
  assign mem[657] = 14'b01100001010111;
  assign mem[658] = 14'b00001000000101;
  assign mem[659] = 14'b10010101011100;
  assign mem[660] = 14'b10110000010001;
  assign mem[661] = 14'b00111100010111;
  assign mem[662] = 14'b00010010111010;
  assign mem[663] = 14'b01000111111100;
  assign mem[664] = 14'b01111111100000;
  assign mem[665] = 14'b10110010110111;
  assign mem[666] = 14'b00000010011001;
  assign mem[667] = 14'b01110000100100;
  assign mem[668] = 14'b01011010000011;
  assign mem[669] = 14'b01001111100001;
  assign mem[670] = 14'b10010000100000;
  assign mem[671] = 14'b10111101111010;
  assign mem[672] = 14'b10110111100100;
  assign mem[673] = 14'b00010101001010;
  assign mem[674] = 14'b01101000010000;
  assign mem[675] = 14'b00000010110011;
  assign mem[676] = 14'b01010110011100;
  assign mem[677] = 14'b00101001010110;
  assign mem[678] = 14'b01011100110101;
  assign mem[679] = 14'b10111110011001;
  assign mem[680] = 14'b00001101011110;
  assign mem[681] = 14'b00110001010110;
  assign mem[682] = 14'b00000111011101;
  assign mem[683] = 14'b01110001101111;
  assign mem[684] = 14'b01011000101110;
  assign mem[685] = 14'b01111011101010;
  assign mem[686] = 14'b01000010011110;
  assign mem[687] = 14'b00000100101110;
  assign mem[688] = 14'b00101101001101;
  assign mem[689] = 14'b10011110000010;
  assign mem[690] = 14'b01101011101010;
  assign mem[691] = 14'b10010101011000;
  assign mem[692] = 14'b10010110101111;
  assign mem[693] = 14'b10111010000001;
  assign mem[694] = 14'b01000000000010;
  assign mem[695] = 14'b10011001100000;
  assign mem[696] = 14'b10100000011101;
  assign mem[697] = 14'b00010101001001;
  assign mem[698] = 14'b10100111011011;
  assign mem[699] = 14'b01010011001101;
  assign mem[700] = 14'b01100001101110;
  assign mem[701] = 14'b00111101101111;
  assign mem[702] = 14'b00011100001111;
  assign mem[703] = 14'b01100100110001;
  assign mem[704] = 14'b01010000100111;
  assign mem[705] = 14'b00010100011100;
  assign mem[706] = 14'b10000001111011;
  assign mem[707] = 14'b00110101001100;
  assign mem[708] = 14'b00011101010101;
  assign mem[709] = 14'b00010011001111;
  assign mem[710] = 14'b00000001110000;
  assign mem[711] = 14'b01100011111110;
  assign mem[712] = 14'b10110111001100;
  assign mem[713] = 14'b10111111110000;
  assign mem[714] = 14'b01110001110110;
  assign mem[715] = 14'b00010110110011;
  assign mem[716] = 14'b10111111110010;
  assign mem[717] = 14'b10011010101000;
  assign mem[718] = 14'b00110110000000;
  assign mem[719] = 14'b00001100100000;
  assign mem[720] = 14'b00010101110101;
  assign mem[721] = 14'b10100110110110;
  assign mem[722] = 14'b00000001100111;
  assign mem[723] = 14'b01110011111100;
  assign mem[724] = 14'b01111100101000;
  assign mem[725] = 14'b00001110101000;
  assign mem[726] = 14'b00001011111100;
  assign mem[727] = 14'b00001001111000;
  assign mem[728] = 14'b01111100111100;
  assign mem[729] = 14'b10000000011111;
  assign mem[730] = 14'b10000011111101;
  assign mem[731] = 14'b01111001001110;
  assign mem[732] = 14'b10101001110110;
  assign mem[733] = 14'b10010101100011;
  assign mem[734] = 14'b00100111001100;
  assign mem[735] = 14'b00011110011010;
  assign mem[736] = 14'b01100101111100;
  assign mem[737] = 14'b10011110101110;
  assign mem[738] = 14'b00010000010100;
  assign mem[739] = 14'b01000011110010;
  assign mem[740] = 14'b00100110011001;
  assign mem[741] = 14'b00111000111001;
  assign mem[742] = 14'b00011001111011;
  assign mem[743] = 14'b01000000101011;
  assign mem[744] = 14'b01001001010000;
  assign mem[745] = 14'b10011000000101;
  assign mem[746] = 14'b10101110001100;
  assign mem[747] = 14'b00111101101010;
  assign mem[748] = 14'b00100000100010;
  assign mem[749] = 14'b01010010001101;
  assign mem[750] = 14'b00011111110100;
  assign mem[751] = 14'b10111001001010;
  assign mem[752] = 14'b01110111010100;
  assign mem[753] = 14'b10111111001100;
  assign mem[754] = 14'b01010011110110;
  assign mem[755] = 14'b00100101001100;
  assign mem[756] = 14'b00010101110111;
  assign mem[757] = 14'b01111000101000;
  assign mem[758] = 14'b00100000110100;
  assign mem[759] = 14'b00110010010001;
  assign mem[760] = 14'b10101010100000;
  assign mem[761] = 14'b10001011000010;
  assign mem[762] = 14'b01110110011010;
  assign mem[763] = 14'b10111011011011;
  assign mem[764] = 14'b00101011100111;
  assign mem[765] = 14'b00010010111111;
  assign mem[766] = 14'b00110100011011;
  assign mem[767] = 14'b00101010010111;
  assign mem[768] = 14'b00100011011011;
  assign mem[769] = 14'b00011111010100;
  assign mem[770] = 14'b10000101111000;
  assign mem[771] = 14'b10011111000000;
  assign mem[772] = 14'b00110010001110;
  assign mem[773] = 14'b00100100100001;
  assign mem[774] = 14'b00011011010110;
  assign mem[775] = 14'b01001001111001;
  assign mem[776] = 14'b01001110000101;
  assign mem[777] = 14'b01110011110111;
  assign mem[778] = 14'b01100010101011;
  assign mem[779] = 14'b10111100001100;
  assign mem[780] = 14'b01000100010110;
  assign mem[781] = 14'b01101111110101;
  assign mem[782] = 14'b01001011101100;
  assign mem[783] = 14'b00000011010011;
  assign mem[784] = 14'b01111101000011;
  assign mem[785] = 14'b10011110101111;
  assign mem[786] = 14'b10010001001010;
  assign mem[787] = 14'b10110011011001;
  assign mem[788] = 14'b00011011000111;
  assign mem[789] = 14'b00100100100000;
  assign mem[790] = 14'b01011010100001;
  assign mem[791] = 14'b10011010010011;
  assign mem[792] = 14'b10000000000000;
  assign mem[793] = 14'b00001111011010;
  assign mem[794] = 14'b01110101100111;
  assign mem[795] = 14'b00010101111001;
  assign mem[796] = 14'b00001101100110;
  assign mem[797] = 14'b00111000011111;
  assign mem[798] = 14'b10000100010001;
  assign mem[799] = 14'b00101011000100;
  assign mem[800] = 14'b10011000101010;
  assign mem[801] = 14'b00011111110010;
  assign mem[802] = 14'b10011110111000;
  assign mem[803] = 14'b00110011000000;
  assign mem[804] = 14'b01011111110100;
  assign mem[805] = 14'b00000000110110;
  assign mem[806] = 14'b00101101000000;
  assign mem[807] = 14'b01001010011011;
  assign mem[808] = 14'b10111000011101;
  assign mem[809] = 14'b00110000000010;
  assign mem[810] = 14'b10000001011110;
  assign mem[811] = 14'b10010011010100;
  assign mem[812] = 14'b01001100010001;
  assign mem[813] = 14'b01101100010101;
  assign mem[814] = 14'b00010001000010;
  assign mem[815] = 14'b10011100110110;
  assign mem[816] = 14'b00101000000111;
  assign mem[817] = 14'b00001011000100;
  assign mem[818] = 14'b00001101111101;
  assign mem[819] = 14'b01100101000001;
  assign mem[820] = 14'b01001101100010;
  assign mem[821] = 14'b10011100101000;
  assign mem[822] = 14'b00100000101010;
  assign mem[823] = 14'b01011001010110;
  assign mem[824] = 14'b10100111110111;
  assign mem[825] = 14'b00001100001100;
  assign mem[826] = 14'b01001001111101;
  assign mem[827] = 14'b01001000001111;
  assign mem[828] = 14'b00100001010110;
  assign mem[829] = 14'b00100000100111;
  assign mem[830] = 14'b01001011000010;
  assign mem[831] = 14'b00001101110100;
  assign mem[832] = 14'b01010011111100;
  assign mem[833] = 14'b01011010100011;
  assign mem[834] = 14'b01011100110010;
  assign mem[835] = 14'b01000011101101;
  assign mem[836] = 14'b01100110011111;
  assign mem[837] = 14'b01110101111101;
  assign mem[838] = 14'b01010010010101;
  assign mem[839] = 14'b10100110101000;
  assign mem[840] = 14'b01000010011100;
  assign mem[841] = 14'b00110010111100;
  assign mem[842] = 14'b01011100011101;
  assign mem[843] = 14'b10101000111110;
  assign mem[844] = 14'b01011010001000;
  assign mem[845] = 14'b10011011111111;
  assign mem[846] = 14'b01111110100000;
  assign mem[847] = 14'b01111001101111;
  assign mem[848] = 14'b01101010010000;
  assign mem[849] = 14'b01110101000011;
  assign mem[850] = 14'b01100010000000;
  assign mem[851] = 14'b00011101110011;
  assign mem[852] = 14'b10101011000011;
  assign mem[853] = 14'b01100010010001;
  assign mem[854] = 14'b10111000011011;
  assign mem[855] = 14'b01011110010000;
  assign mem[856] = 14'b10110010111001;
  assign mem[857] = 14'b00010010010011;
  assign mem[858] = 14'b10001111110001;
  assign mem[859] = 14'b01111011111101;
  assign mem[860] = 14'b00100110101111;
  assign mem[861] = 14'b01111100100010;
  assign mem[862] = 14'b10110001001001;
  assign mem[863] = 14'b01101110010110;
  assign mem[864] = 14'b10001011001111;
  assign mem[865] = 14'b01101001001000;
  assign mem[866] = 14'b01100110001110;
  assign mem[867] = 14'b01111110110010;
  assign mem[868] = 14'b10001001111100;
  assign mem[869] = 14'b01100111000011;
  assign mem[870] = 14'b00110111011001;
  assign mem[871] = 14'b01000011111100;
  assign mem[872] = 14'b01001000000010;
  assign mem[873] = 14'b00100010011101;
  assign mem[874] = 14'b01101101010111;
  assign mem[875] = 14'b01111110101010;
  assign mem[876] = 14'b01010110111000;
  assign mem[877] = 14'b10100010010110;
  assign mem[878] = 14'b10010001101001;
  assign mem[879] = 14'b00100111000011;
  assign mem[880] = 14'b00100101101101;
  assign mem[881] = 14'b01110001101000;
  assign mem[882] = 14'b01101011100001;
  assign mem[883] = 14'b10100101010110;
  assign mem[884] = 14'b10010001011100;
  assign mem[885] = 14'b10010011011101;
  assign mem[886] = 14'b00110111100010;
  assign mem[887] = 14'b00110011111110;
  assign mem[888] = 14'b01011101100111;
  assign mem[889] = 14'b10111011000001;
  assign mem[890] = 14'b00110101010111;
  assign mem[891] = 14'b10111111111011;
  assign mem[892] = 14'b10011001101110;
  assign mem[893] = 14'b10111100011111;
  assign mem[894] = 14'b01000011101100;
  assign mem[895] = 14'b01111010010110;
  assign mem[896] = 14'b10110001000001;
  assign mem[897] = 14'b01100111001101;
  assign mem[898] = 14'b10111111101111;
  assign mem[899] = 14'b00011111111100;
  assign mem[900] = 14'b10110101011011;
  assign mem[901] = 14'b01110010111001;
  assign mem[902] = 14'b10101111000001;
  assign mem[903] = 14'b10110100111110;
  assign mem[904] = 14'b00111010010101;
  assign mem[905] = 14'b10001011101111;
  assign mem[906] = 14'b10011011111010;
  assign mem[907] = 14'b00011001011011;
  assign mem[908] = 14'b01110000000000;
  assign mem[909] = 14'b00111101011111;
  assign mem[910] = 14'b01001110111010;
  assign mem[911] = 14'b00101011001010;
  assign mem[912] = 14'b01110101001000;
  assign mem[913] = 14'b10100010001111;
  assign mem[914] = 14'b00001011110011;
  assign mem[915] = 14'b00011001110110;
  assign mem[916] = 14'b10111100010101;
  assign mem[917] = 14'b01001101011000;
  assign mem[918] = 14'b10011110010110;
  assign mem[919] = 14'b01000100101010;
  assign mem[920] = 14'b01100111000000;
  assign mem[921] = 14'b01111011011010;
  assign mem[922] = 14'b01110101001001;
  assign mem[923] = 14'b10001011001000;
  assign mem[924] = 14'b10111011111101;
  assign mem[925] = 14'b00110111111101;
  assign mem[926] = 14'b10100111111100;
  assign mem[927] = 14'b01011000101010;
  assign mem[928] = 14'b10100001110110;
  assign mem[929] = 14'b01001100100101;
  assign mem[930] = 14'b01110011110110;
  assign mem[931] = 14'b10001001000011;
  assign mem[932] = 14'b00001011000110;
  assign mem[933] = 14'b01101001101100;
  assign mem[934] = 14'b10000100001110;
  assign mem[935] = 14'b01110000011001;
  assign mem[936] = 14'b01010011111011;
  assign mem[937] = 14'b01110001101010;
  assign mem[938] = 14'b10101101001100;
  assign mem[939] = 14'b00000100100010;
  assign mem[940] = 14'b01111010111000;
  assign mem[941] = 14'b01101010101011;
  assign mem[942] = 14'b10111000101110;
  assign mem[943] = 14'b00100111001101;
  assign mem[944] = 14'b01100110110010;
  assign mem[945] = 14'b00111110111010;
  assign mem[946] = 14'b01011010101111;
  assign mem[947] = 14'b00010110110010;
  assign mem[948] = 14'b01011001011001;
  assign mem[949] = 14'b01011010000010;
  assign mem[950] = 14'b01000001010010;
  assign mem[951] = 14'b00100000111001;
  assign mem[952] = 14'b10110101100101;
  assign mem[953] = 14'b01001011110100;
  assign mem[954] = 14'b10001011000001;
  assign mem[955] = 14'b00101100101000;
  assign mem[956] = 14'b10110011110110;
  assign mem[957] = 14'b10010000110000;
  assign mem[958] = 14'b00100111011000;
  assign mem[959] = 14'b10001001001000;
  assign mem[960] = 14'b01101101100011;
  assign mem[961] = 14'b00101001010111;
  assign mem[962] = 14'b00011101101010;
  assign mem[963] = 14'b01101101111111;
  assign mem[964] = 14'b01011100111110;
  assign mem[965] = 14'b10101110011011;
  assign mem[966] = 14'b01010101110000;
  assign mem[967] = 14'b01100010000101;
  assign mem[968] = 14'b10001111011110;
  assign mem[969] = 14'b10110011000000;
  assign mem[970] = 14'b00001001111001;
  assign mem[971] = 14'b10011100111110;
  assign mem[972] = 14'b10110100100010;
  assign mem[973] = 14'b01011000000001;
  assign mem[974] = 14'b10010101110011;
  assign mem[975] = 14'b00100100011101;
  assign mem[976] = 14'b01101101100000;
  assign mem[977] = 14'b01101110101100;
  assign mem[978] = 14'b01001110110111;
  assign mem[979] = 14'b01110000011111;
  assign mem[980] = 14'b10011010001001;
  assign mem[981] = 14'b10001100100101;
  assign mem[982] = 14'b00001000111001;
  assign mem[983] = 14'b01100011110110;
  assign mem[984] = 14'b10101001011101;
  assign mem[985] = 14'b10010111001111;
  assign mem[986] = 14'b10000001001100;
  assign mem[987] = 14'b10110011010000;
  assign mem[988] = 14'b01000001101011;
  assign mem[989] = 14'b00011111001101;
  assign mem[990] = 14'b00000000000010;
  assign mem[991] = 14'b10010001110011;
  assign mem[992] = 14'b00000010100010;
  assign mem[993] = 14'b01100000100110;
  assign mem[994] = 14'b00011111010000;
  assign mem[995] = 14'b00111001000001;
  assign mem[996] = 14'b10011001000000;
  assign mem[997] = 14'b01100011011011;
  assign mem[998] = 14'b01110110000101;
  assign mem[999] = 14'b01100000101011;
  assign mem[1000] = 14'b10000100111110;
  assign mem[1001] = 14'b10011011001111;
  assign mem[1002] = 14'b01010110100000;
  assign mem[1003] = 14'b10001100111011;
  assign mem[1004] = 14'b00111001111010;
  assign mem[1005] = 14'b10111011101001;
  assign mem[1006] = 14'b00010110101100;
  assign mem[1007] = 14'b00101111111011;
  assign mem[1008] = 14'b01010101110110;
  assign mem[1009] = 14'b10010111011100;
  assign mem[1010] = 14'b01001100000001;
  assign mem[1011] = 14'b01011110000011;
  assign mem[1012] = 14'b01101111000010;
  assign mem[1013] = 14'b10010110001010;
  assign mem[1014] = 14'b01000111101100;
  assign mem[1015] = 14'b10011110110101;
  assign mem[1016] = 14'b01100001110101;
  assign mem[1017] = 14'b01011011111111;
  assign mem[1018] = 14'b00101001011100;
  assign mem[1019] = 14'b10011110111100;
  assign mem[1020] = 14'b00011000101100;
  assign mem[1021] = 14'b10100010001011;
  assign mem[1022] = 14'b01001000011110;
  assign mem[1023] = 14'b10011011011101;

  always@(*)
  begin
    data_out_t <= mem[addr_f];
  end

  // Build output registers
  wire [13:0] data_out_reg [n_outreg:0];
  generate if (n_outreg > 0)
  begin
    for( i=n_outreg-1; i >= 1; i=i-1)
    begin: data_out_reg_stage
      mgc_generic_reg #(
        .width(14), 
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_data_out_reg (
        .d(data_out_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(data_out_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(14), 
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_data_out_reg_init (
      .d(data_out_t),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(data_out_reg[0])
    );
    assign data_out = data_out_reg[n_outreg-1];
  end
  else
  begin
    assign data_out = data_out_t;
  end
  endgenerate

endmodule



//------> ./rtl_stagemgc_rom_sync_regout_11_1024_14_1_0_0_1_0_1_0_0_0_1_60.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Sun Oct  6 01:48:34 2024
// ----------------------------------------------------------------------

// 
module stagemgc_rom_sync_regout_11_1024_14_1_0_0_1_0_1_0_0_0_1_60 (addr, data_out,
    clk, s_rst, a_rst, en
);
  input [9:0]addr ;
  output [13:0]data_out ;
  input clk ;
  input s_rst ;
  input a_rst ;
  input en ;


  // Constants for ROM dimensions
  parameter n_width    = 14;
  parameter n_size     = 1024;
  parameter n_numports = 1;
  parameter n_addr_w   = 10;
  parameter n_inreg    = 0;
  parameter n_outreg   = 1;
  wire [9:0] addr_f;

  // Build input address registers
  wire [9:0] addr_reg [n_inreg:0];
  genvar i;
  generate if (n_inreg > 0)
  begin
    for( i=n_inreg-1; i >= 1; i=i-1)
    begin: addr_reg_stage
      mgc_generic_reg #(
        .width(10), 
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_addr_reg (
        .d(addr_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(addr_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(10), 
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_addr_reg_init (
      .d(addr),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(addr_reg[0])
    );
    assign addr_f = addr_reg[n_inreg-1];
  end
  else
  begin
    assign addr_f = addr;
  end
  endgenerate

  // Declare storage for memory elements
  wire [13:0] mem [1023:0];

  // Declare output registers
  reg [13:0] data_out_t;

  // Initialize ROM contents
  assign mem[0] = 14'b00111111111011;
  assign mem[1] = 14'b01000100110001;
  assign mem[2] = 14'b00010000111001;
  assign mem[3] = 14'b00010011001101;
  assign mem[4] = 14'b00100111100010;
  assign mem[5] = 14'b01011101111110;
  assign mem[6] = 14'b01111100001011;
  assign mem[7] = 14'b01010011010001;
  assign mem[8] = 14'b00101000010011;
  assign mem[9] = 14'b01001010001111;
  assign mem[10] = 14'b01100101000000;
  assign mem[11] = 14'b10110110110111;
  assign mem[12] = 14'b01101101101111;
  assign mem[13] = 14'b00101011111100;
  assign mem[14] = 14'b01011100000010;
  assign mem[15] = 14'b10100111001010;
  assign mem[16] = 14'b00110000100101;
  assign mem[17] = 14'b00100001001101;
  assign mem[18] = 14'b00011110101000;
  assign mem[19] = 14'b10101010101101;
  assign mem[20] = 14'b10100101101001;
  assign mem[21] = 14'b10100010100100;
  assign mem[22] = 14'b01000001011101;
  assign mem[23] = 14'b00011101010011;
  assign mem[24] = 14'b01011011010111;
  assign mem[25] = 14'b10000101100010;
  assign mem[26] = 14'b01001000000111;
  assign mem[27] = 14'b01010001000110;
  assign mem[28] = 14'b10110000111100;
  assign mem[29] = 14'b10100101010010;
  assign mem[30] = 14'b01011011111010;
  assign mem[31] = 14'b10101110010011;
  assign mem[32] = 14'b10000011100001;
  assign mem[33] = 14'b10111111110011;
  assign mem[34] = 14'b10100101100111;
  assign mem[35] = 14'b01110100010110;
  assign mem[36] = 14'b01011001010111;
  assign mem[37] = 14'b00110111110001;
  assign mem[38] = 14'b01011101011101;
  assign mem[39] = 14'b10011101111100;
  assign mem[40] = 14'b01000101001010;
  assign mem[41] = 14'b10000001110010;
  assign mem[42] = 14'b10101000000011;
  assign mem[43] = 14'b01001001000111;
  assign mem[44] = 14'b10101100101100;
  assign mem[45] = 14'b00011000000010;
  assign mem[46] = 14'b10111001010001;
  assign mem[47] = 14'b00000001100100;
  assign mem[48] = 14'b10000000110111;
  assign mem[49] = 14'b01100111100001;
  assign mem[50] = 14'b10010111111101;
  assign mem[51] = 14'b01010000011001;
  assign mem[52] = 14'b00110101010100;
  assign mem[53] = 14'b01111010110010;
  assign mem[54] = 14'b01011011000111;
  assign mem[55] = 14'b10010011110100;
  assign mem[56] = 14'b01010001100001;
  assign mem[57] = 14'b10100111110100;
  assign mem[58] = 14'b01111011001010;
  assign mem[59] = 14'b01110101010010;
  assign mem[60] = 14'b10111110001100;
  assign mem[61] = 14'b10110000011100;
  assign mem[62] = 14'b01011110100001;
  assign mem[63] = 14'b00000001001111;
  assign mem[64] = 14'b00000000001101;
  assign mem[65] = 14'b01101100011010;
  assign mem[66] = 14'b10001010110110;
  assign mem[67] = 14'b01010101001101;
  assign mem[68] = 14'b01000111101010;
  assign mem[69] = 14'b10110010111111;
  assign mem[70] = 14'b00101101010111;
  assign mem[71] = 14'b01001001000100;
  assign mem[72] = 14'b10011001110011;
  assign mem[73] = 14'b01110111000101;
  assign mem[74] = 14'b10001001110110;
  assign mem[75] = 14'b10001110010101;
  assign mem[76] = 14'b00100000100011;
  assign mem[77] = 14'b10000100111011;
  assign mem[78] = 14'b10000111101101;
  assign mem[79] = 14'b00110000100110;
  assign mem[80] = 14'b01101101100111;
  assign mem[81] = 14'b00110011000101;
  assign mem[82] = 14'b00010101010111;
  assign mem[83] = 14'b01100011111101;
  assign mem[84] = 14'b10100000010011;
  assign mem[85] = 14'b10000011110011;
  assign mem[86] = 14'b10100100011111;
  assign mem[87] = 14'b10110100100111;
  assign mem[88] = 14'b10101101010110;
  assign mem[89] = 14'b00100010100011;
  assign mem[90] = 14'b00011100010000;
  assign mem[91] = 14'b01110010010111;
  assign mem[92] = 14'b00000000110000;
  assign mem[93] = 14'b10010101001011;
  assign mem[94] = 14'b00101000000000;
  assign mem[95] = 14'b00010011001100;
  assign mem[96] = 14'b10010011011110;
  assign mem[97] = 14'b10101000100011;
  assign mem[98] = 14'b10111000011000;
  assign mem[99] = 14'b00011100011100;
  assign mem[100] = 14'b10110010001110;
  assign mem[101] = 14'b10001100000110;
  assign mem[102] = 14'b01100000001111;
  assign mem[103] = 14'b00101111000100;
  assign mem[104] = 14'b01011111011101;
  assign mem[105] = 14'b00101011101100;
  assign mem[106] = 14'b00100010011011;
  assign mem[107] = 14'b00011001110100;
  assign mem[108] = 14'b00001011000111;
  assign mem[109] = 14'b01101101011100;
  assign mem[110] = 14'b00010000011101;
  assign mem[111] = 14'b10001100001101;
  assign mem[112] = 14'b01010001111100;
  assign mem[113] = 14'b00010111101101;
  assign mem[114] = 14'b10010001101010;
  assign mem[115] = 14'b10110000000101;
  assign mem[116] = 14'b00001110000100;
  assign mem[117] = 14'b00111100110000;
  assign mem[118] = 14'b10101101111101;
  assign mem[119] = 14'b10100111110000;
  assign mem[120] = 14'b01001101010101;
  assign mem[121] = 14'b01110111000000;
  assign mem[122] = 14'b10011011110110;
  assign mem[123] = 14'b01001010001010;
  assign mem[124] = 14'b10100000011110;
  assign mem[125] = 14'b00000001111110;
  assign mem[126] = 14'b00101101101001;
  assign mem[127] = 14'b01101001000000;
  assign mem[128] = 14'b01100111101011;
  assign mem[129] = 14'b01100110001111;
  assign mem[130] = 14'b00011000101110;
  assign mem[131] = 14'b01001100000100;
  assign mem[132] = 14'b00000000101010;
  assign mem[133] = 14'b00001010100001;
  assign mem[134] = 14'b00100011000000;
  assign mem[135] = 14'b01110000110011;
  assign mem[136] = 14'b00010100010000;
  assign mem[137] = 14'b10111011010101;
  assign mem[138] = 14'b01110111111011;
  assign mem[139] = 14'b10000110000010;
  assign mem[140] = 14'b10111010101101;
  assign mem[141] = 14'b00001111011101;
  assign mem[142] = 14'b10100100101101;
  assign mem[143] = 14'b01111000000111;
  assign mem[144] = 14'b01101110101101;
  assign mem[145] = 14'b10000100100111;
  assign mem[146] = 14'b00001111101100;
  assign mem[147] = 14'b10011111111100;
  assign mem[148] = 14'b01001001011111;
  assign mem[149] = 14'b00000010100011;
  assign mem[150] = 14'b10001110110111;
  assign mem[151] = 14'b01000111110101;
  assign mem[152] = 14'b01100100011111;
  assign mem[153] = 14'b10111100010100;
  assign mem[154] = 14'b00101110101111;
  assign mem[155] = 14'b10111010100010;
  assign mem[156] = 14'b01001000100111;
  assign mem[157] = 14'b00110100100010;
  assign mem[158] = 14'b00100000001100;
  assign mem[159] = 14'b10110001011101;
  assign mem[160] = 14'b10111011101011;
  assign mem[161] = 14'b01101000001000;
  assign mem[162] = 14'b01011000010111;
  assign mem[163] = 14'b01110000111001;
  assign mem[164] = 14'b01011100011010;
  assign mem[165] = 14'b10010001101111;
  assign mem[166] = 14'b00111111111100;
  assign mem[167] = 14'b01011011111000;
  assign mem[168] = 14'b01101100010100;
  assign mem[169] = 14'b00110101001010;
  assign mem[170] = 14'b01010000001101;
  assign mem[171] = 14'b10010010110010;
  assign mem[172] = 14'b10101111011101;
  assign mem[173] = 14'b01010010000100;
  assign mem[174] = 14'b10001100110000;
  assign mem[175] = 14'b00011000010100;
  assign mem[176] = 14'b01101011111100;
  assign mem[177] = 14'b01001010100101;
  assign mem[178] = 14'b00111100001101;
  assign mem[179] = 14'b10001001001100;
  assign mem[180] = 14'b10100001010101;
  assign mem[181] = 14'b01111000111001;
  assign mem[182] = 14'b00011011011110;
  assign mem[183] = 14'b01101110111111;
  assign mem[184] = 14'b10110001101111;
  assign mem[185] = 14'b10111111110001;
  assign mem[186] = 14'b10000110011010;
  assign mem[187] = 14'b00110010101011;
  assign mem[188] = 14'b01100110001000;
  assign mem[189] = 14'b01110110100110;
  assign mem[190] = 14'b10000110001111;
  assign mem[191] = 14'b10110100100000;
  assign mem[192] = 14'b01011111010101;
  assign mem[193] = 14'b00110010110101;
  assign mem[194] = 14'b10011011110001;
  assign mem[195] = 14'b10010110101000;
  assign mem[196] = 14'b01000110011010;
  assign mem[197] = 14'b00111010011000;
  assign mem[198] = 14'b01101010101101;
  assign mem[199] = 14'b10101001000110;
  assign mem[200] = 14'b10001110101010;
  assign mem[201] = 14'b10011011011100;
  assign mem[202] = 14'b00110111101110;
  assign mem[203] = 14'b00100001010101;
  assign mem[204] = 14'b00111100111101;
  assign mem[205] = 14'b01011110010110;
  assign mem[206] = 14'b01110010100101;
  assign mem[207] = 14'b01100111010001;
  assign mem[208] = 14'b00110110001100;
  assign mem[209] = 14'b01001000110011;
  assign mem[210] = 14'b00001001110001;
  assign mem[211] = 14'b00101010001100;
  assign mem[212] = 14'b01111000111010;
  assign mem[213] = 14'b00110101110011;
  assign mem[214] = 14'b00101111110100;
  assign mem[215] = 14'b00110100111100;
  assign mem[216] = 14'b00110111000110;
  assign mem[217] = 14'b01000101000010;
  assign mem[218] = 14'b10111010000111;
  assign mem[219] = 14'b01100001011000;
  assign mem[220] = 14'b00011011000010;
  assign mem[221] = 14'b00100111111110;
  assign mem[222] = 14'b10100001100100;
  assign mem[223] = 14'b01010011100000;
  assign mem[224] = 14'b01010010100110;
  assign mem[225] = 14'b00100010001110;
  assign mem[226] = 14'b10110100101010;
  assign mem[227] = 14'b01100000110111;
  assign mem[228] = 14'b00100110110010;
  assign mem[229] = 14'b10001000110100;
  assign mem[230] = 14'b01010100001011;
  assign mem[231] = 14'b01000000000101;
  assign mem[232] = 14'b01001000000001;
  assign mem[233] = 14'b10000110011101;
  assign mem[234] = 14'b10000000100010;
  assign mem[235] = 14'b00000010010000;
  assign mem[236] = 14'b01011000011000;
  assign mem[237] = 14'b10001000000000;
  assign mem[238] = 14'b00101000111101;
  assign mem[239] = 14'b01010100110000;
  assign mem[240] = 14'b10101000111100;
  assign mem[241] = 14'b00101110001111;
  assign mem[242] = 14'b10110001010010;
  assign mem[243] = 14'b01100001101001;
  assign mem[244] = 14'b00011010110011;
  assign mem[245] = 14'b01001101010111;
  assign mem[246] = 14'b10010101000100;
  assign mem[247] = 14'b00011101100000;
  assign mem[248] = 14'b00111010110100;
  assign mem[249] = 14'b00000000100111;
  assign mem[250] = 14'b10000000011011;
  assign mem[251] = 14'b00100000100000;
  assign mem[252] = 14'b00100111000110;
  assign mem[253] = 14'b00010110111101;
  assign mem[254] = 14'b10100100110110;
  assign mem[255] = 14'b10001000000101;
  assign mem[256] = 14'b01010111100001;
  assign mem[257] = 14'b00010001000101;
  assign mem[258] = 14'b00111011001000;
  assign mem[259] = 14'b01001110110001;
  assign mem[260] = 14'b00100000001010;
  assign mem[261] = 14'b10000011001111;
  assign mem[262] = 14'b10110010111000;
  assign mem[263] = 14'b10010110100111;
  assign mem[264] = 14'b00100000001011;
  assign mem[265] = 14'b10011010010110;
  assign mem[266] = 14'b01110011101101;
  assign mem[267] = 14'b00100111000000;
  assign mem[268] = 14'b01111011101110;
  assign mem[269] = 14'b10110101001010;
  assign mem[270] = 14'b00000101110011;
  assign mem[271] = 14'b01111100111001;
  assign mem[272] = 14'b00110000000001;
  assign mem[273] = 14'b10100001010110;
  assign mem[274] = 14'b00000000101000;
  assign mem[275] = 14'b10011100010100;
  assign mem[276] = 14'b10010000011101;
  assign mem[277] = 14'b01111100110011;
  assign mem[278] = 14'b01010111100011;
  assign mem[279] = 14'b00111111010011;
  assign mem[280] = 14'b01111011010110;
  assign mem[281] = 14'b00001010100100;
  assign mem[282] = 14'b10110001110100;
  assign mem[283] = 14'b01110011010011;
  assign mem[284] = 14'b01100101100101;
  assign mem[285] = 14'b01001101110101;
  assign mem[286] = 14'b00101001000100;
  assign mem[287] = 14'b00110110100000;
  assign mem[288] = 14'b10101011001100;
  assign mem[289] = 14'b01101101101110;
  assign mem[290] = 14'b01101001010001;
  assign mem[291] = 14'b10011011001101;
  assign mem[292] = 14'b01101111100011;
  assign mem[293] = 14'b00100100011010;
  assign mem[294] = 14'b00111100101100;
  assign mem[295] = 14'b01010101100001;
  assign mem[296] = 14'b01111010111001;
  assign mem[297] = 14'b01101100011101;
  assign mem[298] = 14'b01011001101001;
  assign mem[299] = 14'b01010111101101;
  assign mem[300] = 14'b10010100100001;
  assign mem[301] = 14'b10110100110000;
  assign mem[302] = 14'b10110000001101;
  assign mem[303] = 14'b00100111001110;
  assign mem[304] = 14'b01101000100001;
  assign mem[305] = 14'b00000110000010;
  assign mem[306] = 14'b01000101101110;
  assign mem[307] = 14'b00000001101001;
  assign mem[308] = 14'b00100000011100;
  assign mem[309] = 14'b10100011001011;
  assign mem[310] = 14'b00000001110111;
  assign mem[311] = 14'b00111101110011;
  assign mem[312] = 14'b01000100010010;
  assign mem[313] = 14'b10110011110001;
  assign mem[314] = 14'b00111001011000;
  assign mem[315] = 14'b10110010101111;
  assign mem[316] = 14'b00001011101110;
  assign mem[317] = 14'b00110010101000;
  assign mem[318] = 14'b00110000111101;
  assign mem[319] = 14'b00001011110010;
  assign mem[320] = 14'b00111110101101;
  assign mem[321] = 14'b10111010011001;
  assign mem[322] = 14'b10001111111010;
  assign mem[323] = 14'b01010100000010;
  assign mem[324] = 14'b10111001101001;
  assign mem[325] = 14'b10101100001010;
  assign mem[326] = 14'b00101100000010;
  assign mem[327] = 14'b00011100111011;
  assign mem[328] = 14'b01001101100110;
  assign mem[329] = 14'b01111111110101;
  assign mem[330] = 14'b00101010000000;
  assign mem[331] = 14'b01100000111101;
  assign mem[332] = 14'b01101010011110;
  assign mem[333] = 14'b00001110011110;
  assign mem[334] = 14'b00101101111000;
  assign mem[335] = 14'b01000011100111;
  assign mem[336] = 14'b10011110111111;
  assign mem[337] = 14'b01101110110001;
  assign mem[338] = 14'b01011110011111;
  assign mem[339] = 14'b10010011000010;
  assign mem[340] = 14'b10100011111100;
  assign mem[341] = 14'b10001011110110;
  assign mem[342] = 14'b00100110101000;
  assign mem[343] = 14'b01100001101111;
  assign mem[344] = 14'b00001011011000;
  assign mem[345] = 14'b01110110010001;
  assign mem[346] = 14'b01011110101000;
  assign mem[347] = 14'b10100011000000;
  assign mem[348] = 14'b10101100011100;
  assign mem[349] = 14'b00100110010100;
  assign mem[350] = 14'b00101011111011;
  assign mem[351] = 14'b00111011001011;
  assign mem[352] = 14'b00001110110001;
  assign mem[353] = 14'b10001100100110;
  assign mem[354] = 14'b00010011011100;
  assign mem[355] = 14'b10001001101111;
  assign mem[356] = 14'b10101100001001;
  assign mem[357] = 14'b10101111010010;
  assign mem[358] = 14'b01011100000110;
  assign mem[359] = 14'b01000011100101;
  assign mem[360] = 14'b01001000011111;
  assign mem[361] = 14'b00111011101011;
  assign mem[362] = 14'b10011001100010;
  assign mem[363] = 14'b01101110010000;
  assign mem[364] = 14'b01101010000010;
  assign mem[365] = 14'b10000111011110;
  assign mem[366] = 14'b01010110100011;
  assign mem[367] = 14'b01111000011011;
  assign mem[368] = 14'b00010101010001;
  assign mem[369] = 14'b10011001010100;
  assign mem[370] = 14'b00101110000101;
  assign mem[371] = 14'b10110000000001;
  assign mem[372] = 14'b10100000111101;
  assign mem[373] = 14'b10001110010100;
  assign mem[374] = 14'b00000111011110;
  assign mem[375] = 14'b01100101011001;
  assign mem[376] = 14'b00000001100101;
  assign mem[377] = 14'b00011101110111;
  assign mem[378] = 14'b10010100001011;
  assign mem[379] = 14'b00111000011000;
  assign mem[380] = 14'b10111011011101;
  assign mem[381] = 14'b10100100101000;
  assign mem[382] = 14'b00001100101100;
  assign mem[383] = 14'b10001011010011;
  assign mem[384] = 14'b00001001111101;
  assign mem[385] = 14'b01111111011111;
  assign mem[386] = 14'b01010010110011;
  assign mem[387] = 14'b10001110101000;
  assign mem[388] = 14'b00110110111000;
  assign mem[389] = 14'b10000001100010;
  assign mem[390] = 14'b01101110011100;
  assign mem[391] = 14'b01111011110010;
  assign mem[392] = 14'b00101111011100;
  assign mem[393] = 14'b01001010010111;
  assign mem[394] = 14'b00100001110011;
  assign mem[395] = 14'b00111101100001;
  assign mem[396] = 14'b00111010101011;
  assign mem[397] = 14'b10110000101010;
  assign mem[398] = 14'b01111000111011;
  assign mem[399] = 14'b01001100111010;
  assign mem[400] = 14'b10111010011100;
  assign mem[401] = 14'b00000110101000;
  assign mem[402] = 14'b01010110100010;
  assign mem[403] = 14'b01100001010100;
  assign mem[404] = 14'b10101101111011;
  assign mem[405] = 14'b01111001100010;
  assign mem[406] = 14'b10111011000110;
  assign mem[407] = 14'b00010001001001;
  assign mem[408] = 14'b00101101001010;
  assign mem[409] = 14'b10011100101011;
  assign mem[410] = 14'b00101000001001;
  assign mem[411] = 14'b00100011001010;
  assign mem[412] = 14'b00100100110000;
  assign mem[413] = 14'b00001100110101;
  assign mem[414] = 14'b00100111110110;
  assign mem[415] = 14'b10101100001000;
  assign mem[416] = 14'b01111001011001;
  assign mem[417] = 14'b00000010001000;
  assign mem[418] = 14'b00001001101001;
  assign mem[419] = 14'b00110001010101;
  assign mem[420] = 14'b01011100000001;
  assign mem[421] = 14'b10010000000011;
  assign mem[422] = 14'b01101011000111;
  assign mem[423] = 14'b00000001111000;
  assign mem[424] = 14'b01000100110101;
  assign mem[425] = 14'b00011100100001;
  assign mem[426] = 14'b10010110100011;
  assign mem[427] = 14'b01110000101110;
  assign mem[428] = 14'b10100000010101;
  assign mem[429] = 14'b10110010000001;
  assign mem[430] = 14'b00100110001001;
  assign mem[431] = 14'b10010101011010;
  assign mem[432] = 14'b10101110101000;
  assign mem[433] = 14'b00001001010111;
  assign mem[434] = 14'b00100000100101;
  assign mem[435] = 14'b10110011001001;
  assign mem[436] = 14'b01110001000001;
  assign mem[437] = 14'b01100000100001;
  assign mem[438] = 14'b01001011000001;
  assign mem[439] = 14'b10011011000110;
  assign mem[440] = 14'b10001100110010;
  assign mem[441] = 14'b01000110100010;
  assign mem[442] = 14'b10010011101111;
  assign mem[443] = 14'b10110001011000;
  assign mem[444] = 14'b10110110010110;
  assign mem[445] = 14'b01100000011110;
  assign mem[446] = 14'b01111100001110;
  assign mem[447] = 14'b10011000100110;
  assign mem[448] = 14'b01101011110000;
  assign mem[449] = 14'b10110101010011;
  assign mem[450] = 14'b00110010001101;
  assign mem[451] = 14'b10000100011001;
  assign mem[452] = 14'b10011010010001;
  assign mem[453] = 14'b00101100010011;
  assign mem[454] = 14'b10100010110110;
  assign mem[455] = 14'b00111010010100;
  assign mem[456] = 14'b01111100011001;
  assign mem[457] = 14'b00010110110001;
  assign mem[458] = 14'b10101001101001;
  assign mem[459] = 14'b01111110000101;
  assign mem[460] = 14'b00001101000000;
  assign mem[461] = 14'b00011001011100;
  assign mem[462] = 14'b00110101010010;
  assign mem[463] = 14'b01001100100100;
  assign mem[464] = 14'b10101001100111;
  assign mem[465] = 14'b01001111110111;
  assign mem[466] = 14'b10010101000111;
  assign mem[467] = 14'b01100010110101;
  assign mem[468] = 14'b01110100000111;
  assign mem[469] = 14'b00111111110011;
  assign mem[470] = 14'b00110000000000;
  assign mem[471] = 14'b10001010001111;
  assign mem[472] = 14'b10011001111101;
  assign mem[473] = 14'b10011110001010;
  assign mem[474] = 14'b01010010001011;
  assign mem[475] = 14'b10110010010101;
  assign mem[476] = 14'b01100110011100;
  assign mem[477] = 14'b00000100101111;
  assign mem[478] = 14'b00010110111001;
  assign mem[479] = 14'b00111100011111;
  assign mem[480] = 14'b01001100001001;
  assign mem[481] = 14'b01011010110101;
  assign mem[482] = 14'b10011100100001;
  assign mem[483] = 14'b01101011110010;
  assign mem[484] = 14'b00110011101111;
  assign mem[485] = 14'b01011100111011;
  assign mem[486] = 14'b10000110111101;
  assign mem[487] = 14'b01011011011100;
  assign mem[488] = 14'b00111100010000;
  assign mem[489] = 14'b00001110100000;
  assign mem[490] = 14'b01001101000101;
  assign mem[491] = 14'b10000101010010;
  assign mem[492] = 14'b00011101001111;
  assign mem[493] = 14'b00100010001000;
  assign mem[494] = 14'b01010111000011;
  assign mem[495] = 14'b01011011110111;
  assign mem[496] = 14'b00110110011001;
  assign mem[497] = 14'b10110101001101;
  assign mem[498] = 14'b10010100100111;
  assign mem[499] = 14'b01111111011001;
  assign mem[500] = 14'b00000000100011;
  assign mem[501] = 14'b00101000110001;
  assign mem[502] = 14'b01011101001011;
  assign mem[503] = 14'b01111110000000;
  assign mem[504] = 14'b00010000111000;
  assign mem[505] = 14'b10111100000111;
  assign mem[506] = 14'b10000011111100;
  assign mem[507] = 14'b00101111101100;
  assign mem[508] = 14'b00111011100101;
  assign mem[509] = 14'b10101100111001;
  assign mem[510] = 14'b01101001010000;
  assign mem[511] = 14'b10000100000110;
  assign mem[512] = 14'b00100100100100;
  assign mem[513] = 14'b01110111100011;
  assign mem[514] = 14'b00011101110110;
  assign mem[515] = 14'b10100111010101;
  assign mem[516] = 14'b00100001000101;
  assign mem[517] = 14'b10010110100101;
  assign mem[518] = 14'b01100100000010;
  assign mem[519] = 14'b01011110001100;
  assign mem[520] = 14'b00100001001100;
  assign mem[521] = 14'b01111000010101;
  assign mem[522] = 14'b00101001110111;
  assign mem[523] = 14'b01010000111111;
  assign mem[524] = 14'b01100001111110;
  assign mem[525] = 14'b01110100000000;
  assign mem[526] = 14'b00101000100101;
  assign mem[527] = 14'b01101010001011;
  assign mem[528] = 14'b10010000000110;
  assign mem[529] = 14'b10101001010101;
  assign mem[530] = 14'b00000100011000;
  assign mem[531] = 14'b10000110000111;
  assign mem[532] = 14'b00110011000110;
  assign mem[533] = 14'b01101001100001;
  assign mem[534] = 14'b00100100110010;
  assign mem[535] = 14'b00111011000011;
  assign mem[536] = 14'b01011111010110;
  assign mem[537] = 14'b01001001111100;
  assign mem[538] = 14'b01011100100110;
  assign mem[539] = 14'b00100111000001;
  assign mem[540] = 14'b10000111000000;
  assign mem[541] = 14'b10100000110001;
  assign mem[542] = 14'b01011111011011;
  assign mem[543] = 14'b10111101011111;
  assign mem[544] = 14'b00101110001110;
  assign mem[545] = 14'b10111111111111;
  assign mem[546] = 14'b10100000110100;
  assign mem[547] = 14'b01111110010110;
  assign mem[548] = 14'b00001100110001;
  assign mem[549] = 14'b00111110110101;
  assign mem[550] = 14'b00101000110010;
  assign mem[551] = 14'b00010110100100;
  assign mem[552] = 14'b01011100001011;
  assign mem[553] = 14'b10110111001000;
  assign mem[554] = 14'b00110011011100;
  assign mem[555] = 14'b00100101111000;
  assign mem[556] = 14'b01001111100010;
  assign mem[557] = 14'b01110001001010;
  assign mem[558] = 14'b01010001010101;
  assign mem[559] = 14'b01010010100001;
  assign mem[560] = 14'b10011011100100;
  assign mem[561] = 14'b00101010001110;
  assign mem[562] = 14'b01101000000000;
  assign mem[563] = 14'b00001011011111;
  assign mem[564] = 14'b00100011000011;
  assign mem[565] = 14'b10110110001000;
  assign mem[566] = 14'b00001101000001;
  assign mem[567] = 14'b00110000100011;
  assign mem[568] = 14'b01011101111100;
  assign mem[569] = 14'b01101010010001;
  assign mem[570] = 14'b00010001100110;
  assign mem[571] = 14'b01100011000011;
  assign mem[572] = 14'b01010010000010;
  assign mem[573] = 14'b10100010010111;
  assign mem[574] = 14'b10010110101010;
  assign mem[575] = 14'b01010010011110;
  assign mem[576] = 14'b00110110111001;
  assign mem[577] = 14'b10011000101001;
  assign mem[578] = 14'b00101111010001;
  assign mem[579] = 14'b00001100001011;
  assign mem[580] = 14'b10010011011001;
  assign mem[581] = 14'b00110101000000;
  assign mem[582] = 14'b01110100001101;
  assign mem[583] = 14'b00001010011100;
  assign mem[584] = 14'b10011111001000;
  assign mem[585] = 14'b01111110101111;
  assign mem[586] = 14'b01100101111111;
  assign mem[587] = 14'b01100110101000;
  assign mem[588] = 14'b10101001001111;
  assign mem[589] = 14'b01100101010010;
  assign mem[590] = 14'b10000001000111;
  assign mem[591] = 14'b01011001001111;
  assign mem[592] = 14'b10011000110100;
  assign mem[593] = 14'b00000111010011;
  assign mem[594] = 14'b01010101010110;
  assign mem[595] = 14'b01000101001001;
  assign mem[596] = 14'b10111011011111;
  assign mem[597] = 14'b00010010110101;
  assign mem[598] = 14'b01001110010111;
  assign mem[599] = 14'b01101100000110;
  assign mem[600] = 14'b01001111101000;
  assign mem[601] = 14'b00111011110011;
  assign mem[602] = 14'b01010110010101;
  assign mem[603] = 14'b10110100111011;
  assign mem[604] = 14'b00110110111110;
  assign mem[605] = 14'b01001100001011;
  assign mem[606] = 14'b01110011011100;
  assign mem[607] = 14'b00011110001011;
  assign mem[608] = 14'b01100111010111;
  assign mem[609] = 14'b00011000000101;
  assign mem[610] = 14'b10001000000100;
  assign mem[611] = 14'b00000100000100;
  assign mem[612] = 14'b00110100111001;
  assign mem[613] = 14'b01001010111000;
  assign mem[614] = 14'b01000100100111;
  assign mem[615] = 14'b01011001000001;
  assign mem[616] = 14'b01111011010111;
  assign mem[617] = 14'b00100001101011;
  assign mem[618] = 14'b01110010101001;
  assign mem[619] = 14'b00000011101100;
  assign mem[620] = 14'b10100110001011;
  assign mem[621] = 14'b10110100001110;
  assign mem[622] = 14'b00011101110010;
  assign mem[623] = 14'b01001010111001;
  assign mem[624] = 14'b10010100110111;
  assign mem[625] = 14'b01110001000111;
  assign mem[626] = 14'b10000010100010;
  assign mem[627] = 14'b01010000000001;
  assign mem[628] = 14'b10100110100110;
  assign mem[629] = 14'b00100100000111;
  assign mem[630] = 14'b00110100010010;
  assign mem[631] = 14'b10000101101100;
  assign mem[632] = 14'b00001011000011;
  assign mem[633] = 14'b00010001000000;
  assign mem[634] = 14'b01001101001000;
  assign mem[635] = 14'b00001010100110;
  assign mem[636] = 14'b10100000000101;
  assign mem[637] = 14'b00000000010010;
  assign mem[638] = 14'b01011000110100;
  assign mem[639] = 14'b00001111000000;
  assign mem[640] = 14'b01000101101011;
  assign mem[641] = 14'b01111100010101;
  assign mem[642] = 14'b00000011100010;
  assign mem[643] = 14'b00100110010011;
  assign mem[644] = 14'b00000000000110;
  assign mem[645] = 14'b10001010101010;
  assign mem[646] = 14'b00000101000000;
  assign mem[647] = 14'b01100010011010;
  assign mem[648] = 14'b10001100000011;
  assign mem[649] = 14'b10001000011111;
  assign mem[650] = 14'b00101100100100;
  assign mem[651] = 14'b00101110100101;
  assign mem[652] = 14'b00011010101011;
  assign mem[653] = 14'b01010100100000;
  assign mem[654] = 14'b01001110011001;
  assign mem[655] = 14'b10011010010100;
  assign mem[656] = 14'b10011000111110;
  assign mem[657] = 14'b00101110011000;
  assign mem[658] = 14'b00011101101011;
  assign mem[659] = 14'b01101001001001;
  assign mem[660] = 14'b01000001010111;
  assign mem[661] = 14'b01010010101010;
  assign mem[662] = 14'b10011101100100;
  assign mem[663] = 14'b01110111111111;
  assign mem[664] = 14'b01111100000101;
  assign mem[665] = 14'b10001000101000;
  assign mem[666] = 14'b01011000111110;
  assign mem[667] = 14'b00110110000101;
  assign mem[668] = 14'b01000001001111;
  assign mem[669] = 14'b01011001110011;
  assign mem[670] = 14'b01010110111001;
  assign mem[671] = 14'b00110100110010;
  assign mem[672] = 14'b01010001101011;
  assign mem[673] = 14'b00001110111000;
  assign mem[674] = 14'b01000011011111;
  assign mem[675] = 14'b10011001010010;
  assign mem[676] = 14'b01000100000100;
  assign mem[677] = 14'b00110000010000;
  assign mem[678] = 14'b10101101101110;
  assign mem[679] = 14'b00001101001000;
  assign mem[680] = 14'b01100001110001;
  assign mem[681] = 14'b00000111100110;
  assign mem[682] = 14'b01011101110000;
  assign mem[683] = 14'b00010100111110;
  assign mem[684] = 14'b10100010001110;
  assign mem[685] = 14'b01011110000001;
  assign mem[686] = 14'b01001010111110;
  assign mem[687] = 14'b01010101110001;
  assign mem[688] = 14'b01000110010010;
  assign mem[689] = 14'b01000001100001;
  assign mem[690] = 14'b00100100000010;
  assign mem[691] = 14'b01100101111001;
  assign mem[692] = 14'b00010111000011;
  assign mem[693] = 14'b01100011100100;
  assign mem[694] = 14'b10001101000101;
  assign mem[695] = 14'b01111101100101;
  assign mem[696] = 14'b00011001011001;
  assign mem[697] = 14'b01101101101100;
  assign mem[698] = 14'b01001010000100;
  assign mem[699] = 14'b01011001100010;
  assign mem[700] = 14'b01111100010100;
  assign mem[701] = 14'b01100011001111;
  assign mem[702] = 14'b01100101011110;
  assign mem[703] = 14'b01101100000101;
  assign mem[704] = 14'b10110010001101;
  assign mem[705] = 14'b01110100111111;
  assign mem[706] = 14'b10011111011010;
  assign mem[707] = 14'b10011110101011;
  assign mem[708] = 14'b01110111110010;
  assign mem[709] = 14'b01110110000100;
  assign mem[710] = 14'b10110011110101;
  assign mem[711] = 14'b00011000001010;
  assign mem[712] = 14'b01100110101011;
  assign mem[713] = 14'b10011111010111;
  assign mem[714] = 14'b00100011011001;
  assign mem[715] = 14'b01110010011111;
  assign mem[716] = 14'b01011011000000;
  assign mem[717] = 14'b10110010000100;
  assign mem[718] = 14'b10110100111101;
  assign mem[719] = 14'b10010111111010;
  assign mem[720] = 14'b00100011001011;
  assign mem[721] = 14'b10101110111111;
  assign mem[722] = 14'b01010011101100;
  assign mem[723] = 14'b01110011110000;
  assign mem[724] = 14'b00101100101101;
  assign mem[725] = 14'b00111110100011;
  assign mem[726] = 14'b10001111111111;
  assign mem[727] = 14'b00000111100100;
  assign mem[728] = 14'b01110101100110;
  assign mem[729] = 14'b10010011000001;
  assign mem[730] = 14'b10111111001011;
  assign mem[731] = 14'b01100000001101;
  assign mem[732] = 14'b10001101000001;
  assign mem[733] = 14'b00100001001001;
  assign mem[734] = 14'b10100000001111;
  assign mem[735] = 14'b00100111010111;
  assign mem[736] = 14'b10010100111101;
  assign mem[737] = 14'b00111011110000;
  assign mem[738] = 14'b10000111100010;
  assign mem[739] = 14'b10110010011011;
  assign mem[740] = 14'b10101010001000;
  assign mem[741] = 14'b01001010011010;
  assign mem[742] = 14'b10110000100111;
  assign mem[743] = 14'b01000000000001;
  assign mem[744] = 14'b00100101101110;
  assign mem[745] = 14'b01100101100000;
  assign mem[746] = 14'b10011011100001;
  assign mem[747] = 14'b10100100111010;
  assign mem[748] = 14'b00001100101000;
  assign mem[749] = 14'b00101110110111;
  assign mem[750] = 14'b00100001010010;
  assign mem[751] = 14'b01000010111110;
  assign mem[752] = 14'b10111100101110;
  assign mem[753] = 14'b01110100010101;
  assign mem[754] = 14'b01010000001100;
  assign mem[755] = 14'b01111011101011;
  assign mem[756] = 14'b00000011110101;
  assign mem[757] = 14'b01011101010110;
  assign mem[758] = 14'b01001100001010;
  assign mem[759] = 14'b01110001111100;
  assign mem[760] = 14'b01110110001000;
  assign mem[761] = 14'b10100100101011;
  assign mem[762] = 14'b10011011100000;
  assign mem[763] = 14'b10001101110011;
  assign mem[764] = 14'b00100001000001;
  assign mem[765] = 14'b00111010001001;
  assign mem[766] = 14'b10100000101101;
  assign mem[767] = 14'b10011100100110;
  assign mem[768] = 14'b10010101101010;
  assign mem[769] = 14'b10001011100110;
  assign mem[770] = 14'b10101101000010;
  assign mem[771] = 14'b10010100011010;
  assign mem[772] = 14'b00000100100110;
  assign mem[773] = 14'b01001001100111;
  assign mem[774] = 14'b00110100111111;
  assign mem[775] = 14'b00010101100001;
  assign mem[776] = 14'b10001101110000;
  assign mem[777] = 14'b10011111001101;
  assign mem[778] = 14'b01000111011001;
  assign mem[779] = 14'b10101010001010;
  assign mem[780] = 14'b10011010110101;
  assign mem[781] = 14'b01101100001011;
  assign mem[782] = 14'b00000000110101;
  assign mem[783] = 14'b01001000101101;
  assign mem[784] = 14'b00000110110111;
  assign mem[785] = 14'b10100000001101;
  assign mem[786] = 14'b01101101110100;
  assign mem[787] = 14'b10011111011111;
  assign mem[788] = 14'b10000010010111;
  assign mem[789] = 14'b00010001110101;
  assign mem[790] = 14'b00100111111100;
  assign mem[791] = 14'b01110110110001;
  assign mem[792] = 14'b01111111010110;
  assign mem[793] = 14'b10100110000110;
  assign mem[794] = 14'b10000111001000;
  assign mem[795] = 14'b10011001101000;
  assign mem[796] = 14'b01111100001111;
  assign mem[797] = 14'b10101111101101;
  assign mem[798] = 14'b00100001010011;
  assign mem[799] = 14'b01011010000101;
  assign mem[800] = 14'b10100001100111;
  assign mem[801] = 14'b10011000110101;
  assign mem[802] = 14'b00101010011110;
  assign mem[803] = 14'b00010110001011;
  assign mem[804] = 14'b01000110110011;
  assign mem[805] = 14'b00111100000100;
  assign mem[806] = 14'b00111111100010;
  assign mem[807] = 14'b01000011000101;
  assign mem[808] = 14'b10110110001001;
  assign mem[809] = 14'b10110100000101;
  assign mem[810] = 14'b10110001011001;
  assign mem[811] = 14'b01000011011001;
  assign mem[812] = 14'b01001100000101;
  assign mem[813] = 14'b10111110011010;
  assign mem[814] = 14'b00011001001011;
  assign mem[815] = 14'b10101010001100;
  assign mem[816] = 14'b10110011100001;
  assign mem[817] = 14'b10001010000001;
  assign mem[818] = 14'b00100101011001;
  assign mem[819] = 14'b00000000001111;
  assign mem[820] = 14'b10101001001110;
  assign mem[821] = 14'b01001110001011;
  assign mem[822] = 14'b00000000010001;
  assign mem[823] = 14'b00001000110101;
  assign mem[824] = 14'b01011100000011;
  assign mem[825] = 14'b10111110010001;
  assign mem[826] = 14'b10101100110010;
  assign mem[827] = 14'b10100010101100;
  assign mem[828] = 14'b10001010110101;
  assign mem[829] = 14'b00111110000110;
  assign mem[830] = 14'b10101011100101;
  assign mem[831] = 14'b01101111011010;
  assign mem[832] = 14'b01011011010000;
  assign mem[833] = 14'b10100011110010;
  assign mem[834] = 14'b10000010010010;
  assign mem[835] = 14'b01011110010011;
  assign mem[836] = 14'b01101100110100;
  assign mem[837] = 14'b00011000100110;
  assign mem[838] = 14'b10101010111000;
  assign mem[839] = 14'b00011111100100;
  assign mem[840] = 14'b00100110100001;
  assign mem[841] = 14'b01111111111111;
  assign mem[842] = 14'b00000110000000;
  assign mem[843] = 14'b00101001010010;
  assign mem[844] = 14'b00101010101001;
  assign mem[845] = 14'b01010100010111;
  assign mem[846] = 14'b00100001111111;
  assign mem[847] = 14'b10010010110100;
  assign mem[848] = 14'b10111011010011;
  assign mem[849] = 14'b01111101100011;
  assign mem[850] = 14'b01000100010111;
  assign mem[851] = 14'b01100111010011;
  assign mem[852] = 14'b01001110010010;
  assign mem[853] = 14'b10111000100100;
  assign mem[854] = 14'b10001110101011;
  assign mem[855] = 14'b10110010100011;
  assign mem[856] = 14'b00000001101000;
  assign mem[857] = 14'b01100011001100;
  assign mem[858] = 14'b10010110101011;
  assign mem[859] = 14'b01101001100101;
  assign mem[860] = 14'b10111101001110;
  assign mem[861] = 14'b01010111110001;
  assign mem[862] = 14'b10101010110111;
  assign mem[863] = 14'b00001000011101;
  assign mem[864] = 14'b00000010000111;
  assign mem[865] = 14'b00101111100001;
  assign mem[866] = 14'b01110000100000;
  assign mem[867] = 14'b01100101111110;
  assign mem[868] = 14'b01001111011101;
  assign mem[869] = 14'b10111101101000;
  assign mem[870] = 14'b00001101001010;
  assign mem[871] = 14'b01000000100001;
  assign mem[872] = 14'b01111000000101;
  assign mem[873] = 14'b10101101000111;
  assign mem[874] = 14'b10000011101010;
  assign mem[875] = 14'b00001111110000;
  assign mem[876] = 14'b00101010100101;
  assign mem[877] = 14'b10110111111100;
  assign mem[878] = 14'b01011110101010;
  assign mem[879] = 14'b00010001001101;
  assign mem[880] = 14'b00011110011110;
  assign mem[881] = 14'b10000011101000;
  assign mem[882] = 14'b01011000111000;
  assign mem[883] = 14'b01101011011100;
  assign mem[884] = 14'b10111011100101;
  assign mem[885] = 14'b10011101011111;
  assign mem[886] = 14'b01010011010111;
  assign mem[887] = 14'b00001110011111;
  assign mem[888] = 14'b00011011101010;
  assign mem[889] = 14'b00000100010001;
  assign mem[890] = 14'b10000010111001;
  assign mem[891] = 14'b00100011011111;
  assign mem[892] = 14'b01010001101001;
  assign mem[893] = 14'b10100000101011;
  assign mem[894] = 14'b00000001110100;
  assign mem[895] = 14'b10111000011111;
  assign mem[896] = 14'b00000001011011;
  assign mem[897] = 14'b10110110110011;
  assign mem[898] = 14'b00001011110101;
  assign mem[899] = 14'b00010100011000;
  assign mem[900] = 14'b01110101100100;
  assign mem[901] = 14'b01100100110011;
  assign mem[902] = 14'b01111101100000;
  assign mem[903] = 14'b01111111011010;
  assign mem[904] = 14'b01110100100000;
  assign mem[905] = 14'b01000001011111;
  assign mem[906] = 14'b00000100110101;
  assign mem[907] = 14'b00100100001110;
  assign mem[908] = 14'b00100011110100;
  assign mem[909] = 14'b10100010011001;
  assign mem[910] = 14'b10110101110111;
  assign mem[911] = 14'b10010100001001;
  assign mem[912] = 14'b10111111001110;
  assign mem[913] = 14'b10100101100010;
  assign mem[914] = 14'b10010101100001;
  assign mem[915] = 14'b01111011101000;
  assign mem[916] = 14'b10100010000000;
  assign mem[917] = 14'b10011010100001;
  assign mem[918] = 14'b10111111010100;
  assign mem[919] = 14'b01110000001011;
  assign mem[920] = 14'b00111101010100;
  assign mem[921] = 14'b00110001110100;
  assign mem[922] = 14'b00000101101111;
  assign mem[923] = 14'b00100000011101;
  assign mem[924] = 14'b00000101010000;
  assign mem[925] = 14'b01010100001000;
  assign mem[926] = 14'b01010111111111;
  assign mem[927] = 14'b10000110010100;
  assign mem[928] = 14'b01001000001101;
  assign mem[929] = 14'b00011011101111;
  assign mem[930] = 14'b10001010100010;
  assign mem[931] = 14'b00000111000011;
  assign mem[932] = 14'b01011111011100;
  assign mem[933] = 14'b00010100100101;
  assign mem[934] = 14'b01100001100110;
  assign mem[935] = 14'b10001001011011;
  assign mem[936] = 14'b01011100001000;
  assign mem[937] = 14'b01110001110011;
  assign mem[938] = 14'b00110000111100;
  assign mem[939] = 14'b10110100101100;
  assign mem[940] = 14'b01001101110001;
  assign mem[941] = 14'b10111110000001;
  assign mem[942] = 14'b01110011001011;
  assign mem[943] = 14'b00010101010110;
  assign mem[944] = 14'b10111101100010;
  assign mem[945] = 14'b10100101111011;
  assign mem[946] = 14'b00111011100001;
  assign mem[947] = 14'b01010000011101;
  assign mem[948] = 14'b01100010011100;
  assign mem[949] = 14'b00101001001110;
  assign mem[950] = 14'b01000001100101;
  assign mem[951] = 14'b00010110001010;
  assign mem[952] = 14'b10011101010001;
  assign mem[953] = 14'b01000000111100;
  assign mem[954] = 14'b10000010110101;
  assign mem[955] = 14'b10000111000100;
  assign mem[956] = 14'b10100011001101;
  assign mem[957] = 14'b00001101110010;
  assign mem[958] = 14'b01111111011110;
  assign mem[959] = 14'b10011110111101;
  assign mem[960] = 14'b10011000100011;
  assign mem[961] = 14'b10111110011111;
  assign mem[962] = 14'b00000111001011;
  assign mem[963] = 14'b00101110010110;
  assign mem[964] = 14'b00110001011110;
  assign mem[965] = 14'b00000110010101;
  assign mem[966] = 14'b01001110001000;
  assign mem[967] = 14'b10010001011111;
  assign mem[968] = 14'b01100100000100;
  assign mem[969] = 14'b10001100011010;
  assign mem[970] = 14'b00011000001111;
  assign mem[971] = 14'b01111111101111;
  assign mem[972] = 14'b00111000101110;
  assign mem[973] = 14'b10101000001110;
  assign mem[974] = 14'b10010000110001;
  assign mem[975] = 14'b00001010111100;
  assign mem[976] = 14'b10000101111101;
  assign mem[977] = 14'b10010100100100;
  assign mem[978] = 14'b01100111100110;
  assign mem[979] = 14'b10110010101101;
  assign mem[980] = 14'b10110101001011;
  assign mem[981] = 14'b01011011011010;
  assign mem[982] = 14'b00111101101110;
  assign mem[983] = 14'b01001010100111;
  assign mem[984] = 14'b10111010100101;
  assign mem[985] = 14'b00010110100110;
  assign mem[986] = 14'b01011110000010;
  assign mem[987] = 14'b00110100111010;
  assign mem[988] = 14'b10110011001110;
  assign mem[989] = 14'b01010010111110;
  assign mem[990] = 14'b01010101100100;
  assign mem[991] = 14'b00001000101001;
  assign mem[992] = 14'b10010100000010;
  assign mem[993] = 14'b00101000011010;
  assign mem[994] = 14'b00010110010111;
  assign mem[995] = 14'b00101010110101;
  assign mem[996] = 14'b00000111011001;
  assign mem[997] = 14'b10110001110111;
  assign mem[998] = 14'b01001010001001;
  assign mem[999] = 14'b00001101000100;
  assign mem[1000] = 14'b00111111011110;
  assign mem[1001] = 14'b10100110101010;
  assign mem[1002] = 14'b01111000101111;
  assign mem[1003] = 14'b10110111101000;
  assign mem[1004] = 14'b01010110011110;
  assign mem[1005] = 14'b00000100111000;
  assign mem[1006] = 14'b01000011010011;
  assign mem[1007] = 14'b01000011111111;
  assign mem[1008] = 14'b01011010000100;
  assign mem[1009] = 14'b10000111100111;
  assign mem[1010] = 14'b10000010111101;
  assign mem[1011] = 14'b01111111111011;
  assign mem[1012] = 14'b00000000000101;
  assign mem[1013] = 14'b01110011100011;
  assign mem[1014] = 14'b01000100001011;
  assign mem[1015] = 14'b00010010000000;
  assign mem[1016] = 14'b01010100101101;
  assign mem[1017] = 14'b01010001101111;
  assign mem[1018] = 14'b01100101001001;
  assign mem[1019] = 14'b00000110110100;
  assign mem[1020] = 14'b01110110001111;
  assign mem[1021] = 14'b10000110011011;
  assign mem[1022] = 14'b01100001010101;
  assign mem[1023] = 14'b10000000100110;

  always@(*)
  begin
    data_out_t <= mem[addr_f];
  end

  // Build output registers
  wire [13:0] data_out_reg [n_outreg:0];
  generate if (n_outreg > 0)
  begin
    for( i=n_outreg-1; i >= 1; i=i-1)
    begin: data_out_reg_stage
      mgc_generic_reg #(
        .width(14), 
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_data_out_reg (
        .d(data_out_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(data_out_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(14), 
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_data_out_reg_init (
      .d(data_out_t),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(data_out_reg[0])
    );
    assign data_out = data_out_reg[n_outreg-1];
  end
  else
  begin
    assign data_out = data_out_t;
  end
  endgenerate

endmodule



//------> ./rtl_stagemgc_rom_sync_regout_10_1024_62_1_0_0_1_0_1_0_0_0_1_60.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Sun Oct  6 01:48:34 2024
// ----------------------------------------------------------------------

// 
module stagemgc_rom_sync_regout_10_1024_62_1_0_0_1_0_1_0_0_0_1_60 (addr, data_out,
    clk, s_rst, a_rst, en
);
  input [9:0]addr ;
  output [61:0]data_out ;
  input clk ;
  input s_rst ;
  input a_rst ;
  input en ;


  // Constants for ROM dimensions
  parameter n_width    = 62;
  parameter n_size     = 1024;
  parameter n_numports = 1;
  parameter n_addr_w   = 10;
  parameter n_inreg    = 0;
  parameter n_outreg   = 1;
  wire [9:0] addr_f;

  // Build input address registers
  wire [9:0] addr_reg [n_inreg:0];
  genvar i;
  generate if (n_inreg > 0)
  begin
    for( i=n_inreg-1; i >= 1; i=i-1)
    begin: addr_reg_stage
      mgc_generic_reg #(
        .width(10), 
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_addr_reg (
        .d(addr_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(addr_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(10), 
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_addr_reg_init (
      .d(addr),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(addr_reg[0])
    );
    assign addr_f = addr_reg[n_inreg-1];
  end
  else
  begin
    assign addr_f = addr;
  end
  endgenerate

  // Declare storage for memory elements
  wire [61:0] mem [1023:0];

  // Declare output registers
  reg [61:0] data_out_t;

  // Initialize ROM contents
  assign mem[0] = 62'b00000000000000000000000000000000000000000000000000000000000000;
  assign mem[1] = 62'b11111111110000000000000000000000000000000000000000000000000000;
  assign mem[2] = 62'b11111111100110101000001001111001100110011111110011101111001101;
  assign mem[3] = 62'b11111111100110101000001001111001100110011111110011101111001101;
  assign mem[4] = 62'b11111111011000011111011110001010100110101011101010100101100011;
  assign mem[5] = 62'b11111111101101100100000110101111001111001100101000110101000110;
  assign mem[6] = 62'b11111111101101100100000110101111001111001100101000110101000110;
  assign mem[7] = 62'b11111111011000011111011110001010100110101011101010100101100011;
  assign mem[8] = 62'b11111111001000111110001011100000111100011010011010011000001011;
  assign mem[9] = 62'b11111111101111011000101001011111001111111101110101110010110000;
  assign mem[10] = 62'b11111111101010100110110110011000101001000011101010000110100011;
  assign mem[11] = 62'b11111111100001110001110011101100111001101011100110100011001000;
  assign mem[12] = 62'b11111111100001110001110011101100111001101011100110100011001000;
  assign mem[13] = 62'b11111111101010100110110110011000101001000011101010000110100011;
  assign mem[14] = 62'b11111111101111011000101001011111001111111101110101110010110000;
  assign mem[15] = 62'b11111111001000111110001011100000111100011010011010011000001011;
  assign mem[16] = 62'b11111110111001000101111010011010111100001010011011010000101100;
  assign mem[17] = 62'b11111111101111110110001000110110100011110100010010010100100110;
  assign mem[18] = 62'b11111111101000101111001000000001101011000101010001011101000001;
  assign mem[19] = 62'b11111111100100010011001111001100100101000010010001110111010110;
  assign mem[20] = 62'b11111111011110001010110101110100111000000001101111011000111011;
  assign mem[21] = 62'b11111111101100001110001011001011110001100000001011110110110001;
  assign mem[22] = 62'b11111111101110100111110100000101010110110001100010110111011010;
  assign mem[23] = 62'b11111111010010100101000000011000101110110101011001111100000110;
  assign mem[24] = 62'b11111111010010100101000000011000101110110101011001111100000110;
  assign mem[25] = 62'b11111111101110100111110100000101010110110001100010110111011010;
  assign mem[26] = 62'b11111111101100001110001011001011110001100000001011110110110001;
  assign mem[27] = 62'b11111111011110001010110101110100111000000001101111011000111011;
  assign mem[28] = 62'b11111111100100010011001111001100100101000010010001110111010110;
  assign mem[29] = 62'b11111111101000101111001000000001101011000101010001011101000001;
  assign mem[30] = 62'b11111111101111110110001000110110100011110100010010010100100110;
  assign mem[31] = 62'b11111110111001000101111010011010111100001010011011010000101100;
  assign mem[32] = 62'b11111110101001000111110110010111110001000011011101100000010100;
  assign mem[33] = 62'b11111111101111111101100010000111100011011110010110110101111110;
  assign mem[34] = 62'b11111111100111101101011101111100100010011010101010111110101111;
  assign mem[35] = 62'b11111111100101011111010110100100110100100011001110110010100000;
  assign mem[36] = 62'b11111111011011010111010001000000001001111000010101110011000000;
  assign mem[37] = 62'b11111111101100111011010111101011110100001111001100011101110011;
  assign mem[38] = 62'b11111111101110001000010010000100000100111101101000011011100101;
  assign mem[39] = 62'b11111111010101100011111001101001110101101010110001111111011101;
  assign mem[40] = 62'b11111111001111000110011111100101111011001000010101111100011011;
  assign mem[41] = 62'b11111111101111000010100111111011111011100100100011000011010111;
  assign mem[42] = 62'b11111111101011011100101000001101000101000110010110111000111110;
  assign mem[43] = 62'b11111111100000011100111000011110011001001000101111111111101110;
  assign mem[44] = 62'b11111111100011000011111111011111111100111000010111000000110101;
  assign mem[45] = 62'b11111111101001101100111110000001000111111100111000011101000001;
  assign mem[46] = 62'b11111111101111101001110101010101111111000010001010010100010111;
  assign mem[47] = 62'b11111111000010110010000001000001101110100011100110000100111010;
  assign mem[48] = 62'b11111111000010110010000001000001101110100011100110000100111010;
  assign mem[49] = 62'b11111111101111101001110101010101111111000010001010010100010111;
  assign mem[50] = 62'b11111111101001101100111110000001000111111100111000011101000001;
  assign mem[51] = 62'b11111111100011000011111111011111111100111000010111000000110101;
  assign mem[52] = 62'b11111111100000011100111000011110011001001000101111111111101110;
  assign mem[53] = 62'b11111111101011011100101000001101000101000110010110111000111110;
  assign mem[54] = 62'b11111111101111000010100111111011111011100100100011000011010111;
  assign mem[55] = 62'b11111111001111000110011111100101111011001000010101111100011011;
  assign mem[56] = 62'b11111111010101100011111001101001110101101010110001111111011101;
  assign mem[57] = 62'b11111111101110001000010010000100000100111101101000011011100101;
  assign mem[58] = 62'b11111111101100111011010111101011110100001111001100011101110011;
  assign mem[59] = 62'b11111111011011010111010001000000001001111000010101110011000000;
  assign mem[60] = 62'b11111111100101011111010110100100110100100011001110110010100000;
  assign mem[61] = 62'b11111111100111101101011101111100100010011010101010111110101111;
  assign mem[62] = 62'b11111111101111111101100010000111100011011110010110110101111110;
  assign mem[63] = 62'b11111110101001000111110110010111110001000011011101100000010100;
  assign mem[64] = 62'b11111110011001001000010101010111110111101000110110011001111110;
  assign mem[65] = 62'b11111111101111111111011000100001100000100001001100110100001101;
  assign mem[66] = 62'b11111111100111001011010000100000110111111011111111111110010110;
  assign mem[67] = 62'b11111111100110000100001011011101010101000111010010110011011111;
  assign mem[68] = 62'b11111111011001111011110111100101000011101010001110110110001010;
  assign mem[69] = 62'b11111111101101010000010011010011010001010011011100100100111010;
  assign mem[70] = 62'b11111111101101110110110001001110110110110011001100001000111100;
  assign mem[71] = 62'b11111111010111000010001000010100110000111110100100010110011111;
  assign mem[72] = 62'b11111111001100000010111000001001101010011111100100111101100011;
  assign mem[73] = 62'b11111111101111001110001111001110101100011001001110010110001001;
  assign mem[74] = 62'b11111111101011000010010000101001011000000101010000001000000000;
  assign mem[75] = 62'b11111111100001000111101011001101010100000110110100101100100011;
  assign mem[76] = 62'b11111111100010011011010000010101001100110111010001001011011111;
  assign mem[77] = 62'b11111111101010001010011010011110100000010001100010011110000010;
  assign mem[78] = 62'b11111111101111100001110110010011111010011100010100101110101001;
  assign mem[79] = 62'b11111111000101111000100001010001000100100010110011111111000110;
  assign mem[80] = 62'b11111110111111010101100100111001010110101010010111001100001110;
  assign mem[81] = 62'b11111111101111110000100110010001110000111000011001111111010011;
  assign mem[82] = 62'b11111111101001001110100010001001001001100100100110001111111011;
  assign mem[83] = 62'b11111111100011101011111111101000101001001000000101000010111001;
  assign mem[84] = 62'b11111111011111100010111010010011011011111110001001101010111010;
  assign mem[85] = 62'b11111111101011110101111100000010101100011011111001010100101010;
  assign mem[86] = 62'b11111111101110110101110100000011100111011010000100100101100011;
  assign mem[87] = 62'b11111111010001000100011101001001100010101100011111011001110111;
  assign mem[88] = 62'b11111111010100000100110101110010010100000101110110011000000001;
  assign mem[89] = 62'b11111111101110011000101000100011101100010010001110000100010010;
  assign mem[90] = 62'b11111111101100100101010100101100100001001101000001000111110101;
  assign mem[91] = 62'b11111111011100110001100110111010011001001100011100010001011110;
  assign mem[92] = 62'b11111111100100111001101100101010111011111000111110010111101001;
  assign mem[93] = 62'b11111111101000001110110000111000001011111111111001011101101110;
  assign mem[94] = 62'b11111111101111111010011100110110101101000000011000100000111010;
  assign mem[95] = 62'b11111110110010110101010010000010010010110011100001100111110110;
  assign mem[96] = 62'b11111110110010110101010010000010010010110011100001100111110110;
  assign mem[97] = 62'b11111111101111111010011100110110101101000000011000100000111010;
  assign mem[98] = 62'b11111111101000001110110000111000001011111111111001011101101110;
  assign mem[99] = 62'b11111111100100111001101100101010111011111000111110010111101001;
  assign mem[100] = 62'b11111111011100110001100110111010011001001100011100010001011110;
  assign mem[101] = 62'b11111111101100100101010100101100100001001101000001000111110101;
  assign mem[102] = 62'b11111111101110011000101000100011101100010010001110000100010010;
  assign mem[103] = 62'b11111111010100000100110101110010010100000101110110011000000001;
  assign mem[104] = 62'b11111111010001000100011101001001100010101100011111011001110111;
  assign mem[105] = 62'b11111111101110110101110100000011100111011010000100100101100011;
  assign mem[106] = 62'b11111111101011110101111100000010101100011011111001010100101010;
  assign mem[107] = 62'b11111111011111100010111010010011011011111110001001101010111010;
  assign mem[108] = 62'b11111111100011101011111111101000101001001000000101000010111001;
  assign mem[109] = 62'b11111111101001001110100010001001001001100100100110001111111011;
  assign mem[110] = 62'b11111111101111110000100110010001110000111000011001111111010011;
  assign mem[111] = 62'b11111110111111010101100100111001010110101010010111001100001110;
  assign mem[112] = 62'b11111111000101111000100001010001000100100010110011111111000110;
  assign mem[113] = 62'b11111111101111100001110110010011111010011100010100101110101001;
  assign mem[114] = 62'b11111111101010001010011010011110100000010001100010011110000010;
  assign mem[115] = 62'b11111111100010011011010000010101001100110111010001001011011111;
  assign mem[116] = 62'b11111111100001000111101011001101010100000110110100101100100011;
  assign mem[117] = 62'b11111111101011000010010000101001011000000101010000001000000000;
  assign mem[118] = 62'b11111111101111001110001111001110101100011001001110010110001001;
  assign mem[119] = 62'b11111111001100000010111000001001101010011111100100111101100011;
  assign mem[120] = 62'b11111111010111000010001000010100110000111110100100010110011111;
  assign mem[121] = 62'b11111111101101110110110001001110110110110011001100001000111100;
  assign mem[122] = 62'b11111111101101010000010011010011010001010011011100100100111010;
  assign mem[123] = 62'b11111111011001111011110111100101000011101010001110110110001010;
  assign mem[124] = 62'b11111111100110000100001011011101010101000111010010110011011111;
  assign mem[125] = 62'b11111111100111001011010000100000110111111011111111111110010110;
  assign mem[126] = 62'b11111111101111111111011000100001100000100001001100110100001101;
  assign mem[127] = 62'b11111110011001001000010101010111110111101000110110011001111110;
  assign mem[128] = 62'b11111110001001001000011101000111111100110111101100011110000100;
  assign mem[129] = 62'b11111111101111111111110110001000010110100110111001001011011011;
  assign mem[130] = 62'b11111111100110111001110100010001010100111010101010100010101111;
  assign mem[131] = 62'b11111111100110010110010001100100100101111100000111100000111101;
  assign mem[132] = 62'b11111111011001001101110010101001100011101111001001001111010111;
  assign mem[133] = 62'b11111111101101011010010110000101110011110010011110011010001011;
  assign mem[134] = 62'b11111111101101101101100101001001100010001110001010000010011011;
  assign mem[135] = 62'b11111111010111110000111010100100110001000111011100110011100111;
  assign mem[136] = 62'b11111111001010100000101010000000100101101100000000010001010001;
  assign mem[137] = 62'b11111111101111010011100110000000111011000010110010111100101101;
  assign mem[138] = 62'b11111111101010110100101011110010011110001000011101010100010001;
  assign mem[139] = 62'b11111111100001011100110100110101100011110111101101101101001001;
  assign mem[140] = 62'b11111111100010000110100111100110011001001100111110101101011001;
  assign mem[141] = 62'b11111111101010011000110000100100011011000000101111101011100010;
  assign mem[142] = 62'b11111111101111011101011001100110100011101000010010000001110111;
  assign mem[143] = 62'b11111111000111011011011101100111011110010100001011111100110001;
  assign mem[144] = 62'b11111110111100001101111000010111000111100111101100001011010101;
  assign mem[145] = 62'b11111111101111110011100001010111111101011011011010011001111011;
  assign mem[146] = 62'b11111111101000111110111100110010100011111011111001010000001101;
  assign mem[147] = 62'b11111111100011111111101101100101010011010001010101011011010100;
  assign mem[148] = 62'b11111111011110110111000001100101010010111011110111100011010110;
  assign mem[149] = 62'b11111111101100000010001100010000100110011100100101010101001001;
  assign mem[150] = 62'b11111111101110101110111101100011001000110111110000101101110100;
  assign mem[151] = 62'b11111111010001110100110100010000111111010011001101101100111110;
  assign mem[152] = 62'b11111111010011010101000001000011000010111000011000000101010010;
  assign mem[153] = 62'b11111111101110100000010111101110101011010011001101000100001101;
  assign mem[154] = 62'b11111111101100011001111000101100110100100010000111001110011011;
  assign mem[155] = 62'b11111111011101011110010111011101011011100001101110001110001001;
  assign mem[156] = 62'b11111111100100100110100100010010011011100110110000100100111001;
  assign mem[157] = 62'b11111111101000011111000100000000001111101110100010111010111111;
  assign mem[158] = 62'b11111111101111111000011100101011111100101111010101101100001001;
  assign mem[159] = 62'b11111110110101111101101101000000001010100110101010010000011001;
  assign mem[160] = 62'b11111110101111011001010110111001111001111110000010000011100000;
  assign mem[161] = 62'b11111111101111111100001001010101100101100011100111000110101101;
  assign mem[162] = 62'b11111111100111111110001110110011100011010101110001011101110001;
  assign mem[163] = 62'b11111111100101001100101000001010010010101000110101010110010110;
  assign mem[164] = 62'b11111111011100000100100100100111011000000000010001111011100111;
  assign mem[165] = 62'b11111111101100110000011111000011110011111111001111110001011100;
  assign mem[166] = 62'b11111111101110010000100110101001001011001010111100000101111110;
  assign mem[167] = 62'b11111111010100110100011110001001000010011110001110011101101010;
  assign mem[168] = 62'b11111111010000010011111011100000001110001101111111110110101110;
  assign mem[169] = 62'b11111111101110111100010111100010100011111001000111001111000010;
  assign mem[170] = 62'b11111111101011101001011010101001100111001101011001000011010010;
  assign mem[171] = 62'b11111111100000000111001111110010000111010011000011111010110111;
  assign mem[172] = 62'b11111111100011011000000101100010110001000001100101100111110011;
  assign mem[173] = 62'b11111111101001011101110111111011110100110001111101011101000010;
  assign mem[174] = 62'b11111111101111101101010111100101110001100101011101011101000001;
  assign mem[175] = 62'b11111111000001001110011111000011001110110110101111010101110111;
  assign mem[176] = 62'b11111111000100010101010111011010110001001010010011111001011010;
  assign mem[177] = 62'b11111111101111100101111111100100100100110010010000100110011011;
  assign mem[178] = 62'b11111111101001111011110100001111101111001010011010111110010100;
  assign mem[179] = 62'b11111111100010101111101101101100100101111110101111001111101010;
  assign mem[180] = 62'b11111111100000110010010111000001001101010111011000100110001111;
  assign mem[181] = 62'b11111111101011001111100100110100111110111101010101011100010010;
  assign mem[182] = 62'b11111111101111001000100101001011110111011101100011101011011010;
  assign mem[183] = 62'b11111111001101100100110100111111100101010001010100001100010001;
  assign mem[184] = 62'b11111111010110010011000111110111011101001111110010011111000110;
  assign mem[185] = 62'b11111111101101111111101010111001100010001011011011111000101011;
  assign mem[186] = 62'b11111111101101000101111110011101110100001111100011010111011100;
  assign mem[187] = 62'b11111111011010101001101100100000101011011011010011111111001010;
  assign mem[188] = 62'b11111111100101110001110111101110111110011001010000000110001100;
  assign mem[189] = 62'b11111111100111011100011110011101011111000000110111001001100001;
  assign mem[190] = 62'b11111111101111111110100111001011101111111111101111011101011101;
  assign mem[191] = 62'b11111110100010110110000110010101110101100101000101010111001101;
  assign mem[192] = 62'b11111110100010110110000110010101110101100101000101010111001101;
  assign mem[193] = 62'b11111111101111111110100111001011101111111111101111011101011101;
  assign mem[194] = 62'b11111111100111011100011110011101011111000000110111001001100001;
  assign mem[195] = 62'b11111111100101110001110111101110111110011001010000000110001100;
  assign mem[196] = 62'b11111111011010101001101100100000101011011011010011111111001010;
  assign mem[197] = 62'b11111111101101000101111110011101110100001111100011010111011100;
  assign mem[198] = 62'b11111111101101111111101010111001100010001011011011111000101011;
  assign mem[199] = 62'b11111111010110010011000111110111011101001111110010011111000110;
  assign mem[200] = 62'b11111111001101100100110100111111100101010001010100001100010001;
  assign mem[201] = 62'b11111111101111001000100101001011110111011101100011101011011010;
  assign mem[202] = 62'b11111111101011001111100100110100111110111101010101011100010010;
  assign mem[203] = 62'b11111111100000110010010111000001001101010111011000100110001111;
  assign mem[204] = 62'b11111111100010101111101101101100100101111110101111001111101010;
  assign mem[205] = 62'b11111111101001111011110100001111101111001010011010111110010100;
  assign mem[206] = 62'b11111111101111100101111111100100100100110010010000100110011011;
  assign mem[207] = 62'b11111111000100010101010111011010110001001010010011111001011010;
  assign mem[208] = 62'b11111111000001001110011111000011001110110110101111010101110111;
  assign mem[209] = 62'b11111111101111101101010111100101110001100101011101011101000001;
  assign mem[210] = 62'b11111111101001011101110111111011110100110001111101011101000010;
  assign mem[211] = 62'b11111111100011011000000101100010110001000001100101100111110011;
  assign mem[212] = 62'b11111111100000000111001111110010000111010011000011111010110111;
  assign mem[213] = 62'b11111111101011101001011010101001100111001101011001000011010010;
  assign mem[214] = 62'b11111111101110111100010111100010100011111001000111001111000010;
  assign mem[215] = 62'b11111111010000010011111011100000001110001101111111110110101110;
  assign mem[216] = 62'b11111111010100110100011110001001000010011110001110011101101010;
  assign mem[217] = 62'b11111111101110010000100110101001001011001010111100000101111110;
  assign mem[218] = 62'b11111111101100110000011111000011110011111111001111110001011100;
  assign mem[219] = 62'b11111111011100000100100100100111011000000000010001111011100111;
  assign mem[220] = 62'b11111111100101001100101000001010010010101000110101010110010110;
  assign mem[221] = 62'b11111111100111111110001110110011100011010101110001011101110001;
  assign mem[222] = 62'b11111111101111111100001001010101100101100011100111000110101101;
  assign mem[223] = 62'b11111110101111011001010110111001111001111110000010000011100000;
  assign mem[224] = 62'b11111110110101111101101101000000001010100110101010010000011001;
  assign mem[225] = 62'b11111111101111111000011100101011111100101111010101101100001001;
  assign mem[226] = 62'b11111111101000011111000100000000001111101110100010111010111111;
  assign mem[227] = 62'b11111111100100100110100100010010011011100110110000100100111001;
  assign mem[228] = 62'b11111111011101011110010111011101011011100001101110001110001001;
  assign mem[229] = 62'b11111111101100011001111000101100110100100010000111001110011011;
  assign mem[230] = 62'b11111111101110100000010111101110101011010011001101000100001101;
  assign mem[231] = 62'b11111111010011010101000001000011000010111000011000000101010010;
  assign mem[232] = 62'b11111111010001110100110100010000111111010011001101101100111110;
  assign mem[233] = 62'b11111111101110101110111101100011001000110111110000101101110100;
  assign mem[234] = 62'b11111111101100000010001100010000100110011100100101010101001001;
  assign mem[235] = 62'b11111111011110110111000001100101010010111011110111100011010110;
  assign mem[236] = 62'b11111111100011111111101101100101010011010001010101011011010100;
  assign mem[237] = 62'b11111111101000111110111100110010100011111011111001010000001101;
  assign mem[238] = 62'b11111111101111110011100001010111111101011011011010011001111011;
  assign mem[239] = 62'b11111110111100001101111000010111000111100111101100001011010101;
  assign mem[240] = 62'b11111111000111011011011101100111011110010100001011111100110001;
  assign mem[241] = 62'b11111111101111011101011001100110100011101000010010000001110111;
  assign mem[242] = 62'b11111111101010011000110000100100011011000000101111101011100010;
  assign mem[243] = 62'b11111111100010000110100111100110011001001100111110101101011001;
  assign mem[244] = 62'b11111111100001011100110100110101100011110111101101101101001001;
  assign mem[245] = 62'b11111111101010110100101011110010011110001000011101010100010001;
  assign mem[246] = 62'b11111111101111010011100110000000111011000010110010111100101101;
  assign mem[247] = 62'b11111111001010100000101010000000100101101100000000010001010001;
  assign mem[248] = 62'b11111111010111110000111010100100110001000111011100110011100111;
  assign mem[249] = 62'b11111111101101101101100101001001100010001110001010000010011011;
  assign mem[250] = 62'b11111111101101011010010110000101110011110010011110011010001011;
  assign mem[251] = 62'b11111111011001001101110010101001100011101111001001001111010111;
  assign mem[252] = 62'b11111111100110010110010001100100100101111100000111100000111101;
  assign mem[253] = 62'b11111111100110111001110100010001010100111010101010100010101111;
  assign mem[254] = 62'b11111111101111111111110110001000010110100110111001001011011011;
  assign mem[255] = 62'b11111110001001001000011101000111111100110111101100011110000100;
  assign mem[256] = 62'b11111101111001001000011111000011111110011001110000000001110001;
  assign mem[257] = 62'b11111111101111111111111101100010000101100011101000101010010010;
  assign mem[258] = 62'b11111111100110110001000000110101110011110000011000001001110101;
  assign mem[259] = 62'b11111111100110011111001111011110000100100100011010111100010000;
  assign mem[260] = 62'b11111111011000110110101010010100101110110010001010010010110000;
  assign mem[261] = 62'b11111111101101011111010000101100000010101110001110110011111001;
  assign mem[262] = 62'b11111111101101101000111000001110101001011001101000100110001000;
  assign mem[263] = 62'b11111111011000001000001110001110110000010011101010101011000100;
  assign mem[264] = 62'b11111111001001101111011100101111110010110111000100001101100110;
  assign mem[265] = 62'b11111111101111010110001010001010110001011110001001111010000100;
  assign mem[266] = 62'b11111111101010101101110011001001011001000101101100000011010100;
  assign mem[267] = 62'b11111111100001100111010101101000001001111100101011100110111000;
  assign mem[268] = 62'b11111111100001111100001111000010001011101111001000011000011011;
  assign mem[269] = 62'b11111111101010011111110101100001010010100111111110011010011101;
  assign mem[270] = 62'b11111111101111011011000011111101111101111101011011101110110111;
  assign mem[271] = 62'b11111111001000001100110110011011101000100111000110010011000110;
  assign mem[272] = 62'b11111110111010101001111011011100100100010010010101110000000011;
  assign mem[273] = 62'b11111111101111110100110111100100010100001000100000101110000100;
  assign mem[274] = 62'b11111111101000110111000100010100110011000101101001100011001100;
  assign mem[275] = 62'b11111111100100001001011111111100010111100011100110101110110001;
  assign mem[276] = 62'b11111111011110100000111110000011101010111110000101000100010100;
  assign mem[277] = 62'b11111111101100001000001101111000111111101010010111000110110000;
  assign mem[278] = 62'b11111111101110101011011011001011101000111001111010100010001110;
  assign mem[279] = 62'b11111111010010001100111011101110101011110000111011101101110001;
  assign mem[280] = 62'b11111111010010111101000010001011011010111011000000001110000111;
  assign mem[281] = 62'b11111111101110100100001000010000110110000111011111011111110010;
  assign mem[282] = 62'b11111111101100010100000100001000000001001010110110100100000111;
  assign mem[283] = 62'b11111111011101110100101000111100010100100000011100110001011000;
  assign mem[284] = 62'b11111111100100011100111011010100011011100110000111001101000111;
  assign mem[285] = 62'b11111111101000100111000111111010011010010011011101010010101010;
  assign mem[286] = 62'b11111111101111110111010101001110011111111100011111010001010110;
  assign mem[287] = 62'b11111110110111100001110101100001101010010111010101101100100001;
  assign mem[288] = 62'b11111110101100010000101000110100010010110000001101011111100011;
  assign mem[289] = 62'b11111111101111111100111000001100001111100011010101011101011100;
  assign mem[290] = 62'b11111111100111110101111000001101101100110000110011110110110010;
  assign mem[291] = 62'b11111111100101010110000001000000111000100101110101000100110111;
  assign mem[292] = 62'b11111111011011101101111100111100100011000001001011110100000001;
  assign mem[293] = 62'b11111111101100110101111101100110001001100010110011001011110110;
  assign mem[294] = 62'b11111111101110001100011110101011101000011100001100111000100101;
  assign mem[295] = 62'b11111111010101001100001101100010000000101011110011110000100100;
  assign mem[296] = 62'b11111111001111110111001101110000011010110111111110110111111001;
  assign mem[297] = 62'b11111111101110111111100010001000001100000010111001010111101100;
  assign mem[298] = 62'b11111111101011100011000011100011010010011101010000010011101001;
  assign mem[299] = 62'b11111111100000010010000101011000100110101011100010001000011010;
  assign mem[300] = 62'b11111111100011001110000100000000001101000011001000111001010111;
  assign mem[301] = 62'b11111111101001100101011100111100101110110110000000110100100010;
  assign mem[302] = 62'b11111111101111101011101000111010001110010001101100111110111011;
  assign mem[303] = 62'b11111111000010000000010001011011010100111011000111101111001111;
  assign mem[304] = 62'b11111111000011100011101101101110110000110011011000110100010100;
  assign mem[305] = 62'b11111111101111100111111100111001010101101011011011001011001000;
  assign mem[306] = 62'b11111111101001110100011011000111110101111010101000000011010101;
  assign mem[307] = 62'b11111111100010111001111000000011100011111010001110101000010111;
  assign mem[308] = 62'b11111111100000100111101001000001110100000101111100010111100001;
  assign mem[309] = 62'b11111111101011010110001000100111111110100100100001010000000101;
  assign mem[310] = 62'b11111111101111000101101000111101010011111101110010000001011101;
  assign mem[311] = 62'b11111111001110010101101100101000011110000100000001101000011011;
  assign mem[312] = 62'b11111111010101111011100010011100110111100111101010011010010011;
  assign mem[313] = 62'b11111111101110000100000000110011001010001010011000000010101100;
  assign mem[314] = 62'b11111111101101000000101101010011111110101100101011110110010010;
  assign mem[315] = 62'b11111111011011000000100000110101101100011111110100000000001001;
  assign mem[316] = 62'b11111111100101101000101000110100101010010111010111001001010000;
  assign mem[317] = 62'b11111111100111100101000000000001010111010011110101010111100101;
  assign mem[318] = 62'b11111111101111111110000111000111011010110110111000000111011111;
  assign mem[319] = 62'b11111110100101111111000000000011010010100100001100110101000011;
  assign mem[320] = 62'b11111110011111011010010011011100110001110100011100111100000001;
  assign mem[321] = 62'b11111111101111111111000010010100011101111100011101001111111000;
  assign mem[322] = 62'b11111111100111010011111001010010001101101010001101001010001101;
  assign mem[323] = 62'b11111111100101111011000011010010010101100000110111000001110100;
  assign mem[324] = 62'b11111111011010010010110100000100100111110111101010000111100101;
  assign mem[325] = 62'b11111111101101001011001011001000100000111000001110111110011111;
  assign mem[326] = 62'b11111111101101111011010000010111110111110111100100011111011010;
  assign mem[327] = 62'b11111111010110101010101001110101111101110001110111111000010111;
  assign mem[328] = 62'b11111111001100110011111000110010110011000100101011001010000110;
  assign mem[329] = 62'b11111111101111001011011100100111001001000010001001101010011101;
  assign mem[330] = 62'b11111111101011001000111100110101000111000000000001001110110100;
  assign mem[331] = 62'b11111111100000111101000010011010111011001010101000111001111110;
  assign mem[332] = 62'b11111111100010100101100000011100100111011000101001110010101000;
  assign mem[333] = 62'b11111111101010000011001001010111101010101110101111100100110111;
  assign mem[334] = 62'b11111111101111100011111101010111111111101011100100000111011011;
  assign mem[335] = 62'b11111111000101000110111101111110000101100101111100010111110010;
  assign mem[336] = 62'b11111111000000011100101010000001000111101110101000001100011101;
  assign mem[337] = 62'b11111111101111101111000001011000010111111001000100000110000110;
  assign mem[338] = 62'b11111111101001010110001110111111100100100011100110110111010111;
  assign mem[339] = 62'b11111111100011100010000100000110000101110111111110101100100010;
  assign mem[340] = 62'b11111111011111111000101111011001001011111001110001001000010000;
  assign mem[341] = 62'b11111111101011101111101101011111000100100100111000000011101010;
  assign mem[342] = 62'b11111111101110111001001000001011100010010110101001110110111100;
  assign mem[343] = 62'b11111111010000101100001101100111001111110110111101101110010000;
  assign mem[344] = 62'b11111111010100011100101011100010100101010101110001000001010100;
  assign mem[345] = 62'b11111111101110010100101001111100000100011100101001111111111100;
  assign mem[346] = 62'b11111111101100101010111100000101101001101000001011100100000000;
  assign mem[347] = 62'b11111111011100011011000111111101001001100101110000000000001011;
  assign mem[348] = 62'b11111111100101000011001100000010011111010110011010000010011011;
  assign mem[349] = 62'b11111111101000000110100001101100110011101101010111101011001100;
  assign mem[350] = 62'b11111111101111111011010101100011101100101101100111001111000100;
  assign mem[351] = 62'b11111110110001010001000000000100110100110101110000100110110011;
  assign mem[352] = 62'b11111110110100011001100001000101111001001001110010000010010110;
  assign mem[353] = 62'b11111111101111111001011111001110101111001011100011100101000000;
  assign mem[354] = 62'b11111111101000010110111100010100011010111010010101100011001100;
  assign mem[355] = 62'b11111111100100110000001010000101000101111011000000000000000100;
  assign mem[356] = 62'b11111111011101001000000001011011101000111010011101101101011011;
  assign mem[357] = 62'b11111111101100011111101000111001010010001000110011110011110011;
  assign mem[358] = 62'b11111111101110011100100010011111011011011010101001011101000100;
  assign mem[359] = 62'b11111111010011101100111100111011111010000001000001010010110111;
  assign mem[360] = 62'b11111111010001011100101010000011010111011101100101000101110111;
  assign mem[361] = 62'b11111111101110110010011011001011010011110000111011111110000100;
  assign mem[362] = 62'b11111111101011111100000110010011100001010100110111011111011101;
  assign mem[363] = 62'b11111111011111001101000000010110010110001111111101000001100111;
  assign mem[364] = 62'b11111111100011110101111000001000111000110001011000001101000100;
  assign mem[365] = 62'b11111111101001000110110001011001101111110101001001110110100010;
  assign mem[366] = 62'b11111111101111110010000110010001101100111111101011011100100001;
  assign mem[367] = 62'b11111110111101110001110000111011001011101011101001111111001001;
  assign mem[368] = 62'b11111111000110101010000001001100000100111101100100101010110010;
  assign mem[369] = 62'b11111111101111011111101010011000101001111001100011110101101110;
  assign mem[370] = 62'b11111111101010010001100111100011001000000100011001101011001000;
  assign mem[371] = 62'b11111111100010010000111101010111111011100110001010110000011111;
  assign mem[372] = 62'b11111111100001010010010001010110101111001100110110110011101011;
  assign mem[373] = 62'b11111111101010111011100000010010110100001111000001010001110100;
  assign mem[374] = 62'b11111111101111010000111101000010000101111111111001001011011101;
  assign mem[375] = 62'b11111111001011010001110011001011101111001111010110011100100010;
  assign mem[376] = 62'b11111111010111011001100011010000001111001001000001100011110110;
  assign mem[377] = 62'b11111111101101110010001101011111001011010000010000001001100000;
  assign mem[378] = 62'b11111111101101010101010110111101010010111010010011111010110001;
  assign mem[379] = 62'b11111111011001100100110111000101100001010000011011110111111111;
  assign mem[380] = 62'b11111111100110001101010000001110100011000111000001101111101001;
  assign mem[381] = 62'b11111111100111000010100100001010110011000101110110110101111010;
  assign mem[382] = 62'b11111111101111111111101001110010110100010010110101000110100001;
  assign mem[383] = 62'b11111110010010110110010011011010111011111000110000111011111101;
  assign mem[384] = 62'b11111110010010110110010011011010111011111000110000111011111101;
  assign mem[385] = 62'b11111111101111111111101001110010110100010010110101000110100001;
  assign mem[386] = 62'b11111111100111000010100100001010110011000101110110110101111010;
  assign mem[387] = 62'b11111111100110001101010000001110100011000111000001101111101001;
  assign mem[388] = 62'b11111111011001100100110111000101100001010000011011110111111111;
  assign mem[389] = 62'b11111111101101010101010110111101010010111010010011111010110001;
  assign mem[390] = 62'b11111111101101110010001101011111001011010000010000001001100000;
  assign mem[391] = 62'b11111111010111011001100011010000001111001001000001100011110110;
  assign mem[392] = 62'b11111111001011010001110011001011101111001111010110011100100010;
  assign mem[393] = 62'b11111111101111010000111101000010000101111111111001001011011101;
  assign mem[394] = 62'b11111111101010111011100000010010110100001111000001010001110100;
  assign mem[395] = 62'b11111111100001010010010001010110101111001100110110110011101011;
  assign mem[396] = 62'b11111111100010010000111101010111111011100110001010110000011111;
  assign mem[397] = 62'b11111111101010010001100111100011001000000100011001101011001000;
  assign mem[398] = 62'b11111111101111011111101010011000101001111001100011110101101110;
  assign mem[399] = 62'b11111111000110101010000001001100000100111101100100101010110010;
  assign mem[400] = 62'b11111110111101110001110000111011001011101011101001111111001001;
  assign mem[401] = 62'b11111111101111110010000110010001101100111111101011011100100001;
  assign mem[402] = 62'b11111111101001000110110001011001101111110101001001110110100010;
  assign mem[403] = 62'b11111111100011110101111000001000111000110001011000001101000100;
  assign mem[404] = 62'b11111111011111001101000000010110010110001111111101000001100111;
  assign mem[405] = 62'b11111111101011111100000110010011100001010100110111011111011101;
  assign mem[406] = 62'b11111111101110110010011011001011010011110000111011111110000100;
  assign mem[407] = 62'b11111111010001011100101010000011010111011101100101000101110111;
  assign mem[408] = 62'b11111111010011101100111100111011111010000001000001010010110111;
  assign mem[409] = 62'b11111111101110011100100010011111011011011010101001011101000100;
  assign mem[410] = 62'b11111111101100011111101000111001010010001000110011110011110011;
  assign mem[411] = 62'b11111111011101001000000001011011101000111010011101101101011011;
  assign mem[412] = 62'b11111111100100110000001010000101000101111011000000000000000100;
  assign mem[413] = 62'b11111111101000010110111100010100011010111010010101100011001100;
  assign mem[414] = 62'b11111111101111111001011111001110101111001011100011100101000000;
  assign mem[415] = 62'b11111110110100011001100001000101111001001001110010000010010110;
  assign mem[416] = 62'b11111110110001010001000000000100110100110101110000100110110011;
  assign mem[417] = 62'b11111111101111111011010101100011101100101101100111001111000100;
  assign mem[418] = 62'b11111111101000000110100001101100110011101101010111101011001100;
  assign mem[419] = 62'b11111111100101000011001100000010011111010110011010000010011011;
  assign mem[420] = 62'b11111111011100011011000111111101001001100101110000000000001011;
  assign mem[421] = 62'b11111111101100101010111100000101101001101000001011100100000000;
  assign mem[422] = 62'b11111111101110010100101001111100000100011100101001111111111100;
  assign mem[423] = 62'b11111111010100011100101011100010100101010101110001000001010100;
  assign mem[424] = 62'b11111111010000101100001101100111001111110110111101101110010000;
  assign mem[425] = 62'b11111111101110111001001000001011100010010110101001110110111100;
  assign mem[426] = 62'b11111111101011101111101101011111000100100100111000000011101010;
  assign mem[427] = 62'b11111111011111111000101111011001001011111001110001001000010000;
  assign mem[428] = 62'b11111111100011100010000100000110000101110111111110101100100010;
  assign mem[429] = 62'b11111111101001010110001110111111100100100011100110110111010111;
  assign mem[430] = 62'b11111111101111101111000001011000010111111001000100000110000110;
  assign mem[431] = 62'b11111111000000011100101010000001000111101110101000001100011101;
  assign mem[432] = 62'b11111111000101000110111101111110000101100101111100010111110010;
  assign mem[433] = 62'b11111111101111100011111101010111111111101011100100000111011011;
  assign mem[434] = 62'b11111111101010000011001001010111101010101110101111100100110111;
  assign mem[435] = 62'b11111111100010100101100000011100100111011000101001110010101000;
  assign mem[436] = 62'b11111111100000111101000010011010111011001010101000111001111110;
  assign mem[437] = 62'b11111111101011001000111100110101000111000000000001001110110100;
  assign mem[438] = 62'b11111111101111001011011100100111001001000010001001101010011101;
  assign mem[439] = 62'b11111111001100110011111000110010110011000100101011001010000110;
  assign mem[440] = 62'b11111111010110101010101001110101111101110001110111111000010111;
  assign mem[441] = 62'b11111111101101111011010000010111110111110111100100011111011010;
  assign mem[442] = 62'b11111111101101001011001011001000100000111000001110111110011111;
  assign mem[443] = 62'b11111111011010010010110100000100100111110111101010000111100101;
  assign mem[444] = 62'b11111111100101111011000011010010010101100000110111000001110100;
  assign mem[445] = 62'b11111111100111010011111001010010001101101010001101001010001101;
  assign mem[446] = 62'b11111111101111111111000010010100011101111100011101001111111000;
  assign mem[447] = 62'b11111110011111011010010011011100110001110100011100111100000001;
  assign mem[448] = 62'b11111110100101111111000000000011010010100100001100110101000011;
  assign mem[449] = 62'b11111111101111111110000111000111011010110110111000000111011111;
  assign mem[450] = 62'b11111111100111100101000000000001010111010011110101010111100101;
  assign mem[451] = 62'b11111111100101101000101000110100101010010111010111001001010000;
  assign mem[452] = 62'b11111111011011000000100000110101101100011111110100000000001001;
  assign mem[453] = 62'b11111111101101000000101101010011111110101100101011110110010010;
  assign mem[454] = 62'b11111111101110000100000000110011001010001010011000000010101100;
  assign mem[455] = 62'b11111111010101111011100010011100110111100111101010011010010011;
  assign mem[456] = 62'b11111111001110010101101100101000011110000100000001101000011011;
  assign mem[457] = 62'b11111111101111000101101000111101010011111101110010000001011101;
  assign mem[458] = 62'b11111111101011010110001000100111111110100100100001010000000101;
  assign mem[459] = 62'b11111111100000100111101001000001110100000101111100010111100001;
  assign mem[460] = 62'b11111111100010111001111000000011100011111010001110101000010111;
  assign mem[461] = 62'b11111111101001110100011011000111110101111010101000000011010101;
  assign mem[462] = 62'b11111111101111100111111100111001010101101011011011001011001000;
  assign mem[463] = 62'b11111111000011100011101101101110110000110011011000110100010100;
  assign mem[464] = 62'b11111111000010000000010001011011010100111011000111101111001111;
  assign mem[465] = 62'b11111111101111101011101000111010001110010001101100111110111011;
  assign mem[466] = 62'b11111111101001100101011100111100101110110110000000110100100010;
  assign mem[467] = 62'b11111111100011001110000100000000001101000011001000111001010111;
  assign mem[468] = 62'b11111111100000010010000101011000100110101011100010001000011010;
  assign mem[469] = 62'b11111111101011100011000011100011010010011101010000010011101001;
  assign mem[470] = 62'b11111111101110111111100010001000001100000010111001010111101100;
  assign mem[471] = 62'b11111111001111110111001101110000011010110111111110110111111001;
  assign mem[472] = 62'b11111111010101001100001101100010000000101011110011110000100100;
  assign mem[473] = 62'b11111111101110001100011110101011101000011100001100111000100101;
  assign mem[474] = 62'b11111111101100110101111101100110001001100010110011001011110110;
  assign mem[475] = 62'b11111111011011101101111100111100100011000001001011110100000001;
  assign mem[476] = 62'b11111111100101010110000001000000111000100101110101000100110111;
  assign mem[477] = 62'b11111111100111110101111000001101101100110000110011110110110010;
  assign mem[478] = 62'b11111111101111111100111000001100001111100011010101011101011100;
  assign mem[479] = 62'b11111110101100010000101000110100010010110000001101011111100011;
  assign mem[480] = 62'b11111110110111100001110101100001101010010111010101101100100001;
  assign mem[481] = 62'b11111111101111110111010101001110011111111100011111010001010110;
  assign mem[482] = 62'b11111111101000100111000111111010011010010011011101010010101010;
  assign mem[483] = 62'b11111111100100011100111011010100011011100110000111001101000111;
  assign mem[484] = 62'b11111111011101110100101000111100010100100000011100110001011000;
  assign mem[485] = 62'b11111111101100010100000100001000000001001010110110100100000111;
  assign mem[486] = 62'b11111111101110100100001000010000110110000111011111011111110010;
  assign mem[487] = 62'b11111111010010111101000010001011011010111011000000001110000111;
  assign mem[488] = 62'b11111111010010001100111011101110101011110000111011101101110001;
  assign mem[489] = 62'b11111111101110101011011011001011101000111001111010100010001110;
  assign mem[490] = 62'b11111111101100001000001101111000111111101010010111000110110000;
  assign mem[491] = 62'b11111111011110100000111110000011101010111110000101000100010100;
  assign mem[492] = 62'b11111111100100001001011111111100010111100011100110101110110001;
  assign mem[493] = 62'b11111111101000110111000100010100110011000101101001100011001100;
  assign mem[494] = 62'b11111111101111110100110111100100010100001000100000101110000100;
  assign mem[495] = 62'b11111110111010101001111011011100100100010010010101110000000011;
  assign mem[496] = 62'b11111111001000001100110110011011101000100111000110010011000110;
  assign mem[497] = 62'b11111111101111011011000011111101111101111101011011101110110111;
  assign mem[498] = 62'b11111111101010011111110101100001010010100111111110011010011101;
  assign mem[499] = 62'b11111111100001111100001111000010001011101111001000011000011011;
  assign mem[500] = 62'b11111111100001100111010101101000001001111100101011100110111000;
  assign mem[501] = 62'b11111111101010101101110011001001011001000101101100000011010100;
  assign mem[502] = 62'b11111111101111010110001010001010110001011110001001111010000100;
  assign mem[503] = 62'b11111111001001101111011100101111110010110111000100001101100110;
  assign mem[504] = 62'b11111111011000001000001110001110110000010011101010101011000100;
  assign mem[505] = 62'b11111111101101101000111000001110101001011001101000100110001000;
  assign mem[506] = 62'b11111111101101011111010000101100000010101110001110110011111001;
  assign mem[507] = 62'b11111111011000110110101010010100101110110010001010010010110000;
  assign mem[508] = 62'b11111111100110011111001111011110000100100100011010111100010000;
  assign mem[509] = 62'b11111111100110110001000000110101110011110000011000001001110101;
  assign mem[510] = 62'b11111111101111111111111101100010000101100011101000101010010010;
  assign mem[511] = 62'b11111101111001001000011111000011111110011001110000000001110001;
  assign mem[512] = 62'b11111101101001001000011111100010111110110011001010010010111010;
  assign mem[513] = 62'b11111111101111111111111111011000100001011000100001110100000010;
  assign mem[514] = 62'b11111111100110101100100101110011101101001011111110001010011100;
  assign mem[515] = 62'b11111111100110100011101101000111101010101000011001110001110001;
  assign mem[516] = 62'b11111111011000101011000100101110000110110101011110110101000100;
  assign mem[517] = 62'b11111111101101100001101100010010000100010001011010010001001111;
  assign mem[518] = 62'b11111111101101100110100000000011011101100010110011110101000110;
  assign mem[519] = 62'b11111111011000010011110110101010101010111100111001000000111111;
  assign mem[520] = 62'b11111111001001010110110100100111101001101101100010101011111010;
  assign mem[521] = 62'b11111111101111010111011010011011101101010000110110100001011101;
  assign mem[522] = 62'b11111111101010101010010101010001111010001011001011100110001110;
  assign mem[523] = 62'b11111111100001101100100101000000010111000100110111001110111111;
  assign mem[524] = 62'b11111111100001110111000001101101100100110111000100100001110010;
  assign mem[525] = 62'b11111111101010100011010110011101101110010101000101101011010010;
  assign mem[526] = 62'b11111111101111011001110111010101010110100010000011110011101110;
  assign mem[527] = 62'b11111111001000100101100001011100100111110001000001100000000100;
  assign mem[528] = 62'b11111110111001110111111011011011101011001001001010100001011100;
  assign mem[529] = 62'b11111111101111110101100000110100101101101001110101110010011110;
  assign mem[530] = 62'b11111111101000110011000110101001110101000110000100011001010101;
  assign mem[531] = 62'b11111111100100001110010111111101011011001010100100001110000000;
  assign mem[532] = 62'b11111111011110010101111010100001101101001111001101100000100101;
  assign mem[533] = 62'b11111111101100001011001101000101001001001100011110001111110001;
  assign mem[534] = 62'b11111111101110101001101000001110010011111001100101100000000000;
  assign mem[535] = 62'b11111111010010011000111110011010011001010101010101010010111010;
  assign mem[536] = 62'b11111111010010110001000001101001001110100101010100010100100000;
  assign mem[537] = 62'b11111111101110100101111110110000110110000000010110101100110000;
  assign mem[538] = 62'b11111111101100010001001000001100110001010000011100000000000100;
  assign mem[539] = 62'b11111111011101111111101111111101100110101010010100000111011110;
  assign mem[540] = 62'b11111111100100011000000101101001101001001010110011001010100010;
  assign mem[541] = 62'b11111111101000101011001000011100011110110111100001110110001000;
  assign mem[542] = 62'b11111111101111110110101111101001110101000101000101001110001100;
  assign mem[543] = 62'b11111110111000010011111000011100010010110000010011000010100001;
  assign mem[544] = 62'b11111110101010101100010000000110111101010111111000001100010111;
  assign mem[545] = 62'b11111111101111111101001101110001010100101100011011111011010011;
  assign mem[546] = 62'b11111111100111110001101011100010011100111000101101001100110011;
  assign mem[547] = 62'b11111111100101011010101100001101010001100101110110010010011111;
  assign mem[548] = 62'b11111111011011100010100111100000010100111111010101011010010011;
  assign mem[549] = 62'b11111111101100111000101011001100100111100110011010000001100000;
  assign mem[550] = 62'b11111111101110001010011000111101000100001110010001100101111010;
  assign mem[551] = 62'b11111111010101011000000100000000010010111101000110011110110100;
  assign mem[552] = 62'b11111111001111011110110111010010000000101111010011100000000010;
  assign mem[553] = 62'b11111111101111000001000101101000010100110011110111001110001100;
  assign mem[554] = 62'b11111111101011011111110110011010000110111001111001001011101001;
  assign mem[555] = 62'b11111111100000010111011111001111101100001100011011100010110111;
  assign mem[556] = 62'b11111111100011001001000010000111101100010010011010011000011111;
  assign mem[557] = 62'b11111111101001101001001101111110100100001010110000011010110010;
  assign mem[558] = 62'b11111111101111101010101111101111001011000011001111110111011100;
  assign mem[559] = 62'b11111111000010011001001001100101001101111111010011010000001001;
  assign mem[560] = 62'b11111111000011001010110111101111111001010001010001011010100111;
  assign mem[561] = 62'b11111111101111101000111001101110101100011110100001011110010001;
  assign mem[562] = 62'b11111111101001110000101101000100010000111100000111010111000010;
  assign mem[563] = 62'b11111111100010111110111100001001001011010001000001000000010101;
  assign mem[564] = 62'b11111111100000100010010001000100100000001100101011000010001100;
  assign mem[565] = 62'b11111111101011011001011000111100010100111111011011110001000111;
  assign mem[566] = 62'b11111111101111000100001001000010111100100010011000111101011111;
  assign mem[567] = 62'b11111111001110101110000110101101000110001011011110001101001000;
  assign mem[568] = 62'b11111111010101101111101110011110001011100111011011001110110110;
  assign mem[569] = 62'b11111111101110000110001010000000101111110111000110011011011001;
  assign mem[570] = 62'b11111111101100111110000011000011101000110011100100011001111011;
  assign mem[571] = 62'b11111111011011001011111001011100011101101100110001100101110010;
  assign mem[572] = 62'b11111111100101100100000000000111010101111101110010001111011111;
  assign mem[573] = 62'b11111111100111101001001111011100000111101111111001011111010010;
  assign mem[574] = 62'b11111111101111111101110101001110111011000110111001000101100100;
  assign mem[575] = 62'b11111110100111100011011011101010100101100001110100011010000110;
  assign mem[576] = 62'b11111110011100010001010100111101001100111001010011101100011101;
  assign mem[577] = 62'b11111111101111111111001110000010011100111000101010011001111001;
  assign mem[578] = 62'b11111111100111001111100101010110001110000001111001100101000010;
  assign mem[579] = 62'b11111111100101111111100111110010111101111001010110101000010000;
  assign mem[580] = 62'b11111111011010000111010110010101000011101101010000101011000000;
  assign mem[581] = 62'b11111111101101001101101111110001111011110010111111101111011100;
  assign mem[582] = 62'b11111111101101111001000001011000001111011011011000110110000001;
  assign mem[583] = 62'b11111111010110110110011001100001100011100010100000110010110110;
  assign mem[584] = 62'b11111111001100011011011001000001010011010111010111010011011101;
  assign mem[585] = 62'b11111111101111001100110110100001011010001110101010111011110000;
  assign mem[586] = 62'b11111111101011000101100111010000101010010011001010001011110101;
  assign mem[587] = 62'b11111111100001000010010111001001001000110100001010100101010111;
  assign mem[588] = 62'b11111111100010100000011000101111101111010011010011110010111010;
  assign mem[589] = 62'b11111111101010000110110010011011010010110000001010011101011110;
  assign mem[590] = 62'b11111111101111100010111010011100110111110010110100101101111000;
  assign mem[591] = 62'b11111111000101011111110000000010000110010101001100101111011110;
  assign mem[592] = 62'b11111111000000000011101110100010101101011011111011100001011011;
  assign mem[593] = 62'b11111111101111101111110100011100001111000010101000110110001000;
  assign mem[594] = 62'b11111111101001010010011001000011100011101011000100101001101100;
  assign mem[595] = 62'b11111111100011100111000010001111100011110101100011000000101001;
  assign mem[596] = 62'b11111111011111101101110101011101011100001001001101001011011110;
  assign mem[597] = 62'b11111111101011110010110101010011001011000011010010001100100111;
  assign mem[598] = 62'b11111111101110110111011110101101101010000001111000011001010001;
  assign mem[599] = 62'b11111111010000111000010101101101001110000101110100100111001110;
  assign mem[600] = 62'b11111111010100010000110001000011011100100010010011011011110000;
  assign mem[601] = 62'b11111111101110010110101001110101010101000001000110011111010011;
  assign mem[602] = 62'b11111111101100101000001000111100011001101110011100010001001001;
  assign mem[603] = 62'b11111111011100100110010111111111000011100001100101001110001001;
  assign mem[604] = 62'b11111111100100111110011100110000100101110011001010010010000110;
  assign mem[605] = 62'b11111111101000001010101001110000010011111101010100010111111111;
  assign mem[606] = 62'b11111111101111111010111001110100100101001100000100000100001111;
  assign mem[607] = 62'b11111110110010000011001001011001110100111011010100010001001101;
  assign mem[608] = 62'b11111110110011100111011001111100010010110001011010001010011001;
  assign mem[609] = 62'b11111111101111111001111110101010000101010010000010110101100000;
  assign mem[610] = 62'b11111111101000010010110111000100010001101011111000001111111010;
  assign mem[611] = 62'b11111111100100110100111011110001101101010110001001111101111111;
  assign mem[612] = 62'b11111111011100111100110100101110101110111000011100110100100001;
  assign mem[613] = 62'b11111111101100100010011111010110000111000000101001110000010011;
  assign mem[614] = 62'b11111111101110011010100110000111000101010111010101001110100111;
  assign mem[615] = 62'b11111111010011111000111001101111101001011011101100001001110001;
  assign mem[616] = 62'b11111111010001010000100011111011101111110001101001001101111000;
  assign mem[617] = 62'b11111111101110110100001000001101011110100110011001000000001001;
  assign mem[618] = 62'b11111111101011111001000001101101100001000100010101010011000001;
  assign mem[619] = 62'b11111111011111010111111101111011100110010101101100110110100011;
  assign mem[620] = 62'b11111111100011110000111100010001001001100000011100010100011000;
  assign mem[621] = 62'b11111111101001001010101010010000011111110001011010100000010101;
  assign mem[622] = 62'b11111111101111110001010110111000111011011111011001101011110110;
  assign mem[623] = 62'b11111110111110100011101011011111111101111001001010101000111111;
  assign mem[624] = 62'b11111111000110010001010001101010000011000111011000001100001101;
  assign mem[625] = 62'b11111111101111100000110000111101001010010000001100011000001100;
  assign mem[626] = 62'b11111111101010001110000001100001001010010110010011101111000110;
  assign mem[627] = 62'b11111111100010010110000111001101001100101110110111000100010000;
  assign mem[628] = 62'b11111111100001001100111110100111001111111011100010010101001111;
  assign mem[629] = 62'b11111111101010111110111000111111011000100111110101011110110110;
  assign mem[630] = 62'b11111111101111001111100110101110111100000110111011110001100101;
  assign mem[631] = 62'b11111111001011101010010110001100110100111100010101110110101101;
  assign mem[632] = 62'b11111111010111001101110110001111001001001001100001000010010010;
  assign mem[633] = 62'b11111111101101110100011111111011110011100010101001000101011010;
  assign mem[634] = 62'b11111111101101010010110101101100011011000110000111010100100100;
  assign mem[635] = 62'b11111111011001110000010111110101000100000011011111100111110010;
  assign mem[636] = 62'b11111111100110001000101110010001001111111011000010001011111111;
  assign mem[637] = 62'b11111111100111000110111010110010010110000011100100000110111111;
  assign mem[638] = 62'b11111111101111111111100001110001101000011100001100101101110111;
  assign mem[639] = 62'b11111110010101111111010100110100100001111110101011001000100110;
  assign mem[640] = 62'b11111110001111011010100010100101101010101110011001011111001011;
  assign mem[641] = 62'b11111111101111111111110000100101000011110001010011101111010001;
  assign mem[642] = 62'b11111111100110111110001100101010011001110010010101101101110101;
  assign mem[643] = 62'b11111111100110010001110001010101000011011111110101001101011011;
  assign mem[644] = 62'b11111111011001011001010101010110110111101010111001010010001111;
  assign mem[645] = 62'b11111111101101010111110111000101110010100010001000101001111111;
  assign mem[646] = 62'b11111111101101101111111001111001000011100101010111010110011010;
  assign mem[647] = 62'b11111111010111100101001111010111100110000100111101111110101110;
  assign mem[648] = 62'b11111111001010111001001111000111010101111100111011100110101011;
  assign mem[649] = 62'b11111111101111010010010010001000000110101111001010101110110100;
  assign mem[650] = 62'b11111111101010111000000110100011110011010001011110110011101111;
  assign mem[651] = 62'b11111111100001010111100011011011100100110110111110001010111100;
  assign mem[652] = 62'b11111111100010001011110010110101100110001011000001001111100010;
  assign mem[653] = 62'b11111111101010010101001100100100010000100100001111010100100011;
  assign mem[654] = 62'b11111111101111011110100010100110011100000110100011001000101010;
  assign mem[655] = 62'b11111111000111000010101111110110001101000010001100010011111111;
  assign mem[656] = 62'b11111110111100111111110101001100111011001100000111110111000001;
  assign mem[657] = 62'b11111111101111110010110100011100000011100100010100001101010100;
  assign mem[658] = 62'b11111111101001000010110111100101000011010101110101111011111110;
  assign mem[659] = 62'b11111111100011111010110011001111101010101111100000011010000000;
  assign mem[660] = 62'b11111111011111000010000001100100000110101111111111011111111110;
  assign mem[661] = 62'b11111111101011111111001001110100100101101000011011000101000111;
  assign mem[662] = 62'b11111111101110110000101100111101001011000110101111011010110010;
  assign mem[663] = 62'b11111111010001101000101111011111111011111010001111001001000011;
  assign mem[664] = 62'b11111111010011100000111111010111100011010100111011011010101011;
  assign mem[665] = 62'b11111111101110011110011101101100101001101001010001011001011010;
  assign mem[666] = 62'b11111111101100011100110001010110001001100111101010101011010111;
  assign mem[667] = 62'b11111111011101010011001101000000101011101010000110000010011101;
  assign mem[668] = 62'b11111111100100101011010111100101010001011001110010001011110001;
  assign mem[669] = 62'b11111111101000011011000000101000011101100110101010000110010101;
  assign mem[670] = 62'b11111111101111111000111110100100101011111010011101100010000110;
  assign mem[671] = 62'b11111110110101001011100111011101001010010011010100110100001010;
  assign mem[672] = 62'b11111110110000011110110110000101001110010001100011000001100100;
  assign mem[673] = 62'b11111111101111111011110000000100000010100000100110000110010001;
  assign mem[674] = 62'b11111111101000000010011000101101110101011011100101001011111010;
  assign mem[675] = 62'b11111111100101000111111010100000011100110110011001101010100110;
  assign mem[676] = 62'b11111111011100001111110110110101000111001001100011000100101001;
  assign mem[677] = 62'b11111111101100101101101110001000001010000000001101101010011001;
  assign mem[678] = 62'b11111111101110010010101000110111111111100000011100111001011110;
  assign mem[679] = 62'b11111111010100101000100101001111010001000110111000001011110011;
  assign mem[680] = 62'b11111111010000100000000100111000000101111010110110011000011110;
  assign mem[681] = 62'b11111111101110111010110000011101001100010100001010010101000100;
  assign mem[682] = 62'b11111111101011101100100100100110100000101101101100010000001101;
  assign mem[683] = 62'b11111111100000000001110100000011001000001010111000001011100001;
  assign mem[684] = 62'b11111111100011011101000101001100011011100000010111111110001101;
  assign mem[685] = 62'b11111111101001011010000011111101000010101111010111111111100001;
  assign mem[686] = 62'b11111111101111101110001101000110001101011001101010110110110111;
  assign mem[687] = 62'b11111111000000110101100100110110111100101100100110011110000110;
  assign mem[688] = 62'b11111111000100101110001011000101111111011110011111101010001000;
  assign mem[689] = 62'b11111111101111100100111111000101001111100001011010110000001000;
  assign mem[690] = 62'b11111111101001111111011111010011110001001100010100100111011110;
  assign mem[691] = 62'b11111111100010101010100111011011101000011110101110101101011000;
  assign mem[692] = 62'b11111111100000110111101101000010111000010010111100010010110110;
  assign mem[693] = 62'b11111111101011001100010001010110100101111100110111101111110011;
  assign mem[694] = 62'b11111111101111001010000001011111111100010001100000100111001110;
  assign mem[695] = 62'b11111111001101001100010111011101001101001011001011110111101110;
  assign mem[696] = 62'b11111111010110011110111001010010011100101011010110001111001011;
  assign mem[697] = 62'b11111111101101111101011110001101101010100110111010010110011100;
  assign mem[698] = 62'b11111111101101001000100101010111000110111001011010010011100001;
  assign mem[699] = 62'b11111111011010011110010000110011010011110110111111001100011011;
  assign mem[700] = 62'b11111111100101110110011101111011100111001111100011010001011100;
  assign mem[701] = 62'b11111111100111011000001100010100101100001100000100011101100100;
  assign mem[702] = 62'b11111111101111111110110101010111100100001001011111110110101110;
  assign mem[703] = 62'b11111110100001010001101000010111011011010000101100000101111111;
  assign mem[704] = 62'b11111110100100011010100011100101101111111110000110000101111001;
  assign mem[705] = 62'b11111111101111111110010111110001000010000010001100000000010100;
  assign mem[706] = 62'b11111111100111100000101111101100011011100100001011001101011011;
  assign mem[707] = 62'b11111111100101101101010000101100100110010011110111010001001000;
  assign mem[708] = 62'b11111111011010110101000111001100010010010111001101110000001001;
  assign mem[709] = 62'b11111111101101000011010110011100101111010110011101001010111001;
  assign mem[710] = 62'b11111111101110000001110110011011011001001010000000111101010100;
  assign mem[711] = 62'b11111111010110000111010101100101011100100010001100001000000010;
  assign mem[712] = 62'b11111111001101111101010001011000111111000000010000100110011010;
  assign mem[713] = 62'b11111111101111000111000111101010111110001010000100011100001000;
  assign mem[714] = 62'b11111111101011010010110111010000001001110111100111100100100101;
  assign mem[715] = 62'b11111111100000101101000000010110000111100011111000010111101100;
  assign mem[716] = 62'b11111111100010110100110011001111010011010011101001101110111000;
  assign mem[717] = 62'b11111111101001111000001000001011101101101101000010010001110010;
  assign mem[718] = 62'b11111111101111100110111110110101111100111110111101111000101001;
  assign mem[719] = 62'b11111111000011111100100010111101010111110110110100100010010011;
  assign mem[720] = 62'b11111111000001100111011000100101000000101111100010010011100111;
  assign mem[721] = 62'b11111111101111101100100000110111000110100000011101010101001101;
  assign mem[722] = 62'b11111111101001100001101010111011110001010001010111010110010100;
  assign mem[723] = 62'b11111111100011010011000101001001010010110000010100110111100001;
  assign mem[724] = 62'b11111111100000001100101010111001010101111011011011110110010110;
  assign mem[725] = 62'b11111111101011100110001111101000011111110110010001010101011110;
  assign mem[726] = 62'b11111111101110111101111101011011100101000111001010001111000000;
  assign mem[727] = 62'b11111111010000000111110001100000000110101110011111110111010010;
  assign mem[728] = 62'b11111111010101000000010110001111011100000110010111000001001000;
  assign mem[729] = 62'b11111111101110001110100011001111101100011101011100111010000101;
  assign mem[730] = 62'b11111111101100110011001110111000100000110000101101111010100000;
  assign mem[731] = 62'b11111111011011111001010001010100010111111111111100000011011001;
  assign mem[732] = 62'b11111111100101010001010100111111110101000101011001110111111100;
  assign mem[733] = 62'b11111111100111111010000011111110000111101100000011011010000110;
  assign mem[734] = 62'b11111111101111111100100001011000010100111000010011000111101101;
  assign mem[735] = 62'b11111110101101110101000000011011111001100000001000111011001001;
  assign mem[736] = 62'b11111110110110101111110001101100111110011110011011000100101001;
  assign mem[737] = 62'b11111111101111110111111001100100100010111101110011001100000111;
  assign mem[738] = 62'b11111111101000100011000110011011100111010010000001101110100001;
  assign mem[739] = 62'b11111111100100100001110000001100110000011000001001000111111111;
  assign mem[740] = 62'b11111111011101101001100000110001011100111110100001000011011001;
  assign mem[741] = 62'b11111111101100010110111110111101011001111111101111100001011010;
  assign mem[742] = 62'b11111111101110100010010000100101011011101011010110000000100101;
  assign mem[743] = 62'b11111111010011001001000001111110110110001110001011101010101111;
  assign mem[744] = 62'b11111111010010000000111000010110000011110101110010011110111110;
  assign mem[745] = 62'b11111111101110101101001100111101010001010110111000100000010001;
  assign mem[746] = 62'b11111111101100000101001101100111011100010001100101111001010111;
  assign mem[747] = 62'b11111111011110101100000000011010010101111100100101011000100000;
  assign mem[748] = 62'b11111111100100000100100111001001100110001111010001000010001100;
  assign mem[749] = 62'b11111111101000111011000001000010011011010010000110110001001001;
  assign mem[750] = 62'b11111111101111110100001101000101011000110110000110000010000111;
  assign mem[751] = 62'b11111110111011011011111010011011101100001110001111011001001100;
  assign mem[752] = 62'b11111111000111110100001010011110111011110100101100101100011100;
  assign mem[753] = 62'b11111111101111011100001111011001000011010010110111111010110111;
  assign mem[754] = 62'b11111111101010011100010011100011011110100111010110000011110101;
  assign mem[755] = 62'b11111111100010000001011011101010100001011101010110000011010110;
  assign mem[756] = 62'b11111111100001100010000101100100011111001110100100011011100101;
  assign mem[757] = 62'b11111111101010110001001111111110111101001111101111101011001000;
  assign mem[758] = 62'b11111111101111010100111000101100011111101011110010110100000111;
  assign mem[759] = 62'b11111111001010001000000011111000011011000110000011000111011010;
  assign mem[760] = 62'b11111111010111111100100100110111010011011100110100000111100100;
  assign mem[761] = 62'b11111111101101101011001111010000101100111001101000101010111001;
  assign mem[762] = 62'b11111111101101011100110011111101010000100011000000110111111111;
  assign mem[763] = 62'b11111111011001000010001110111110000001111011110111101111010001;
  assign mem[764] = 62'b11111111100110011010110000111100111111010100101011001110000110;
  assign mem[765] = 62'b11111111100110110101011010111111101111010010101010111111001101;
  assign mem[766] = 62'b11111111101111111111111010011100101100100101111000110001001111;
  assign mem[767] = 62'b11111110000010110110010110101100001110010100001001011100000011;
  assign mem[768] = 62'b11111110000010110110010110101100001110010100001001011100000011;
  assign mem[769] = 62'b11111111101111111111111010011100101100100101111000110001001111;
  assign mem[770] = 62'b11111111100110110101011010111111101111010010101010111111001101;
  assign mem[771] = 62'b11111111100110011010110000111100111111010100101011001110000110;
  assign mem[772] = 62'b11111111011001000010001110111110000001111011110111101111010001;
  assign mem[773] = 62'b11111111101101011100110011111101010000100011000000110111111111;
  assign mem[774] = 62'b11111111101101101011001111010000101100111001101000101010111001;
  assign mem[775] = 62'b11111111010111111100100100110111010011011100110100000111100100;
  assign mem[776] = 62'b11111111001010001000000011111000011011000110000011000111011010;
  assign mem[777] = 62'b11111111101111010100111000101100011111101011110010110100000111;
  assign mem[778] = 62'b11111111101010110001001111111110111101001111101111101011001000;
  assign mem[779] = 62'b11111111100001100010000101100100011111001110100100011011100101;
  assign mem[780] = 62'b11111111100010000001011011101010100001011101010110000011010110;
  assign mem[781] = 62'b11111111101010011100010011100011011110100111010110000011110101;
  assign mem[782] = 62'b11111111101111011100001111011001000011010010110111111010110111;
  assign mem[783] = 62'b11111111000111110100001010011110111011110100101100101100011100;
  assign mem[784] = 62'b11111110111011011011111010011011101100001110001111011001001100;
  assign mem[785] = 62'b11111111101111110100001101000101011000110110000110000010000111;
  assign mem[786] = 62'b11111111101000111011000001000010011011010010000110110001001001;
  assign mem[787] = 62'b11111111100100000100100111001001100110001111010001000010001100;
  assign mem[788] = 62'b11111111011110101100000000011010010101111100100101011000100000;
  assign mem[789] = 62'b11111111101100000101001101100111011100010001100101111001010111;
  assign mem[790] = 62'b11111111101110101101001100111101010001010110111000100000010001;
  assign mem[791] = 62'b11111111010010000000111000010110000011110101110010011110111110;
  assign mem[792] = 62'b11111111010011001001000001111110110110001110001011101010101111;
  assign mem[793] = 62'b11111111101110100010010000100101011011101011010110000000100101;
  assign mem[794] = 62'b11111111101100010110111110111101011001111111101111100001011010;
  assign mem[795] = 62'b11111111011101101001100000110001011100111110100001000011011001;
  assign mem[796] = 62'b11111111100100100001110000001100110000011000001001000111111111;
  assign mem[797] = 62'b11111111101000100011000110011011100111010010000001101110100001;
  assign mem[798] = 62'b11111111101111110111111001100100100010111101110011001100000111;
  assign mem[799] = 62'b11111110110110101111110001101100111110011110011011000100101001;
  assign mem[800] = 62'b11111110101101110101000000011011111001100000001000111011001001;
  assign mem[801] = 62'b11111111101111111100100001011000010100111000010011000111101101;
  assign mem[802] = 62'b11111111100111111010000011111110000111101100000011011010000110;
  assign mem[803] = 62'b11111111100101010001010100111111110101000101011001110111111100;
  assign mem[804] = 62'b11111111011011111001010001010100010111111111111100000011011001;
  assign mem[805] = 62'b11111111101100110011001110111000100000110000101101111010100000;
  assign mem[806] = 62'b11111111101110001110100011001111101100011101011100111010000101;
  assign mem[807] = 62'b11111111010101000000010110001111011100000110010111000001001000;
  assign mem[808] = 62'b11111111010000000111110001100000000110101110011111110111010010;
  assign mem[809] = 62'b11111111101110111101111101011011100101000111001010001111000000;
  assign mem[810] = 62'b11111111101011100110001111101000011111110110010001010101011110;
  assign mem[811] = 62'b11111111100000001100101010111001010101111011011011110110010110;
  assign mem[812] = 62'b11111111100011010011000101001001010010110000010100110111100001;
  assign mem[813] = 62'b11111111101001100001101010111011110001010001010111010110010100;
  assign mem[814] = 62'b11111111101111101100100000110111000110100000011101010101001101;
  assign mem[815] = 62'b11111111000001100111011000100101000000101111100010010011100111;
  assign mem[816] = 62'b11111111000011111100100010111101010111110110110100100010010011;
  assign mem[817] = 62'b11111111101111100110111110110101111100111110111101111000101001;
  assign mem[818] = 62'b11111111101001111000001000001011101101101101000010010001110010;
  assign mem[819] = 62'b11111111100010110100110011001111010011010011101001101110111000;
  assign mem[820] = 62'b11111111100000101101000000010110000111100011111000010111101100;
  assign mem[821] = 62'b11111111101011010010110111010000001001110111100111100100100101;
  assign mem[822] = 62'b11111111101111000111000111101010111110001010000100011100001000;
  assign mem[823] = 62'b11111111001101111101010001011000111111000000010000100110011010;
  assign mem[824] = 62'b11111111010110000111010101100101011100100010001100001000000010;
  assign mem[825] = 62'b11111111101110000001110110011011011001001010000000111101010100;
  assign mem[826] = 62'b11111111101101000011010110011100101111010110011101001010111001;
  assign mem[827] = 62'b11111111011010110101000111001100010010010111001101110000001001;
  assign mem[828] = 62'b11111111100101101101010000101100100110010011110111010001001000;
  assign mem[829] = 62'b11111111100111100000101111101100011011100100001011001101011011;
  assign mem[830] = 62'b11111111101111111110010111110001000010000010001100000000010100;
  assign mem[831] = 62'b11111110100100011010100011100101101111111110000110000101111001;
  assign mem[832] = 62'b11111110100001010001101000010111011011010000101100000101111111;
  assign mem[833] = 62'b11111111101111111110110101010111100100001001011111110110101110;
  assign mem[834] = 62'b11111111100111011000001100010100101100001100000100011101100100;
  assign mem[835] = 62'b11111111100101110110011101111011100111001111100011010001011100;
  assign mem[836] = 62'b11111111011010011110010000110011010011110110111111001100011011;
  assign mem[837] = 62'b11111111101101001000100101010111000110111001011010010011100001;
  assign mem[838] = 62'b11111111101101111101011110001101101010100110111010010110011100;
  assign mem[839] = 62'b11111111010110011110111001010010011100101011010110001111001011;
  assign mem[840] = 62'b11111111001101001100010111011101001101001011001011110111101110;
  assign mem[841] = 62'b11111111101111001010000001011111111100010001100000100111001110;
  assign mem[842] = 62'b11111111101011001100010001010110100101111100110111101111110011;
  assign mem[843] = 62'b11111111100000110111101101000010111000010010111100010010110110;
  assign mem[844] = 62'b11111111100010101010100111011011101000011110101110101101011000;
  assign mem[845] = 62'b11111111101001111111011111010011110001001100010100100111011110;
  assign mem[846] = 62'b11111111101111100100111111000101001111100001011010110000001000;
  assign mem[847] = 62'b11111111000100101110001011000101111111011110011111101010001000;
  assign mem[848] = 62'b11111111000000110101100100110110111100101100100110011110000110;
  assign mem[849] = 62'b11111111101111101110001101000110001101011001101010110110110111;
  assign mem[850] = 62'b11111111101001011010000011111101000010101111010111111111100001;
  assign mem[851] = 62'b11111111100011011101000101001100011011100000010111111110001101;
  assign mem[852] = 62'b11111111100000000001110100000011001000001010111000001011100001;
  assign mem[853] = 62'b11111111101011101100100100100110100000101101101100010000001101;
  assign mem[854] = 62'b11111111101110111010110000011101001100010100001010010101000100;
  assign mem[855] = 62'b11111111010000100000000100111000000101111010110110011000011110;
  assign mem[856] = 62'b11111111010100101000100101001111010001000110111000001011110011;
  assign mem[857] = 62'b11111111101110010010101000110111111111100000011100111001011110;
  assign mem[858] = 62'b11111111101100101101101110001000001010000000001101101010011001;
  assign mem[859] = 62'b11111111011100001111110110110101000111001001100011000100101001;
  assign mem[860] = 62'b11111111100101000111111010100000011100110110011001101010100110;
  assign mem[861] = 62'b11111111101000000010011000101101110101011011100101001011111010;
  assign mem[862] = 62'b11111111101111111011110000000100000010100000100110000110010001;
  assign mem[863] = 62'b11111110110000011110110110000101001110010001100011000001100100;
  assign mem[864] = 62'b11111110110101001011100111011101001010010011010100110100001010;
  assign mem[865] = 62'b11111111101111111000111110100100101011111010011101100010000110;
  assign mem[866] = 62'b11111111101000011011000000101000011101100110101010000110010101;
  assign mem[867] = 62'b11111111100100101011010111100101010001011001110010001011110001;
  assign mem[868] = 62'b11111111011101010011001101000000101011101010000110000010011101;
  assign mem[869] = 62'b11111111101100011100110001010110001001100111101010101011010111;
  assign mem[870] = 62'b11111111101110011110011101101100101001101001010001011001011010;
  assign mem[871] = 62'b11111111010011100000111111010111100011010100111011011010101011;
  assign mem[872] = 62'b11111111010001101000101111011111111011111010001111001001000011;
  assign mem[873] = 62'b11111111101110110000101100111101001011000110101111011010110010;
  assign mem[874] = 62'b11111111101011111111001001110100100101101000011011000101000111;
  assign mem[875] = 62'b11111111011111000010000001100100000110101111111111011111111110;
  assign mem[876] = 62'b11111111100011111010110011001111101010101111100000011010000000;
  assign mem[877] = 62'b11111111101001000010110111100101000011010101110101111011111110;
  assign mem[878] = 62'b11111111101111110010110100011100000011100100010100001101010100;
  assign mem[879] = 62'b11111110111100111111110101001100111011001100000111110111000001;
  assign mem[880] = 62'b11111111000111000010101111110110001101000010001100010011111111;
  assign mem[881] = 62'b11111111101111011110100010100110011100000110100011001000101010;
  assign mem[882] = 62'b11111111101010010101001100100100010000100100001111010100100011;
  assign mem[883] = 62'b11111111100010001011110010110101100110001011000001001111100010;
  assign mem[884] = 62'b11111111100001010111100011011011100100110110111110001010111100;
  assign mem[885] = 62'b11111111101010111000000110100011110011010001011110110011101111;
  assign mem[886] = 62'b11111111101111010010010010001000000110101111001010101110110100;
  assign mem[887] = 62'b11111111001010111001001111000111010101111100111011100110101011;
  assign mem[888] = 62'b11111111010111100101001111010111100110000100111101111110101110;
  assign mem[889] = 62'b11111111101101101111111001111001000011100101010111010110011010;
  assign mem[890] = 62'b11111111101101010111110111000101110010100010001000101001111111;
  assign mem[891] = 62'b11111111011001011001010101010110110111101010111001010010001111;
  assign mem[892] = 62'b11111111100110010001110001010101000011011111110101001101011011;
  assign mem[893] = 62'b11111111100110111110001100101010011001110010010101101101110101;
  assign mem[894] = 62'b11111111101111111111110000100101000011110001010011101111010001;
  assign mem[895] = 62'b11111110001111011010100010100101101010101110011001011111001011;
  assign mem[896] = 62'b11111110010101111111010100110100100001111110101011001000100110;
  assign mem[897] = 62'b11111111101111111111100001110001101000011100001100101101110111;
  assign mem[898] = 62'b11111111100111000110111010110010010110000011100100000110111111;
  assign mem[899] = 62'b11111111100110001000101110010001001111111011000010001011111111;
  assign mem[900] = 62'b11111111011001110000010111110101000100000011011111100111110010;
  assign mem[901] = 62'b11111111101101010010110101101100011011000110000111010100100100;
  assign mem[902] = 62'b11111111101101110100011111111011110011100010101001000101011010;
  assign mem[903] = 62'b11111111010111001101110110001111001001001001100001000010010010;
  assign mem[904] = 62'b11111111001011101010010110001100110100111100010101110110101101;
  assign mem[905] = 62'b11111111101111001111100110101110111100000110111011110001100101;
  assign mem[906] = 62'b11111111101010111110111000111111011000100111110101011110110110;
  assign mem[907] = 62'b11111111100001001100111110100111001111111011100010010101001111;
  assign mem[908] = 62'b11111111100010010110000111001101001100101110110111000100010000;
  assign mem[909] = 62'b11111111101010001110000001100001001010010110010011101111000110;
  assign mem[910] = 62'b11111111101111100000110000111101001010010000001100011000001100;
  assign mem[911] = 62'b11111111000110010001010001101010000011000111011000001100001101;
  assign mem[912] = 62'b11111110111110100011101011011111111101111001001010101000111111;
  assign mem[913] = 62'b11111111101111110001010110111000111011011111011001101011110110;
  assign mem[914] = 62'b11111111101001001010101010010000011111110001011010100000010101;
  assign mem[915] = 62'b11111111100011110000111100010001001001100000011100010100011000;
  assign mem[916] = 62'b11111111011111010111111101111011100110010101101100110110100011;
  assign mem[917] = 62'b11111111101011111001000001101101100001000100010101010011000001;
  assign mem[918] = 62'b11111111101110110100001000001101011110100110011001000000001001;
  assign mem[919] = 62'b11111111010001010000100011111011101111110001101001001101111000;
  assign mem[920] = 62'b11111111010011111000111001101111101001011011101100001001110001;
  assign mem[921] = 62'b11111111101110011010100110000111000101010111010101001110100111;
  assign mem[922] = 62'b11111111101100100010011111010110000111000000101001110000010011;
  assign mem[923] = 62'b11111111011100111100110100101110101110111000011100110100100001;
  assign mem[924] = 62'b11111111100100110100111011110001101101010110001001111101111111;
  assign mem[925] = 62'b11111111101000010010110111000100010001101011111000001111111010;
  assign mem[926] = 62'b11111111101111111001111110101010000101010010000010110101100000;
  assign mem[927] = 62'b11111110110011100111011001111100010010110001011010001010011001;
  assign mem[928] = 62'b11111110110010000011001001011001110100111011010100010001001101;
  assign mem[929] = 62'b11111111101111111010111001110100100101001100000100000100001111;
  assign mem[930] = 62'b11111111101000001010101001110000010011111101010100010111111111;
  assign mem[931] = 62'b11111111100100111110011100110000100101110011001010010010000110;
  assign mem[932] = 62'b11111111011100100110010111111111000011100001100101001110001001;
  assign mem[933] = 62'b11111111101100101000001000111100011001101110011100010001001001;
  assign mem[934] = 62'b11111111101110010110101001110101010101000001000110011111010011;
  assign mem[935] = 62'b11111111010100010000110001000011011100100010010011011011110000;
  assign mem[936] = 62'b11111111010000111000010101101101001110000101110100100111001110;
  assign mem[937] = 62'b11111111101110110111011110101101101010000001111000011001010001;
  assign mem[938] = 62'b11111111101011110010110101010011001011000011010010001100100111;
  assign mem[939] = 62'b11111111011111101101110101011101011100001001001101001011011110;
  assign mem[940] = 62'b11111111100011100111000010001111100011110101100011000000101001;
  assign mem[941] = 62'b11111111101001010010011001000011100011101011000100101001101100;
  assign mem[942] = 62'b11111111101111101111110100011100001111000010101000110110001000;
  assign mem[943] = 62'b11111111000000000011101110100010101101011011111011100001011011;
  assign mem[944] = 62'b11111111000101011111110000000010000110010101001100101111011110;
  assign mem[945] = 62'b11111111101111100010111010011100110111110010110100101101111000;
  assign mem[946] = 62'b11111111101010000110110010011011010010110000001010011101011110;
  assign mem[947] = 62'b11111111100010100000011000101111101111010011010011110010111010;
  assign mem[948] = 62'b11111111100001000010010111001001001000110100001010100101010111;
  assign mem[949] = 62'b11111111101011000101100111010000101010010011001010001011110101;
  assign mem[950] = 62'b11111111101111001100110110100001011010001110101010111011110000;
  assign mem[951] = 62'b11111111001100011011011001000001010011010111010111010011011101;
  assign mem[952] = 62'b11111111010110110110011001100001100011100010100000110010110110;
  assign mem[953] = 62'b11111111101101111001000001011000001111011011011000110110000001;
  assign mem[954] = 62'b11111111101101001101101111110001111011110010111111101111011100;
  assign mem[955] = 62'b11111111011010000111010110010101000011101101010000101011000000;
  assign mem[956] = 62'b11111111100101111111100111110010111101111001010110101000010000;
  assign mem[957] = 62'b11111111100111001111100101010110001110000001111001100101000010;
  assign mem[958] = 62'b11111111101111111111001110000010011100111000101010011001111001;
  assign mem[959] = 62'b11111110011100010001010100111101001100111001010011101100011101;
  assign mem[960] = 62'b11111110100111100011011011101010100101100001110100011010000110;
  assign mem[961] = 62'b11111111101111111101110101001110111011000110111001000101100100;
  assign mem[962] = 62'b11111111100111101001001111011100000111101111111001011111010010;
  assign mem[963] = 62'b11111111100101100100000000000111010101111101110010001111011111;
  assign mem[964] = 62'b11111111011011001011111001011100011101101100110001100101110010;
  assign mem[965] = 62'b11111111101100111110000011000011101000110011100100011001111011;
  assign mem[966] = 62'b11111111101110000110001010000000101111110111000110011011011001;
  assign mem[967] = 62'b11111111010101101111101110011110001011100111011011001110110110;
  assign mem[968] = 62'b11111111001110101110000110101101000110001011011110001101001000;
  assign mem[969] = 62'b11111111101111000100001001000010111100100010011000111101011111;
  assign mem[970] = 62'b11111111101011011001011000111100010100111111011011110001000111;
  assign mem[971] = 62'b11111111100000100010010001000100100000001100101011000010001100;
  assign mem[972] = 62'b11111111100010111110111100001001001011010001000001000000010101;
  assign mem[973] = 62'b11111111101001110000101101000100010000111100000111010111000010;
  assign mem[974] = 62'b11111111101111101000111001101110101100011110100001011110010001;
  assign mem[975] = 62'b11111111000011001010110111101111111001010001010001011010100111;
  assign mem[976] = 62'b11111111000010011001001001100101001101111111010011010000001001;
  assign mem[977] = 62'b11111111101111101010101111101111001011000011001111110111011100;
  assign mem[978] = 62'b11111111101001101001001101111110100100001010110000011010110010;
  assign mem[979] = 62'b11111111100011001001000010000111101100010010011010011000011111;
  assign mem[980] = 62'b11111111100000010111011111001111101100001100011011100010110111;
  assign mem[981] = 62'b11111111101011011111110110011010000110111001111001001011101001;
  assign mem[982] = 62'b11111111101111000001000101101000010100110011110111001110001100;
  assign mem[983] = 62'b11111111001111011110110111010010000000101111010011100000000010;
  assign mem[984] = 62'b11111111010101011000000100000000010010111101000110011110110100;
  assign mem[985] = 62'b11111111101110001010011000111101000100001110010001100101111010;
  assign mem[986] = 62'b11111111101100111000101011001100100111100110011010000001100000;
  assign mem[987] = 62'b11111111011011100010100111100000010100111111010101011010010011;
  assign mem[988] = 62'b11111111100101011010101100001101010001100101110110010010011111;
  assign mem[989] = 62'b11111111100111110001101011100010011100111000101101001100110011;
  assign mem[990] = 62'b11111111101111111101001101110001010100101100011011111011010011;
  assign mem[991] = 62'b11111110101010101100010000000110111101010111111000001100010111;
  assign mem[992] = 62'b11111110111000010011111000011100010010110000010011000010100001;
  assign mem[993] = 62'b11111111101111110110101111101001110101000101000101001110001100;
  assign mem[994] = 62'b11111111101000101011001000011100011110110111100001110110001000;
  assign mem[995] = 62'b11111111100100011000000101101001101001001010110011001010100010;
  assign mem[996] = 62'b11111111011101111111101111111101100110101010010100000111011110;
  assign mem[997] = 62'b11111111101100010001001000001100110001010000011100000000000100;
  assign mem[998] = 62'b11111111101110100101111110110000110110000000010110101100110000;
  assign mem[999] = 62'b11111111010010110001000001101001001110100101010100010100100000;
  assign mem[1000] = 62'b11111111010010011000111110011010011001010101010101010010111010;
  assign mem[1001] = 62'b11111111101110101001101000001110010011111001100101100000000000;
  assign mem[1002] = 62'b11111111101100001011001101000101001001001100011110001111110001;
  assign mem[1003] = 62'b11111111011110010101111010100001101101001111001101100000100101;
  assign mem[1004] = 62'b11111111100100001110010111111101011011001010100100001110000000;
  assign mem[1005] = 62'b11111111101000110011000110101001110101000110000100011001010101;
  assign mem[1006] = 62'b11111111101111110101100000110100101101101001110101110010011110;
  assign mem[1007] = 62'b11111110111001110111111011011011101011001001001010100001011100;
  assign mem[1008] = 62'b11111111001000100101100001011100100111110001000001100000000100;
  assign mem[1009] = 62'b11111111101111011001110111010101010110100010000011110011101110;
  assign mem[1010] = 62'b11111111101010100011010110011101101110010101000101101011010010;
  assign mem[1011] = 62'b11111111100001110111000001101101100100110111000100100001110010;
  assign mem[1012] = 62'b11111111100001101100100101000000010111000100110111001110111111;
  assign mem[1013] = 62'b11111111101010101010010101010001111010001011001011100110001110;
  assign mem[1014] = 62'b11111111101111010111011010011011101101010000110110100001011101;
  assign mem[1015] = 62'b11111111001001010110110100100111101001101101100010101011111010;
  assign mem[1016] = 62'b11111111011000010011110110101010101010111100111001000000111111;
  assign mem[1017] = 62'b11111111101101100110100000000011011101100010110011110101000110;
  assign mem[1018] = 62'b11111111101101100001101100010010000100010001011010010001001111;
  assign mem[1019] = 62'b11111111011000101011000100101110000110110101011110110101000100;
  assign mem[1020] = 62'b11111111100110100011101101000111101010101000011001110001110001;
  assign mem[1021] = 62'b11111111100110101100100101110011101101001011111110001010011100;
  assign mem[1022] = 62'b11111111101111111111111111011000100001011000100001110100000010;
  assign mem[1023] = 62'b11111101101001001000011111100010111110110011001010010010111010;

  always@(*)
  begin
    data_out_t <= mem[addr_f];
  end

  // Build output registers
  wire [61:0] data_out_reg [n_outreg:0];
  generate if (n_outreg > 0)
  begin
    for( i=n_outreg-1; i >= 1; i=i-1)
    begin: data_out_reg_stage
      mgc_generic_reg #(
        .width(62), 
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_data_out_reg (
        .d(data_out_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(data_out_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(62), 
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_data_out_reg_init (
      .d(data_out_t),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(data_out_reg[0])
    );
    assign data_out = data_out_reg[n_outreg-1];
  end
  else
  begin
    assign data_out = data_out_t;
  end
  endgenerate

endmodule



//------> ./rtl_stagemgc_rom_sync_regout_9_1024_64_1_0_0_1_0_1_0_0_0_1_60.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Sun Oct  6 01:48:34 2024
// ----------------------------------------------------------------------

// 
module stagemgc_rom_sync_regout_9_1024_64_1_0_0_1_0_1_0_0_0_1_60 (addr, data_out,
    clk, s_rst, a_rst, en
);
  input [9:0]addr ;
  output [63:0]data_out ;
  input clk ;
  input s_rst ;
  input a_rst ;
  input en ;


  // Constants for ROM dimensions
  parameter n_width    = 64;
  parameter n_size     = 1024;
  parameter n_numports = 1;
  parameter n_addr_w   = 10;
  parameter n_inreg    = 0;
  parameter n_outreg   = 1;
  wire [9:0] addr_f;

  // Build input address registers
  wire [9:0] addr_reg [n_inreg:0];
  genvar i;
  generate if (n_inreg > 0)
  begin
    for( i=n_inreg-1; i >= 1; i=i-1)
    begin: addr_reg_stage
      mgc_generic_reg #(
        .width(10), 
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_addr_reg (
        .d(addr_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(addr_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(10), 
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_addr_reg_init (
      .d(addr),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(addr_reg[0])
    );
    assign addr_f = addr_reg[n_inreg-1];
  end
  else
  begin
    assign addr_f = addr;
  end
  endgenerate

  // Declare storage for memory elements
  wire [63:0] mem [1023:0];

  // Declare output registers
  reg [63:0] data_out_t;

  // Initialize ROM contents
  assign mem[0] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  assign mem[1] = 64'b1000000000000000000000000000000000000000000000000000000000000000;
  assign mem[2] = 64'b0011111111100110101000001001111001100110011111110011101111001101;
  assign mem[3] = 64'b1011111111100110101000001001111001100110011111110011101111001101;
  assign mem[4] = 64'b0011111111101101100100000110101111001111001100101000110101000110;
  assign mem[5] = 64'b1011111111011000011111011110001010100110101011101010100101100011;
  assign mem[6] = 64'b0011111111011000011111011110001010100110101011101010100101100011;
  assign mem[7] = 64'b1011111111101101100100000110101111001111001100101000110101000110;
  assign mem[8] = 64'b0011111111101111011000101001011111001111111101110101110010110000;
  assign mem[9] = 64'b1011111111001000111110001011100000111100011010011010011000001011;
  assign mem[10] = 64'b0011111111100001110001110011101100111001101011100110100011001000;
  assign mem[11] = 64'b1011111111101010100110110110011000101001000011101010000110100011;
  assign mem[12] = 64'b0011111111101010100110110110011000101001000011101010000110100011;
  assign mem[13] = 64'b1011111111100001110001110011101100111001101011100110100011001000;
  assign mem[14] = 64'b0011111111001000111110001011100000111100011010011010011000001011;
  assign mem[15] = 64'b1011111111101111011000101001011111001111111101110101110010110000;
  assign mem[16] = 64'b0011111111101111110110001000110110100011110100010010010100100110;
  assign mem[17] = 64'b1011111110111001000101111010011010111100001010011011010000101100;
  assign mem[18] = 64'b0011111111100100010011001111001100100101000010010001110111010110;
  assign mem[19] = 64'b1011111111101000101111001000000001101011000101010001011101000001;
  assign mem[20] = 64'b0011111111101100001110001011001011110001100000001011110110110001;
  assign mem[21] = 64'b1011111111011110001010110101110100111000000001101111011000111011;
  assign mem[22] = 64'b0011111111010010100101000000011000101110110101011001111100000110;
  assign mem[23] = 64'b1011111111101110100111110100000101010110110001100010110111011010;
  assign mem[24] = 64'b0011111111101110100111110100000101010110110001100010110111011010;
  assign mem[25] = 64'b1011111111010010100101000000011000101110110101011001111100000110;
  assign mem[26] = 64'b0011111111011110001010110101110100111000000001101111011000111011;
  assign mem[27] = 64'b1011111111101100001110001011001011110001100000001011110110110001;
  assign mem[28] = 64'b0011111111101000101111001000000001101011000101010001011101000001;
  assign mem[29] = 64'b1011111111100100010011001111001100100101000010010001110111010110;
  assign mem[30] = 64'b0011111110111001000101111010011010111100001010011011010000101100;
  assign mem[31] = 64'b1011111111101111110110001000110110100011110100010010010100100110;
  assign mem[32] = 64'b0011111111101111111101100010000111100011011110010110110101111110;
  assign mem[33] = 64'b1011111110101001000111110110010111110001000011011101100000010100;
  assign mem[34] = 64'b0011111111100101011111010110100100110100100011001110110010100000;
  assign mem[35] = 64'b1011111111100111101101011101111100100010011010101010111110101111;
  assign mem[36] = 64'b0011111111101100111011010111101011110100001111001100011101110011;
  assign mem[37] = 64'b1011111111011011010111010001000000001001111000010101110011000000;
  assign mem[38] = 64'b0011111111010101100011111001101001110101101010110001111111011101;
  assign mem[39] = 64'b1011111111101110001000010010000100000100111101101000011011100101;
  assign mem[40] = 64'b0011111111101111000010100111111011111011100100100011000011010111;
  assign mem[41] = 64'b1011111111001111000110011111100101111011001000010101111100011011;
  assign mem[42] = 64'b0011111111100000011100111000011110011001001000101111111111101110;
  assign mem[43] = 64'b1011111111101011011100101000001101000101000110010110111000111110;
  assign mem[44] = 64'b0011111111101001101100111110000001000111111100111000011101000001;
  assign mem[45] = 64'b1011111111100011000011111111011111111100111000010111000000110101;
  assign mem[46] = 64'b0011111111000010110010000001000001101110100011100110000100111010;
  assign mem[47] = 64'b1011111111101111101001110101010101111111000010001010010100010111;
  assign mem[48] = 64'b0011111111101111101001110101010101111111000010001010010100010111;
  assign mem[49] = 64'b1011111111000010110010000001000001101110100011100110000100111010;
  assign mem[50] = 64'b0011111111100011000011111111011111111100111000010111000000110101;
  assign mem[51] = 64'b1011111111101001101100111110000001000111111100111000011101000001;
  assign mem[52] = 64'b0011111111101011011100101000001101000101000110010110111000111110;
  assign mem[53] = 64'b1011111111100000011100111000011110011001001000101111111111101110;
  assign mem[54] = 64'b0011111111001111000110011111100101111011001000010101111100011011;
  assign mem[55] = 64'b1011111111101111000010100111111011111011100100100011000011010111;
  assign mem[56] = 64'b0011111111101110001000010010000100000100111101101000011011100101;
  assign mem[57] = 64'b1011111111010101100011111001101001110101101010110001111111011101;
  assign mem[58] = 64'b0011111111011011010111010001000000001001111000010101110011000000;
  assign mem[59] = 64'b1011111111101100111011010111101011110100001111001100011101110011;
  assign mem[60] = 64'b0011111111100111101101011101111100100010011010101010111110101111;
  assign mem[61] = 64'b1011111111100101011111010110100100110100100011001110110010100000;
  assign mem[62] = 64'b0011111110101001000111110110010111110001000011011101100000010100;
  assign mem[63] = 64'b1011111111101111111101100010000111100011011110010110110101111110;
  assign mem[64] = 64'b0011111111101111111111011000100001100000100001001100110100001101;
  assign mem[65] = 64'b1011111110011001001000010101010111110111101000110110011001111110;
  assign mem[66] = 64'b0011111111100110000100001011011101010101000111010010110011011111;
  assign mem[67] = 64'b1011111111100111001011010000100000110111111011111111111110010110;
  assign mem[68] = 64'b0011111111101101010000010011010011010001010011011100100100111010;
  assign mem[69] = 64'b1011111111011001111011110111100101000011101010001110110110001010;
  assign mem[70] = 64'b0011111111010111000010001000010100110000111110100100010110011111;
  assign mem[71] = 64'b1011111111101101110110110001001110110110110011001100001000111100;
  assign mem[72] = 64'b0011111111101111001110001111001110101100011001001110010110001001;
  assign mem[73] = 64'b1011111111001100000010111000001001101010011111100100111101100011;
  assign mem[74] = 64'b0011111111100001000111101011001101010100000110110100101100100011;
  assign mem[75] = 64'b1011111111101011000010010000101001011000000101010000001000000000;
  assign mem[76] = 64'b0011111111101010001010011010011110100000010001100010011110000010;
  assign mem[77] = 64'b1011111111100010011011010000010101001100110111010001001011011111;
  assign mem[78] = 64'b0011111111000101111000100001010001000100100010110011111111000110;
  assign mem[79] = 64'b1011111111101111100001110110010011111010011100010100101110101001;
  assign mem[80] = 64'b0011111111101111110000100110010001110000111000011001111111010011;
  assign mem[81] = 64'b1011111110111111010101100100111001010110101010010111001100001110;
  assign mem[82] = 64'b0011111111100011101011111111101000101001001000000101000010111001;
  assign mem[83] = 64'b1011111111101001001110100010001001001001100100100110001111111011;
  assign mem[84] = 64'b0011111111101011110101111100000010101100011011111001010100101010;
  assign mem[85] = 64'b1011111111011111100010111010010011011011111110001001101010111010;
  assign mem[86] = 64'b0011111111010001000100011101001001100010101100011111011001110111;
  assign mem[87] = 64'b1011111111101110110101110100000011100111011010000100100101100011;
  assign mem[88] = 64'b0011111111101110011000101000100011101100010010001110000100010010;
  assign mem[89] = 64'b1011111111010100000100110101110010010100000101110110011000000001;
  assign mem[90] = 64'b0011111111011100110001100110111010011001001100011100010001011110;
  assign mem[91] = 64'b1011111111101100100101010100101100100001001101000001000111110101;
  assign mem[92] = 64'b0011111111101000001110110000111000001011111111111001011101101110;
  assign mem[93] = 64'b1011111111100100111001101100101010111011111000111110010111101001;
  assign mem[94] = 64'b0011111110110010110101010010000010010010110011100001100111110110;
  assign mem[95] = 64'b1011111111101111111010011100110110101101000000011000100000111010;
  assign mem[96] = 64'b0011111111101111111010011100110110101101000000011000100000111010;
  assign mem[97] = 64'b1011111110110010110101010010000010010010110011100001100111110110;
  assign mem[98] = 64'b0011111111100100111001101100101010111011111000111110010111101001;
  assign mem[99] = 64'b1011111111101000001110110000111000001011111111111001011101101110;
  assign mem[100] = 64'b0011111111101100100101010100101100100001001101000001000111110101;
  assign mem[101] = 64'b1011111111011100110001100110111010011001001100011100010001011110;
  assign mem[102] = 64'b0011111111010100000100110101110010010100000101110110011000000001;
  assign mem[103] = 64'b1011111111101110011000101000100011101100010010001110000100010010;
  assign mem[104] = 64'b0011111111101110110101110100000011100111011010000100100101100011;
  assign mem[105] = 64'b1011111111010001000100011101001001100010101100011111011001110111;
  assign mem[106] = 64'b0011111111011111100010111010010011011011111110001001101010111010;
  assign mem[107] = 64'b1011111111101011110101111100000010101100011011111001010100101010;
  assign mem[108] = 64'b0011111111101001001110100010001001001001100100100110001111111011;
  assign mem[109] = 64'b1011111111100011101011111111101000101001001000000101000010111001;
  assign mem[110] = 64'b0011111110111111010101100100111001010110101010010111001100001110;
  assign mem[111] = 64'b1011111111101111110000100110010001110000111000011001111111010011;
  assign mem[112] = 64'b0011111111101111100001110110010011111010011100010100101110101001;
  assign mem[113] = 64'b1011111111000101111000100001010001000100100010110011111111000110;
  assign mem[114] = 64'b0011111111100010011011010000010101001100110111010001001011011111;
  assign mem[115] = 64'b1011111111101010001010011010011110100000010001100010011110000010;
  assign mem[116] = 64'b0011111111101011000010010000101001011000000101010000001000000000;
  assign mem[117] = 64'b1011111111100001000111101011001101010100000110110100101100100011;
  assign mem[118] = 64'b0011111111001100000010111000001001101010011111100100111101100011;
  assign mem[119] = 64'b1011111111101111001110001111001110101100011001001110010110001001;
  assign mem[120] = 64'b0011111111101101110110110001001110110110110011001100001000111100;
  assign mem[121] = 64'b1011111111010111000010001000010100110000111110100100010110011111;
  assign mem[122] = 64'b0011111111011001111011110111100101000011101010001110110110001010;
  assign mem[123] = 64'b1011111111101101010000010011010011010001010011011100100100111010;
  assign mem[124] = 64'b0011111111100111001011010000100000110111111011111111111110010110;
  assign mem[125] = 64'b1011111111100110000100001011011101010101000111010010110011011111;
  assign mem[126] = 64'b0011111110011001001000010101010111110111101000110110011001111110;
  assign mem[127] = 64'b1011111111101111111111011000100001100000100001001100110100001101;
  assign mem[128] = 64'b0011111111101111111111110110001000010110100110111001001011011011;
  assign mem[129] = 64'b1011111110001001001000011101000111111100110111101100011110000100;
  assign mem[130] = 64'b0011111111100110010110010001100100100101111100000111100000111101;
  assign mem[131] = 64'b1011111111100110111001110100010001010100111010101010100010101111;
  assign mem[132] = 64'b0011111111101101011010010110000101110011110010011110011010001011;
  assign mem[133] = 64'b1011111111011001001101110010101001100011101111001001001111010111;
  assign mem[134] = 64'b0011111111010111110000111010100100110001000111011100110011100111;
  assign mem[135] = 64'b1011111111101101101101100101001001100010001110001010000010011011;
  assign mem[136] = 64'b0011111111101111010011100110000000111011000010110010111100101101;
  assign mem[137] = 64'b1011111111001010100000101010000000100101101100000000010001010001;
  assign mem[138] = 64'b0011111111100001011100110100110101100011110111101101101101001001;
  assign mem[139] = 64'b1011111111101010110100101011110010011110001000011101010100010001;
  assign mem[140] = 64'b0011111111101010011000110000100100011011000000101111101011100010;
  assign mem[141] = 64'b1011111111100010000110100111100110011001001100111110101101011001;
  assign mem[142] = 64'b0011111111000111011011011101100111011110010100001011111100110001;
  assign mem[143] = 64'b1011111111101111011101011001100110100011101000010010000001110111;
  assign mem[144] = 64'b0011111111101111110011100001010111111101011011011010011001111011;
  assign mem[145] = 64'b1011111110111100001101111000010111000111100111101100001011010101;
  assign mem[146] = 64'b0011111111100011111111101101100101010011010001010101011011010100;
  assign mem[147] = 64'b1011111111101000111110111100110010100011111011111001010000001101;
  assign mem[148] = 64'b0011111111101100000010001100010000100110011100100101010101001001;
  assign mem[149] = 64'b1011111111011110110111000001100101010010111011110111100011010110;
  assign mem[150] = 64'b0011111111010001110100110100010000111111010011001101101100111110;
  assign mem[151] = 64'b1011111111101110101110111101100011001000110111110000101101110100;
  assign mem[152] = 64'b0011111111101110100000010111101110101011010011001101000100001101;
  assign mem[153] = 64'b1011111111010011010101000001000011000010111000011000000101010010;
  assign mem[154] = 64'b0011111111011101011110010111011101011011100001101110001110001001;
  assign mem[155] = 64'b1011111111101100011001111000101100110100100010000111001110011011;
  assign mem[156] = 64'b0011111111101000011111000100000000001111101110100010111010111111;
  assign mem[157] = 64'b1011111111100100100110100100010010011011100110110000100100111001;
  assign mem[158] = 64'b0011111110110101111101101101000000001010100110101010010000011001;
  assign mem[159] = 64'b1011111111101111111000011100101011111100101111010101101100001001;
  assign mem[160] = 64'b0011111111101111111100001001010101100101100011100111000110101101;
  assign mem[161] = 64'b1011111110101111011001010110111001111001111110000010000011100000;
  assign mem[162] = 64'b0011111111100101001100101000001010010010101000110101010110010110;
  assign mem[163] = 64'b1011111111100111111110001110110011100011010101110001011101110001;
  assign mem[164] = 64'b0011111111101100110000011111000011110011111111001111110001011100;
  assign mem[165] = 64'b1011111111011100000100100100100111011000000000010001111011100111;
  assign mem[166] = 64'b0011111111010100110100011110001001000010011110001110011101101010;
  assign mem[167] = 64'b1011111111101110010000100110101001001011001010111100000101111110;
  assign mem[168] = 64'b0011111111101110111100010111100010100011111001000111001111000010;
  assign mem[169] = 64'b1011111111010000010011111011100000001110001101111111110110101110;
  assign mem[170] = 64'b0011111111100000000111001111110010000111010011000011111010110111;
  assign mem[171] = 64'b1011111111101011101001011010101001100111001101011001000011010010;
  assign mem[172] = 64'b0011111111101001011101110111111011110100110001111101011101000010;
  assign mem[173] = 64'b1011111111100011011000000101100010110001000001100101100111110011;
  assign mem[174] = 64'b0011111111000001001110011111000011001110110110101111010101110111;
  assign mem[175] = 64'b1011111111101111101101010111100101110001100101011101011101000001;
  assign mem[176] = 64'b0011111111101111100101111111100100100100110010010000100110011011;
  assign mem[177] = 64'b1011111111000100010101010111011010110001001010010011111001011010;
  assign mem[178] = 64'b0011111111100010101111101101101100100101111110101111001111101010;
  assign mem[179] = 64'b1011111111101001111011110100001111101111001010011010111110010100;
  assign mem[180] = 64'b0011111111101011001111100100110100111110111101010101011100010010;
  assign mem[181] = 64'b1011111111100000110010010111000001001101010111011000100110001111;
  assign mem[182] = 64'b0011111111001101100100110100111111100101010001010100001100010001;
  assign mem[183] = 64'b1011111111101111001000100101001011110111011101100011101011011010;
  assign mem[184] = 64'b0011111111101101111111101010111001100010001011011011111000101011;
  assign mem[185] = 64'b1011111111010110010011000111110111011101001111110010011111000110;
  assign mem[186] = 64'b0011111111011010101001101100100000101011011011010011111111001010;
  assign mem[187] = 64'b1011111111101101000101111110011101110100001111100011010111011100;
  assign mem[188] = 64'b0011111111100111011100011110011101011111000000110111001001100001;
  assign mem[189] = 64'b1011111111100101110001110111101110111110011001010000000110001100;
  assign mem[190] = 64'b0011111110100010110110000110010101110101100101000101010111001101;
  assign mem[191] = 64'b1011111111101111111110100111001011101111111111101111011101011101;
  assign mem[192] = 64'b0011111111101111111110100111001011101111111111101111011101011101;
  assign mem[193] = 64'b1011111110100010110110000110010101110101100101000101010111001101;
  assign mem[194] = 64'b0011111111100101110001110111101110111110011001010000000110001100;
  assign mem[195] = 64'b1011111111100111011100011110011101011111000000110111001001100001;
  assign mem[196] = 64'b0011111111101101000101111110011101110100001111100011010111011100;
  assign mem[197] = 64'b1011111111011010101001101100100000101011011011010011111111001010;
  assign mem[198] = 64'b0011111111010110010011000111110111011101001111110010011111000110;
  assign mem[199] = 64'b1011111111101101111111101010111001100010001011011011111000101011;
  assign mem[200] = 64'b0011111111101111001000100101001011110111011101100011101011011010;
  assign mem[201] = 64'b1011111111001101100100110100111111100101010001010100001100010001;
  assign mem[202] = 64'b0011111111100000110010010111000001001101010111011000100110001111;
  assign mem[203] = 64'b1011111111101011001111100100110100111110111101010101011100010010;
  assign mem[204] = 64'b0011111111101001111011110100001111101111001010011010111110010100;
  assign mem[205] = 64'b1011111111100010101111101101101100100101111110101111001111101010;
  assign mem[206] = 64'b0011111111000100010101010111011010110001001010010011111001011010;
  assign mem[207] = 64'b1011111111101111100101111111100100100100110010010000100110011011;
  assign mem[208] = 64'b0011111111101111101101010111100101110001100101011101011101000001;
  assign mem[209] = 64'b1011111111000001001110011111000011001110110110101111010101110111;
  assign mem[210] = 64'b0011111111100011011000000101100010110001000001100101100111110011;
  assign mem[211] = 64'b1011111111101001011101110111111011110100110001111101011101000010;
  assign mem[212] = 64'b0011111111101011101001011010101001100111001101011001000011010010;
  assign mem[213] = 64'b1011111111100000000111001111110010000111010011000011111010110111;
  assign mem[214] = 64'b0011111111010000010011111011100000001110001101111111110110101110;
  assign mem[215] = 64'b1011111111101110111100010111100010100011111001000111001111000010;
  assign mem[216] = 64'b0011111111101110010000100110101001001011001010111100000101111110;
  assign mem[217] = 64'b1011111111010100110100011110001001000010011110001110011101101010;
  assign mem[218] = 64'b0011111111011100000100100100100111011000000000010001111011100111;
  assign mem[219] = 64'b1011111111101100110000011111000011110011111111001111110001011100;
  assign mem[220] = 64'b0011111111100111111110001110110011100011010101110001011101110001;
  assign mem[221] = 64'b1011111111100101001100101000001010010010101000110101010110010110;
  assign mem[222] = 64'b0011111110101111011001010110111001111001111110000010000011100000;
  assign mem[223] = 64'b1011111111101111111100001001010101100101100011100111000110101101;
  assign mem[224] = 64'b0011111111101111111000011100101011111100101111010101101100001001;
  assign mem[225] = 64'b1011111110110101111101101101000000001010100110101010010000011001;
  assign mem[226] = 64'b0011111111100100100110100100010010011011100110110000100100111001;
  assign mem[227] = 64'b1011111111101000011111000100000000001111101110100010111010111111;
  assign mem[228] = 64'b0011111111101100011001111000101100110100100010000111001110011011;
  assign mem[229] = 64'b1011111111011101011110010111011101011011100001101110001110001001;
  assign mem[230] = 64'b0011111111010011010101000001000011000010111000011000000101010010;
  assign mem[231] = 64'b1011111111101110100000010111101110101011010011001101000100001101;
  assign mem[232] = 64'b0011111111101110101110111101100011001000110111110000101101110100;
  assign mem[233] = 64'b1011111111010001110100110100010000111111010011001101101100111110;
  assign mem[234] = 64'b0011111111011110110111000001100101010010111011110111100011010110;
  assign mem[235] = 64'b1011111111101100000010001100010000100110011100100101010101001001;
  assign mem[236] = 64'b0011111111101000111110111100110010100011111011111001010000001101;
  assign mem[237] = 64'b1011111111100011111111101101100101010011010001010101011011010100;
  assign mem[238] = 64'b0011111110111100001101111000010111000111100111101100001011010101;
  assign mem[239] = 64'b1011111111101111110011100001010111111101011011011010011001111011;
  assign mem[240] = 64'b0011111111101111011101011001100110100011101000010010000001110111;
  assign mem[241] = 64'b1011111111000111011011011101100111011110010100001011111100110001;
  assign mem[242] = 64'b0011111111100010000110100111100110011001001100111110101101011001;
  assign mem[243] = 64'b1011111111101010011000110000100100011011000000101111101011100010;
  assign mem[244] = 64'b0011111111101010110100101011110010011110001000011101010100010001;
  assign mem[245] = 64'b1011111111100001011100110100110101100011110111101101101101001001;
  assign mem[246] = 64'b0011111111001010100000101010000000100101101100000000010001010001;
  assign mem[247] = 64'b1011111111101111010011100110000000111011000010110010111100101101;
  assign mem[248] = 64'b0011111111101101101101100101001001100010001110001010000010011011;
  assign mem[249] = 64'b1011111111010111110000111010100100110001000111011100110011100111;
  assign mem[250] = 64'b0011111111011001001101110010101001100011101111001001001111010111;
  assign mem[251] = 64'b1011111111101101011010010110000101110011110010011110011010001011;
  assign mem[252] = 64'b0011111111100110111001110100010001010100111010101010100010101111;
  assign mem[253] = 64'b1011111111100110010110010001100100100101111100000111100000111101;
  assign mem[254] = 64'b0011111110001001001000011101000111111100110111101100011110000100;
  assign mem[255] = 64'b1011111111101111111111110110001000010110100110111001001011011011;
  assign mem[256] = 64'b0011111111101111111111111101100010000101100011101000101010010010;
  assign mem[257] = 64'b1011111101111001001000011111000011111110011001110000000001110001;
  assign mem[258] = 64'b0011111111100110011111001111011110000100100100011010111100010000;
  assign mem[259] = 64'b1011111111100110110001000000110101110011110000011000001001110101;
  assign mem[260] = 64'b0011111111101101011111010000101100000010101110001110110011111001;
  assign mem[261] = 64'b1011111111011000110110101010010100101110110010001010010010110000;
  assign mem[262] = 64'b0011111111011000001000001110001110110000010011101010101011000100;
  assign mem[263] = 64'b1011111111101101101000111000001110101001011001101000100110001000;
  assign mem[264] = 64'b0011111111101111010110001010001010110001011110001001111010000100;
  assign mem[265] = 64'b1011111111001001101111011100101111110010110111000100001101100110;
  assign mem[266] = 64'b0011111111100001100111010101101000001001111100101011100110111000;
  assign mem[267] = 64'b1011111111101010101101110011001001011001000101101100000011010100;
  assign mem[268] = 64'b0011111111101010011111110101100001010010100111111110011010011101;
  assign mem[269] = 64'b1011111111100001111100001111000010001011101111001000011000011011;
  assign mem[270] = 64'b0011111111001000001100110110011011101000100111000110010011000110;
  assign mem[271] = 64'b1011111111101111011011000011111101111101111101011011101110110111;
  assign mem[272] = 64'b0011111111101111110100110111100100010100001000100000101110000100;
  assign mem[273] = 64'b1011111110111010101001111011011100100100010010010101110000000011;
  assign mem[274] = 64'b0011111111100100001001011111111100010111100011100110101110110001;
  assign mem[275] = 64'b1011111111101000110111000100010100110011000101101001100011001100;
  assign mem[276] = 64'b0011111111101100001000001101111000111111101010010111000110110000;
  assign mem[277] = 64'b1011111111011110100000111110000011101010111110000101000100010100;
  assign mem[278] = 64'b0011111111010010001100111011101110101011110000111011101101110001;
  assign mem[279] = 64'b1011111111101110101011011011001011101000111001111010100010001110;
  assign mem[280] = 64'b0011111111101110100100001000010000110110000111011111011111110010;
  assign mem[281] = 64'b1011111111010010111101000010001011011010111011000000001110000111;
  assign mem[282] = 64'b0011111111011101110100101000111100010100100000011100110001011000;
  assign mem[283] = 64'b1011111111101100010100000100001000000001001010110110100100000111;
  assign mem[284] = 64'b0011111111101000100111000111111010011010010011011101010010101010;
  assign mem[285] = 64'b1011111111100100011100111011010100011011100110000111001101000111;
  assign mem[286] = 64'b0011111110110111100001110101100001101010010111010101101100100001;
  assign mem[287] = 64'b1011111111101111110111010101001110011111111100011111010001010110;
  assign mem[288] = 64'b0011111111101111111100111000001100001111100011010101011101011100;
  assign mem[289] = 64'b1011111110101100010000101000110100010010110000001101011111100011;
  assign mem[290] = 64'b0011111111100101010110000001000000111000100101110101000100110111;
  assign mem[291] = 64'b1011111111100111110101111000001101101100110000110011110110110010;
  assign mem[292] = 64'b0011111111101100110101111101100110001001100010110011001011110110;
  assign mem[293] = 64'b1011111111011011101101111100111100100011000001001011110100000001;
  assign mem[294] = 64'b0011111111010101001100001101100010000000101011110011110000100100;
  assign mem[295] = 64'b1011111111101110001100011110101011101000011100001100111000100101;
  assign mem[296] = 64'b0011111111101110111111100010001000001100000010111001010111101100;
  assign mem[297] = 64'b1011111111001111110111001101110000011010110111111110110111111001;
  assign mem[298] = 64'b0011111111100000010010000101011000100110101011100010001000011010;
  assign mem[299] = 64'b1011111111101011100011000011100011010010011101010000010011101001;
  assign mem[300] = 64'b0011111111101001100101011100111100101110110110000000110100100010;
  assign mem[301] = 64'b1011111111100011001110000100000000001101000011001000111001010111;
  assign mem[302] = 64'b0011111111000010000000010001011011010100111011000111101111001111;
  assign mem[303] = 64'b1011111111101111101011101000111010001110010001101100111110111011;
  assign mem[304] = 64'b0011111111101111100111111100111001010101101011011011001011001000;
  assign mem[305] = 64'b1011111111000011100011101101101110110000110011011000110100010100;
  assign mem[306] = 64'b0011111111100010111001111000000011100011111010001110101000010111;
  assign mem[307] = 64'b1011111111101001110100011011000111110101111010101000000011010101;
  assign mem[308] = 64'b0011111111101011010110001000100111111110100100100001010000000101;
  assign mem[309] = 64'b1011111111100000100111101001000001110100000101111100010111100001;
  assign mem[310] = 64'b0011111111001110010101101100101000011110000100000001101000011011;
  assign mem[311] = 64'b1011111111101111000101101000111101010011111101110010000001011101;
  assign mem[312] = 64'b0011111111101110000100000000110011001010001010011000000010101100;
  assign mem[313] = 64'b1011111111010101111011100010011100110111100111101010011010010011;
  assign mem[314] = 64'b0011111111011011000000100000110101101100011111110100000000001001;
  assign mem[315] = 64'b1011111111101101000000101101010011111110101100101011110110010010;
  assign mem[316] = 64'b0011111111100111100101000000000001010111010011110101010111100101;
  assign mem[317] = 64'b1011111111100101101000101000110100101010010111010111001001010000;
  assign mem[318] = 64'b0011111110100101111111000000000011010010100100001100110101000011;
  assign mem[319] = 64'b1011111111101111111110000111000111011010110110111000000111011111;
  assign mem[320] = 64'b0011111111101111111111000010010100011101111100011101001111111000;
  assign mem[321] = 64'b1011111110011111011010010011011100110001110100011100111100000001;
  assign mem[322] = 64'b0011111111100101111011000011010010010101100000110111000001110100;
  assign mem[323] = 64'b1011111111100111010011111001010010001101101010001101001010001101;
  assign mem[324] = 64'b0011111111101101001011001011001000100000111000001110111110011111;
  assign mem[325] = 64'b1011111111011010010010110100000100100111110111101010000111100101;
  assign mem[326] = 64'b0011111111010110101010101001110101111101110001110111111000010111;
  assign mem[327] = 64'b1011111111101101111011010000010111110111110111100100011111011010;
  assign mem[328] = 64'b0011111111101111001011011100100111001001000010001001101010011101;
  assign mem[329] = 64'b1011111111001100110011111000110010110011000100101011001010000110;
  assign mem[330] = 64'b0011111111100000111101000010011010111011001010101000111001111110;
  assign mem[331] = 64'b1011111111101011001000111100110101000111000000000001001110110100;
  assign mem[332] = 64'b0011111111101010000011001001010111101010101110101111100100110111;
  assign mem[333] = 64'b1011111111100010100101100000011100100111011000101001110010101000;
  assign mem[334] = 64'b0011111111000101000110111101111110000101100101111100010111110010;
  assign mem[335] = 64'b1011111111101111100011111101010111111111101011100100000111011011;
  assign mem[336] = 64'b0011111111101111101111000001011000010111111001000100000110000110;
  assign mem[337] = 64'b1011111111000000011100101010000001000111101110101000001100011101;
  assign mem[338] = 64'b0011111111100011100010000100000110000101110111111110101100100010;
  assign mem[339] = 64'b1011111111101001010110001110111111100100100011100110110111010111;
  assign mem[340] = 64'b0011111111101011101111101101011111000100100100111000000011101010;
  assign mem[341] = 64'b1011111111011111111000101111011001001011111001110001001000010000;
  assign mem[342] = 64'b0011111111010000101100001101100111001111110110111101101110010000;
  assign mem[343] = 64'b1011111111101110111001001000001011100010010110101001110110111100;
  assign mem[344] = 64'b0011111111101110010100101001111100000100011100101001111111111100;
  assign mem[345] = 64'b1011111111010100011100101011100010100101010101110001000001010100;
  assign mem[346] = 64'b0011111111011100011011000111111101001001100101110000000000001011;
  assign mem[347] = 64'b1011111111101100101010111100000101101001101000001011100100000000;
  assign mem[348] = 64'b0011111111101000000110100001101100110011101101010111101011001100;
  assign mem[349] = 64'b1011111111100101000011001100000010011111010110011010000010011011;
  assign mem[350] = 64'b0011111110110001010001000000000100110100110101110000100110110011;
  assign mem[351] = 64'b1011111111101111111011010101100011101100101101100111001111000100;
  assign mem[352] = 64'b0011111111101111111001011111001110101111001011100011100101000000;
  assign mem[353] = 64'b1011111110110100011001100001000101111001001001110010000010010110;
  assign mem[354] = 64'b0011111111100100110000001010000101000101111011000000000000000100;
  assign mem[355] = 64'b1011111111101000010110111100010100011010111010010101100011001100;
  assign mem[356] = 64'b0011111111101100011111101000111001010010001000110011110011110011;
  assign mem[357] = 64'b1011111111011101001000000001011011101000111010011101101101011011;
  assign mem[358] = 64'b0011111111010011101100111100111011111010000001000001010010110111;
  assign mem[359] = 64'b1011111111101110011100100010011111011011011010101001011101000100;
  assign mem[360] = 64'b0011111111101110110010011011001011010011110000111011111110000100;
  assign mem[361] = 64'b1011111111010001011100101010000011010111011101100101000101110111;
  assign mem[362] = 64'b0011111111011111001101000000010110010110001111111101000001100111;
  assign mem[363] = 64'b1011111111101011111100000110010011100001010100110111011111011101;
  assign mem[364] = 64'b0011111111101001000110110001011001101111110101001001110110100010;
  assign mem[365] = 64'b1011111111100011110101111000001000111000110001011000001101000100;
  assign mem[366] = 64'b0011111110111101110001110000111011001011101011101001111111001001;
  assign mem[367] = 64'b1011111111101111110010000110010001101100111111101011011100100001;
  assign mem[368] = 64'b0011111111101111011111101010011000101001111001100011110101101110;
  assign mem[369] = 64'b1011111111000110101010000001001100000100111101100100101010110010;
  assign mem[370] = 64'b0011111111100010010000111101010111111011100110001010110000011111;
  assign mem[371] = 64'b1011111111101010010001100111100011001000000100011001101011001000;
  assign mem[372] = 64'b0011111111101010111011100000010010110100001111000001010001110100;
  assign mem[373] = 64'b1011111111100001010010010001010110101111001100110110110011101011;
  assign mem[374] = 64'b0011111111001011010001110011001011101111001111010110011100100010;
  assign mem[375] = 64'b1011111111101111010000111101000010000101111111111001001011011101;
  assign mem[376] = 64'b0011111111101101110010001101011111001011010000010000001001100000;
  assign mem[377] = 64'b1011111111010111011001100011010000001111001001000001100011110110;
  assign mem[378] = 64'b0011111111011001100100110111000101100001010000011011110111111111;
  assign mem[379] = 64'b1011111111101101010101010110111101010010111010010011111010110001;
  assign mem[380] = 64'b0011111111100111000010100100001010110011000101110110110101111010;
  assign mem[381] = 64'b1011111111100110001101010000001110100011000111000001101111101001;
  assign mem[382] = 64'b0011111110010010110110010011011010111011111000110000111011111101;
  assign mem[383] = 64'b1011111111101111111111101001110010110100010010110101000110100001;
  assign mem[384] = 64'b0011111111101111111111101001110010110100010010110101000110100001;
  assign mem[385] = 64'b1011111110010010110110010011011010111011111000110000111011111101;
  assign mem[386] = 64'b0011111111100110001101010000001110100011000111000001101111101001;
  assign mem[387] = 64'b1011111111100111000010100100001010110011000101110110110101111010;
  assign mem[388] = 64'b0011111111101101010101010110111101010010111010010011111010110001;
  assign mem[389] = 64'b1011111111011001100100110111000101100001010000011011110111111111;
  assign mem[390] = 64'b0011111111010111011001100011010000001111001001000001100011110110;
  assign mem[391] = 64'b1011111111101101110010001101011111001011010000010000001001100000;
  assign mem[392] = 64'b0011111111101111010000111101000010000101111111111001001011011101;
  assign mem[393] = 64'b1011111111001011010001110011001011101111001111010110011100100010;
  assign mem[394] = 64'b0011111111100001010010010001010110101111001100110110110011101011;
  assign mem[395] = 64'b1011111111101010111011100000010010110100001111000001010001110100;
  assign mem[396] = 64'b0011111111101010010001100111100011001000000100011001101011001000;
  assign mem[397] = 64'b1011111111100010010000111101010111111011100110001010110000011111;
  assign mem[398] = 64'b0011111111000110101010000001001100000100111101100100101010110010;
  assign mem[399] = 64'b1011111111101111011111101010011000101001111001100011110101101110;
  assign mem[400] = 64'b0011111111101111110010000110010001101100111111101011011100100001;
  assign mem[401] = 64'b1011111110111101110001110000111011001011101011101001111111001001;
  assign mem[402] = 64'b0011111111100011110101111000001000111000110001011000001101000100;
  assign mem[403] = 64'b1011111111101001000110110001011001101111110101001001110110100010;
  assign mem[404] = 64'b0011111111101011111100000110010011100001010100110111011111011101;
  assign mem[405] = 64'b1011111111011111001101000000010110010110001111111101000001100111;
  assign mem[406] = 64'b0011111111010001011100101010000011010111011101100101000101110111;
  assign mem[407] = 64'b1011111111101110110010011011001011010011110000111011111110000100;
  assign mem[408] = 64'b0011111111101110011100100010011111011011011010101001011101000100;
  assign mem[409] = 64'b1011111111010011101100111100111011111010000001000001010010110111;
  assign mem[410] = 64'b0011111111011101001000000001011011101000111010011101101101011011;
  assign mem[411] = 64'b1011111111101100011111101000111001010010001000110011110011110011;
  assign mem[412] = 64'b0011111111101000010110111100010100011010111010010101100011001100;
  assign mem[413] = 64'b1011111111100100110000001010000101000101111011000000000000000100;
  assign mem[414] = 64'b0011111110110100011001100001000101111001001001110010000010010110;
  assign mem[415] = 64'b1011111111101111111001011111001110101111001011100011100101000000;
  assign mem[416] = 64'b0011111111101111111011010101100011101100101101100111001111000100;
  assign mem[417] = 64'b1011111110110001010001000000000100110100110101110000100110110011;
  assign mem[418] = 64'b0011111111100101000011001100000010011111010110011010000010011011;
  assign mem[419] = 64'b1011111111101000000110100001101100110011101101010111101011001100;
  assign mem[420] = 64'b0011111111101100101010111100000101101001101000001011100100000000;
  assign mem[421] = 64'b1011111111011100011011000111111101001001100101110000000000001011;
  assign mem[422] = 64'b0011111111010100011100101011100010100101010101110001000001010100;
  assign mem[423] = 64'b1011111111101110010100101001111100000100011100101001111111111100;
  assign mem[424] = 64'b0011111111101110111001001000001011100010010110101001110110111100;
  assign mem[425] = 64'b1011111111010000101100001101100111001111110110111101101110010000;
  assign mem[426] = 64'b0011111111011111111000101111011001001011111001110001001000010000;
  assign mem[427] = 64'b1011111111101011101111101101011111000100100100111000000011101010;
  assign mem[428] = 64'b0011111111101001010110001110111111100100100011100110110111010111;
  assign mem[429] = 64'b1011111111100011100010000100000110000101110111111110101100100010;
  assign mem[430] = 64'b0011111111000000011100101010000001000111101110101000001100011101;
  assign mem[431] = 64'b1011111111101111101111000001011000010111111001000100000110000110;
  assign mem[432] = 64'b0011111111101111100011111101010111111111101011100100000111011011;
  assign mem[433] = 64'b1011111111000101000110111101111110000101100101111100010111110010;
  assign mem[434] = 64'b0011111111100010100101100000011100100111011000101001110010101000;
  assign mem[435] = 64'b1011111111101010000011001001010111101010101110101111100100110111;
  assign mem[436] = 64'b0011111111101011001000111100110101000111000000000001001110110100;
  assign mem[437] = 64'b1011111111100000111101000010011010111011001010101000111001111110;
  assign mem[438] = 64'b0011111111001100110011111000110010110011000100101011001010000110;
  assign mem[439] = 64'b1011111111101111001011011100100111001001000010001001101010011101;
  assign mem[440] = 64'b0011111111101101111011010000010111110111110111100100011111011010;
  assign mem[441] = 64'b1011111111010110101010101001110101111101110001110111111000010111;
  assign mem[442] = 64'b0011111111011010010010110100000100100111110111101010000111100101;
  assign mem[443] = 64'b1011111111101101001011001011001000100000111000001110111110011111;
  assign mem[444] = 64'b0011111111100111010011111001010010001101101010001101001010001101;
  assign mem[445] = 64'b1011111111100101111011000011010010010101100000110111000001110100;
  assign mem[446] = 64'b0011111110011111011010010011011100110001110100011100111100000001;
  assign mem[447] = 64'b1011111111101111111111000010010100011101111100011101001111111000;
  assign mem[448] = 64'b0011111111101111111110000111000111011010110110111000000111011111;
  assign mem[449] = 64'b1011111110100101111111000000000011010010100100001100110101000011;
  assign mem[450] = 64'b0011111111100101101000101000110100101010010111010111001001010000;
  assign mem[451] = 64'b1011111111100111100101000000000001010111010011110101010111100101;
  assign mem[452] = 64'b0011111111101101000000101101010011111110101100101011110110010010;
  assign mem[453] = 64'b1011111111011011000000100000110101101100011111110100000000001001;
  assign mem[454] = 64'b0011111111010101111011100010011100110111100111101010011010010011;
  assign mem[455] = 64'b1011111111101110000100000000110011001010001010011000000010101100;
  assign mem[456] = 64'b0011111111101111000101101000111101010011111101110010000001011101;
  assign mem[457] = 64'b1011111111001110010101101100101000011110000100000001101000011011;
  assign mem[458] = 64'b0011111111100000100111101001000001110100000101111100010111100001;
  assign mem[459] = 64'b1011111111101011010110001000100111111110100100100001010000000101;
  assign mem[460] = 64'b0011111111101001110100011011000111110101111010101000000011010101;
  assign mem[461] = 64'b1011111111100010111001111000000011100011111010001110101000010111;
  assign mem[462] = 64'b0011111111000011100011101101101110110000110011011000110100010100;
  assign mem[463] = 64'b1011111111101111100111111100111001010101101011011011001011001000;
  assign mem[464] = 64'b0011111111101111101011101000111010001110010001101100111110111011;
  assign mem[465] = 64'b1011111111000010000000010001011011010100111011000111101111001111;
  assign mem[466] = 64'b0011111111100011001110000100000000001101000011001000111001010111;
  assign mem[467] = 64'b1011111111101001100101011100111100101110110110000000110100100010;
  assign mem[468] = 64'b0011111111101011100011000011100011010010011101010000010011101001;
  assign mem[469] = 64'b1011111111100000010010000101011000100110101011100010001000011010;
  assign mem[470] = 64'b0011111111001111110111001101110000011010110111111110110111111001;
  assign mem[471] = 64'b1011111111101110111111100010001000001100000010111001010111101100;
  assign mem[472] = 64'b0011111111101110001100011110101011101000011100001100111000100101;
  assign mem[473] = 64'b1011111111010101001100001101100010000000101011110011110000100100;
  assign mem[474] = 64'b0011111111011011101101111100111100100011000001001011110100000001;
  assign mem[475] = 64'b1011111111101100110101111101100110001001100010110011001011110110;
  assign mem[476] = 64'b0011111111100111110101111000001101101100110000110011110110110010;
  assign mem[477] = 64'b1011111111100101010110000001000000111000100101110101000100110111;
  assign mem[478] = 64'b0011111110101100010000101000110100010010110000001101011111100011;
  assign mem[479] = 64'b1011111111101111111100111000001100001111100011010101011101011100;
  assign mem[480] = 64'b0011111111101111110111010101001110011111111100011111010001010110;
  assign mem[481] = 64'b1011111110110111100001110101100001101010010111010101101100100001;
  assign mem[482] = 64'b0011111111100100011100111011010100011011100110000111001101000111;
  assign mem[483] = 64'b1011111111101000100111000111111010011010010011011101010010101010;
  assign mem[484] = 64'b0011111111101100010100000100001000000001001010110110100100000111;
  assign mem[485] = 64'b1011111111011101110100101000111100010100100000011100110001011000;
  assign mem[486] = 64'b0011111111010010111101000010001011011010111011000000001110000111;
  assign mem[487] = 64'b1011111111101110100100001000010000110110000111011111011111110010;
  assign mem[488] = 64'b0011111111101110101011011011001011101000111001111010100010001110;
  assign mem[489] = 64'b1011111111010010001100111011101110101011110000111011101101110001;
  assign mem[490] = 64'b0011111111011110100000111110000011101010111110000101000100010100;
  assign mem[491] = 64'b1011111111101100001000001101111000111111101010010111000110110000;
  assign mem[492] = 64'b0011111111101000110111000100010100110011000101101001100011001100;
  assign mem[493] = 64'b1011111111100100001001011111111100010111100011100110101110110001;
  assign mem[494] = 64'b0011111110111010101001111011011100100100010010010101110000000011;
  assign mem[495] = 64'b1011111111101111110100110111100100010100001000100000101110000100;
  assign mem[496] = 64'b0011111111101111011011000011111101111101111101011011101110110111;
  assign mem[497] = 64'b1011111111001000001100110110011011101000100111000110010011000110;
  assign mem[498] = 64'b0011111111100001111100001111000010001011101111001000011000011011;
  assign mem[499] = 64'b1011111111101010011111110101100001010010100111111110011010011101;
  assign mem[500] = 64'b0011111111101010101101110011001001011001000101101100000011010100;
  assign mem[501] = 64'b1011111111100001100111010101101000001001111100101011100110111000;
  assign mem[502] = 64'b0011111111001001101111011100101111110010110111000100001101100110;
  assign mem[503] = 64'b1011111111101111010110001010001010110001011110001001111010000100;
  assign mem[504] = 64'b0011111111101101101000111000001110101001011001101000100110001000;
  assign mem[505] = 64'b1011111111011000001000001110001110110000010011101010101011000100;
  assign mem[506] = 64'b0011111111011000110110101010010100101110110010001010010010110000;
  assign mem[507] = 64'b1011111111101101011111010000101100000010101110001110110011111001;
  assign mem[508] = 64'b0011111111100110110001000000110101110011110000011000001001110101;
  assign mem[509] = 64'b1011111111100110011111001111011110000100100100011010111100010000;
  assign mem[510] = 64'b0011111101111001001000011111000011111110011001110000000001110001;
  assign mem[511] = 64'b1011111111101111111111111101100010000101100011101000101010010010;
  assign mem[512] = 64'b0011111111101111111111111111011000100001011000100001110100000010;
  assign mem[513] = 64'b1011111101101001001000011111100010111110110011001010010010111010;
  assign mem[514] = 64'b0011111111100110100011101101000111101010101000011001110001110001;
  assign mem[515] = 64'b1011111111100110101100100101110011101101001011111110001010011100;
  assign mem[516] = 64'b0011111111101101100001101100010010000100010001011010010001001111;
  assign mem[517] = 64'b1011111111011000101011000100101110000110110101011110110101000100;
  assign mem[518] = 64'b0011111111011000010011110110101010101010111100111001000000111111;
  assign mem[519] = 64'b1011111111101101100110100000000011011101100010110011110101000110;
  assign mem[520] = 64'b0011111111101111010111011010011011101101010000110110100001011101;
  assign mem[521] = 64'b1011111111001001010110110100100111101001101101100010101011111010;
  assign mem[522] = 64'b0011111111100001101100100101000000010111000100110111001110111111;
  assign mem[523] = 64'b1011111111101010101010010101010001111010001011001011100110001110;
  assign mem[524] = 64'b0011111111101010100011010110011101101110010101000101101011010010;
  assign mem[525] = 64'b1011111111100001110111000001101101100100110111000100100001110010;
  assign mem[526] = 64'b0011111111001000100101100001011100100111110001000001100000000100;
  assign mem[527] = 64'b1011111111101111011001110111010101010110100010000011110011101110;
  assign mem[528] = 64'b0011111111101111110101100000110100101101101001110101110010011110;
  assign mem[529] = 64'b1011111110111001110111111011011011101011001001001010100001011100;
  assign mem[530] = 64'b0011111111100100001110010111111101011011001010100100001110000000;
  assign mem[531] = 64'b1011111111101000110011000110101001110101000110000100011001010101;
  assign mem[532] = 64'b0011111111101100001011001101000101001001001100011110001111110001;
  assign mem[533] = 64'b1011111111011110010101111010100001101101001111001101100000100101;
  assign mem[534] = 64'b0011111111010010011000111110011010011001010101010101010010111010;
  assign mem[535] = 64'b1011111111101110101001101000001110010011111001100101100000000000;
  assign mem[536] = 64'b0011111111101110100101111110110000110110000000010110101100110000;
  assign mem[537] = 64'b1011111111010010110001000001101001001110100101010100010100100000;
  assign mem[538] = 64'b0011111111011101111111101111111101100110101010010100000111011110;
  assign mem[539] = 64'b1011111111101100010001001000001100110001010000011100000000000100;
  assign mem[540] = 64'b0011111111101000101011001000011100011110110111100001110110001000;
  assign mem[541] = 64'b1011111111100100011000000101101001101001001010110011001010100010;
  assign mem[542] = 64'b0011111110111000010011111000011100010010110000010011000010100001;
  assign mem[543] = 64'b1011111111101111110110101111101001110101000101000101001110001100;
  assign mem[544] = 64'b0011111111101111111101001101110001010100101100011011111011010011;
  assign mem[545] = 64'b1011111110101010101100010000000110111101010111111000001100010111;
  assign mem[546] = 64'b0011111111100101011010101100001101010001100101110110010010011111;
  assign mem[547] = 64'b1011111111100111110001101011100010011100111000101101001100110011;
  assign mem[548] = 64'b0011111111101100111000101011001100100111100110011010000001100000;
  assign mem[549] = 64'b1011111111011011100010100111100000010100111111010101011010010011;
  assign mem[550] = 64'b0011111111010101011000000100000000010010111101000110011110110100;
  assign mem[551] = 64'b1011111111101110001010011000111101000100001110010001100101111010;
  assign mem[552] = 64'b0011111111101111000001000101101000010100110011110111001110001100;
  assign mem[553] = 64'b1011111111001111011110110111010010000000101111010011100000000010;
  assign mem[554] = 64'b0011111111100000010111011111001111101100001100011011100010110111;
  assign mem[555] = 64'b1011111111101011011111110110011010000110111001111001001011101001;
  assign mem[556] = 64'b0011111111101001101001001101111110100100001010110000011010110010;
  assign mem[557] = 64'b1011111111100011001001000010000111101100010010011010011000011111;
  assign mem[558] = 64'b0011111111000010011001001001100101001101111111010011010000001001;
  assign mem[559] = 64'b1011111111101111101010101111101111001011000011001111110111011100;
  assign mem[560] = 64'b0011111111101111101000111001101110101100011110100001011110010001;
  assign mem[561] = 64'b1011111111000011001010110111101111111001010001010001011010100111;
  assign mem[562] = 64'b0011111111100010111110111100001001001011010001000001000000010101;
  assign mem[563] = 64'b1011111111101001110000101101000100010000111100000111010111000010;
  assign mem[564] = 64'b0011111111101011011001011000111100010100111111011011110001000111;
  assign mem[565] = 64'b1011111111100000100010010001000100100000001100101011000010001100;
  assign mem[566] = 64'b0011111111001110101110000110101101000110001011011110001101001000;
  assign mem[567] = 64'b1011111111101111000100001001000010111100100010011000111101011111;
  assign mem[568] = 64'b0011111111101110000110001010000000101111110111000110011011011001;
  assign mem[569] = 64'b1011111111010101101111101110011110001011100111011011001110110110;
  assign mem[570] = 64'b0011111111011011001011111001011100011101101100110001100101110010;
  assign mem[571] = 64'b1011111111101100111110000011000011101000110011100100011001111011;
  assign mem[572] = 64'b0011111111100111101001001111011100000111101111111001011111010010;
  assign mem[573] = 64'b1011111111100101100100000000000111010101111101110010001111011111;
  assign mem[574] = 64'b0011111110100111100011011011101010100101100001110100011010000110;
  assign mem[575] = 64'b1011111111101111111101110101001110111011000110111001000101100100;
  assign mem[576] = 64'b0011111111101111111111001110000010011100111000101010011001111001;
  assign mem[577] = 64'b1011111110011100010001010100111101001100111001010011101100011101;
  assign mem[578] = 64'b0011111111100101111111100111110010111101111001010110101000010000;
  assign mem[579] = 64'b1011111111100111001111100101010110001110000001111001100101000010;
  assign mem[580] = 64'b0011111111101101001101101111110001111011110010111111101111011100;
  assign mem[581] = 64'b1011111111011010000111010110010101000011101101010000101011000000;
  assign mem[582] = 64'b0011111111010110110110011001100001100011100010100000110010110110;
  assign mem[583] = 64'b1011111111101101111001000001011000001111011011011000110110000001;
  assign mem[584] = 64'b0011111111101111001100110110100001011010001110101010111011110000;
  assign mem[585] = 64'b1011111111001100011011011001000001010011010111010111010011011101;
  assign mem[586] = 64'b0011111111100001000010010111001001001000110100001010100101010111;
  assign mem[587] = 64'b1011111111101011000101100111010000101010010011001010001011110101;
  assign mem[588] = 64'b0011111111101010000110110010011011010010110000001010011101011110;
  assign mem[589] = 64'b1011111111100010100000011000101111101111010011010011110010111010;
  assign mem[590] = 64'b0011111111000101011111110000000010000110010101001100101111011110;
  assign mem[591] = 64'b1011111111101111100010111010011100110111110010110100101101111000;
  assign mem[592] = 64'b0011111111101111101111110100011100001111000010101000110110001000;
  assign mem[593] = 64'b1011111111000000000011101110100010101101011011111011100001011011;
  assign mem[594] = 64'b0011111111100011100111000010001111100011110101100011000000101001;
  assign mem[595] = 64'b1011111111101001010010011001000011100011101011000100101001101100;
  assign mem[596] = 64'b0011111111101011110010110101010011001011000011010010001100100111;
  assign mem[597] = 64'b1011111111011111101101110101011101011100001001001101001011011110;
  assign mem[598] = 64'b0011111111010000111000010101101101001110000101110100100111001110;
  assign mem[599] = 64'b1011111111101110110111011110101101101010000001111000011001010001;
  assign mem[600] = 64'b0011111111101110010110101001110101010101000001000110011111010011;
  assign mem[601] = 64'b1011111111010100010000110001000011011100100010010011011011110000;
  assign mem[602] = 64'b0011111111011100100110010111111111000011100001100101001110001001;
  assign mem[603] = 64'b1011111111101100101000001000111100011001101110011100010001001001;
  assign mem[604] = 64'b0011111111101000001010101001110000010011111101010100010111111111;
  assign mem[605] = 64'b1011111111100100111110011100110000100101110011001010010010000110;
  assign mem[606] = 64'b0011111110110010000011001001011001110100111011010100010001001101;
  assign mem[607] = 64'b1011111111101111111010111001110100100101001100000100000100001111;
  assign mem[608] = 64'b0011111111101111111001111110101010000101010010000010110101100000;
  assign mem[609] = 64'b1011111110110011100111011001111100010010110001011010001010011001;
  assign mem[610] = 64'b0011111111100100110100111011110001101101010110001001111101111111;
  assign mem[611] = 64'b1011111111101000010010110111000100010001101011111000001111111010;
  assign mem[612] = 64'b0011111111101100100010011111010110000111000000101001110000010011;
  assign mem[613] = 64'b1011111111011100111100110100101110101110111000011100110100100001;
  assign mem[614] = 64'b0011111111010011111000111001101111101001011011101100001001110001;
  assign mem[615] = 64'b1011111111101110011010100110000111000101010111010101001110100111;
  assign mem[616] = 64'b0011111111101110110100001000001101011110100110011001000000001001;
  assign mem[617] = 64'b1011111111010001010000100011111011101111110001101001001101111000;
  assign mem[618] = 64'b0011111111011111010111111101111011100110010101101100110110100011;
  assign mem[619] = 64'b1011111111101011111001000001101101100001000100010101010011000001;
  assign mem[620] = 64'b0011111111101001001010101010010000011111110001011010100000010101;
  assign mem[621] = 64'b1011111111100011110000111100010001001001100000011100010100011000;
  assign mem[622] = 64'b0011111110111110100011101011011111111101111001001010101000111111;
  assign mem[623] = 64'b1011111111101111110001010110111000111011011111011001101011110110;
  assign mem[624] = 64'b0011111111101111100000110000111101001010010000001100011000001100;
  assign mem[625] = 64'b1011111111000110010001010001101010000011000111011000001100001101;
  assign mem[626] = 64'b0011111111100010010110000111001101001100101110110111000100010000;
  assign mem[627] = 64'b1011111111101010001110000001100001001010010110010011101111000110;
  assign mem[628] = 64'b0011111111101010111110111000111111011000100111110101011110110110;
  assign mem[629] = 64'b1011111111100001001100111110100111001111111011100010010101001111;
  assign mem[630] = 64'b0011111111001011101010010110001100110100111100010101110110101101;
  assign mem[631] = 64'b1011111111101111001111100110101110111100000110111011110001100101;
  assign mem[632] = 64'b0011111111101101110100011111111011110011100010101001000101011010;
  assign mem[633] = 64'b1011111111010111001101110110001111001001001001100001000010010010;
  assign mem[634] = 64'b0011111111011001110000010111110101000100000011011111100111110010;
  assign mem[635] = 64'b1011111111101101010010110101101100011011000110000111010100100100;
  assign mem[636] = 64'b0011111111100111000110111010110010010110000011100100000110111111;
  assign mem[637] = 64'b1011111111100110001000101110010001001111111011000010001011111111;
  assign mem[638] = 64'b0011111110010101111111010100110100100001111110101011001000100110;
  assign mem[639] = 64'b1011111111101111111111100001110001101000011100001100101101110111;
  assign mem[640] = 64'b0011111111101111111111110000100101000011110001010011101111010001;
  assign mem[641] = 64'b1011111110001111011010100010100101101010101110011001011111001011;
  assign mem[642] = 64'b0011111111100110010001110001010101000011011111110101001101011011;
  assign mem[643] = 64'b1011111111100110111110001100101010011001110010010101101101110101;
  assign mem[644] = 64'b0011111111101101010111110111000101110010100010001000101001111111;
  assign mem[645] = 64'b1011111111011001011001010101010110110111101010111001010010001111;
  assign mem[646] = 64'b0011111111010111100101001111010111100110000100111101111110101110;
  assign mem[647] = 64'b1011111111101101101111111001111001000011100101010111010110011010;
  assign mem[648] = 64'b0011111111101111010010010010001000000110101111001010101110110100;
  assign mem[649] = 64'b1011111111001010111001001111000111010101111100111011100110101011;
  assign mem[650] = 64'b0011111111100001010111100011011011100100110110111110001010111100;
  assign mem[651] = 64'b1011111111101010111000000110100011110011010001011110110011101111;
  assign mem[652] = 64'b0011111111101010010101001100100100010000100100001111010100100011;
  assign mem[653] = 64'b1011111111100010001011110010110101100110001011000001001111100010;
  assign mem[654] = 64'b0011111111000111000010101111110110001101000010001100010011111111;
  assign mem[655] = 64'b1011111111101111011110100010100110011100000110100011001000101010;
  assign mem[656] = 64'b0011111111101111110010110100011100000011100100010100001101010100;
  assign mem[657] = 64'b1011111110111100111111110101001100111011001100000111110111000001;
  assign mem[658] = 64'b0011111111100011111010110011001111101010101111100000011010000000;
  assign mem[659] = 64'b1011111111101001000010110111100101000011010101110101111011111110;
  assign mem[660] = 64'b0011111111101011111111001001110100100101101000011011000101000111;
  assign mem[661] = 64'b1011111111011111000010000001100100000110101111111111011111111110;
  assign mem[662] = 64'b0011111111010001101000101111011111111011111010001111001001000011;
  assign mem[663] = 64'b1011111111101110110000101100111101001011000110101111011010110010;
  assign mem[664] = 64'b0011111111101110011110011101101100101001101001010001011001011010;
  assign mem[665] = 64'b1011111111010011100000111111010111100011010100111011011010101011;
  assign mem[666] = 64'b0011111111011101010011001101000000101011101010000110000010011101;
  assign mem[667] = 64'b1011111111101100011100110001010110001001100111101010101011010111;
  assign mem[668] = 64'b0011111111101000011011000000101000011101100110101010000110010101;
  assign mem[669] = 64'b1011111111100100101011010111100101010001011001110010001011110001;
  assign mem[670] = 64'b0011111110110101001011100111011101001010010011010100110100001010;
  assign mem[671] = 64'b1011111111101111111000111110100100101011111010011101100010000110;
  assign mem[672] = 64'b0011111111101111111011110000000100000010100000100110000110010001;
  assign mem[673] = 64'b1011111110110000011110110110000101001110010001100011000001100100;
  assign mem[674] = 64'b0011111111100101000111111010100000011100110110011001101010100110;
  assign mem[675] = 64'b1011111111101000000010011000101101110101011011100101001011111010;
  assign mem[676] = 64'b0011111111101100101101101110001000001010000000001101101010011001;
  assign mem[677] = 64'b1011111111011100001111110110110101000111001001100011000100101001;
  assign mem[678] = 64'b0011111111010100101000100101001111010001000110111000001011110011;
  assign mem[679] = 64'b1011111111101110010010101000110111111111100000011100111001011110;
  assign mem[680] = 64'b0011111111101110111010110000011101001100010100001010010101000100;
  assign mem[681] = 64'b1011111111010000100000000100111000000101111010110110011000011110;
  assign mem[682] = 64'b0011111111100000000001110100000011001000001010111000001011100001;
  assign mem[683] = 64'b1011111111101011101100100100100110100000101101101100010000001101;
  assign mem[684] = 64'b0011111111101001011010000011111101000010101111010111111111100001;
  assign mem[685] = 64'b1011111111100011011101000101001100011011100000010111111110001101;
  assign mem[686] = 64'b0011111111000000110101100100110110111100101100100110011110000110;
  assign mem[687] = 64'b1011111111101111101110001101000110001101011001101010110110110111;
  assign mem[688] = 64'b0011111111101111100100111111000101001111100001011010110000001000;
  assign mem[689] = 64'b1011111111000100101110001011000101111111011110011111101010001000;
  assign mem[690] = 64'b0011111111100010101010100111011011101000011110101110101101011000;
  assign mem[691] = 64'b1011111111101001111111011111010011110001001100010100100111011110;
  assign mem[692] = 64'b0011111111101011001100010001010110100101111100110111101111110011;
  assign mem[693] = 64'b1011111111100000110111101101000010111000010010111100010010110110;
  assign mem[694] = 64'b0011111111001101001100010111011101001101001011001011110111101110;
  assign mem[695] = 64'b1011111111101111001010000001011111111100010001100000100111001110;
  assign mem[696] = 64'b0011111111101101111101011110001101101010100110111010010110011100;
  assign mem[697] = 64'b1011111111010110011110111001010010011100101011010110001111001011;
  assign mem[698] = 64'b0011111111011010011110010000110011010011110110111111001100011011;
  assign mem[699] = 64'b1011111111101101001000100101010111000110111001011010010011100001;
  assign mem[700] = 64'b0011111111100111011000001100010100101100001100000100011101100100;
  assign mem[701] = 64'b1011111111100101110110011101111011100111001111100011010001011100;
  assign mem[702] = 64'b0011111110100001010001101000010111011011010000101100000101111111;
  assign mem[703] = 64'b1011111111101111111110110101010111100100001001011111110110101110;
  assign mem[704] = 64'b0011111111101111111110010111110001000010000010001100000000010100;
  assign mem[705] = 64'b1011111110100100011010100011100101101111111110000110000101111001;
  assign mem[706] = 64'b0011111111100101101101010000101100100110010011110111010001001000;
  assign mem[707] = 64'b1011111111100111100000101111101100011011100100001011001101011011;
  assign mem[708] = 64'b0011111111101101000011010110011100101111010110011101001010111001;
  assign mem[709] = 64'b1011111111011010110101000111001100010010010111001101110000001001;
  assign mem[710] = 64'b0011111111010110000111010101100101011100100010001100001000000010;
  assign mem[711] = 64'b1011111111101110000001110110011011011001001010000000111101010100;
  assign mem[712] = 64'b0011111111101111000111000111101010111110001010000100011100001000;
  assign mem[713] = 64'b1011111111001101111101010001011000111111000000010000100110011010;
  assign mem[714] = 64'b0011111111100000101101000000010110000111100011111000010111101100;
  assign mem[715] = 64'b1011111111101011010010110111010000001001110111100111100100100101;
  assign mem[716] = 64'b0011111111101001111000001000001011101101101101000010010001110010;
  assign mem[717] = 64'b1011111111100010110100110011001111010011010011101001101110111000;
  assign mem[718] = 64'b0011111111000011111100100010111101010111110110110100100010010011;
  assign mem[719] = 64'b1011111111101111100110111110110101111100111110111101111000101001;
  assign mem[720] = 64'b0011111111101111101100100000110111000110100000011101010101001101;
  assign mem[721] = 64'b1011111111000001100111011000100101000000101111100010010011100111;
  assign mem[722] = 64'b0011111111100011010011000101001001010010110000010100110111100001;
  assign mem[723] = 64'b1011111111101001100001101010111011110001010001010111010110010100;
  assign mem[724] = 64'b0011111111101011100110001111101000011111110110010001010101011110;
  assign mem[725] = 64'b1011111111100000001100101010111001010101111011011011110110010110;
  assign mem[726] = 64'b0011111111010000000111110001100000000110101110011111110111010010;
  assign mem[727] = 64'b1011111111101110111101111101011011100101000111001010001111000000;
  assign mem[728] = 64'b0011111111101110001110100011001111101100011101011100111010000101;
  assign mem[729] = 64'b1011111111010101000000010110001111011100000110010111000001001000;
  assign mem[730] = 64'b0011111111011011111001010001010100010111111111111100000011011001;
  assign mem[731] = 64'b1011111111101100110011001110111000100000110000101101111010100000;
  assign mem[732] = 64'b0011111111100111111010000011111110000111101100000011011010000110;
  assign mem[733] = 64'b1011111111100101010001010100111111110101000101011001110111111100;
  assign mem[734] = 64'b0011111110101101110101000000011011111001100000001000111011001001;
  assign mem[735] = 64'b1011111111101111111100100001011000010100111000010011000111101101;
  assign mem[736] = 64'b0011111111101111110111111001100100100010111101110011001100000111;
  assign mem[737] = 64'b1011111110110110101111110001101100111110011110011011000100101001;
  assign mem[738] = 64'b0011111111100100100001110000001100110000011000001001000111111111;
  assign mem[739] = 64'b1011111111101000100011000110011011100111010010000001101110100001;
  assign mem[740] = 64'b0011111111101100010110111110111101011001111111101111100001011010;
  assign mem[741] = 64'b1011111111011101101001100000110001011100111110100001000011011001;
  assign mem[742] = 64'b0011111111010011001001000001111110110110001110001011101010101111;
  assign mem[743] = 64'b1011111111101110100010010000100101011011101011010110000000100101;
  assign mem[744] = 64'b0011111111101110101101001100111101010001010110111000100000010001;
  assign mem[745] = 64'b1011111111010010000000111000010110000011110101110010011110111110;
  assign mem[746] = 64'b0011111111011110101100000000011010010101111100100101011000100000;
  assign mem[747] = 64'b1011111111101100000101001101100111011100010001100101111001010111;
  assign mem[748] = 64'b0011111111101000111011000001000010011011010010000110110001001001;
  assign mem[749] = 64'b1011111111100100000100100111001001100110001111010001000010001100;
  assign mem[750] = 64'b0011111110111011011011111010011011101100001110001111011001001100;
  assign mem[751] = 64'b1011111111101111110100001101000101011000110110000110000010000111;
  assign mem[752] = 64'b0011111111101111011100001111011001000011010010110111111010110111;
  assign mem[753] = 64'b1011111111000111110100001010011110111011110100101100101100011100;
  assign mem[754] = 64'b0011111111100010000001011011101010100001011101010110000011010110;
  assign mem[755] = 64'b1011111111101010011100010011100011011110100111010110000011110101;
  assign mem[756] = 64'b0011111111101010110001001111111110111101001111101111101011001000;
  assign mem[757] = 64'b1011111111100001100010000101100100011111001110100100011011100101;
  assign mem[758] = 64'b0011111111001010001000000011111000011011000110000011000111011010;
  assign mem[759] = 64'b1011111111101111010100111000101100011111101011110010110100000111;
  assign mem[760] = 64'b0011111111101101101011001111010000101100111001101000101010111001;
  assign mem[761] = 64'b1011111111010111111100100100110111010011011100110100000111100100;
  assign mem[762] = 64'b0011111111011001000010001110111110000001111011110111101111010001;
  assign mem[763] = 64'b1011111111101101011100110011111101010000100011000000110111111111;
  assign mem[764] = 64'b0011111111100110110101011010111111101111010010101010111111001101;
  assign mem[765] = 64'b1011111111100110011010110000111100111111010100101011001110000110;
  assign mem[766] = 64'b0011111110000010110110010110101100001110010100001001011100000011;
  assign mem[767] = 64'b1011111111101111111111111010011100101100100101111000110001001111;
  assign mem[768] = 64'b0011111111101111111111111010011100101100100101111000110001001111;
  assign mem[769] = 64'b1011111110000010110110010110101100001110010100001001011100000011;
  assign mem[770] = 64'b0011111111100110011010110000111100111111010100101011001110000110;
  assign mem[771] = 64'b1011111111100110110101011010111111101111010010101010111111001101;
  assign mem[772] = 64'b0011111111101101011100110011111101010000100011000000110111111111;
  assign mem[773] = 64'b1011111111011001000010001110111110000001111011110111101111010001;
  assign mem[774] = 64'b0011111111010111111100100100110111010011011100110100000111100100;
  assign mem[775] = 64'b1011111111101101101011001111010000101100111001101000101010111001;
  assign mem[776] = 64'b0011111111101111010100111000101100011111101011110010110100000111;
  assign mem[777] = 64'b1011111111001010001000000011111000011011000110000011000111011010;
  assign mem[778] = 64'b0011111111100001100010000101100100011111001110100100011011100101;
  assign mem[779] = 64'b1011111111101010110001001111111110111101001111101111101011001000;
  assign mem[780] = 64'b0011111111101010011100010011100011011110100111010110000011110101;
  assign mem[781] = 64'b1011111111100010000001011011101010100001011101010110000011010110;
  assign mem[782] = 64'b0011111111000111110100001010011110111011110100101100101100011100;
  assign mem[783] = 64'b1011111111101111011100001111011001000011010010110111111010110111;
  assign mem[784] = 64'b0011111111101111110100001101000101011000110110000110000010000111;
  assign mem[785] = 64'b1011111110111011011011111010011011101100001110001111011001001100;
  assign mem[786] = 64'b0011111111100100000100100111001001100110001111010001000010001100;
  assign mem[787] = 64'b1011111111101000111011000001000010011011010010000110110001001001;
  assign mem[788] = 64'b0011111111101100000101001101100111011100010001100101111001010111;
  assign mem[789] = 64'b1011111111011110101100000000011010010101111100100101011000100000;
  assign mem[790] = 64'b0011111111010010000000111000010110000011110101110010011110111110;
  assign mem[791] = 64'b1011111111101110101101001100111101010001010110111000100000010001;
  assign mem[792] = 64'b0011111111101110100010010000100101011011101011010110000000100101;
  assign mem[793] = 64'b1011111111010011001001000001111110110110001110001011101010101111;
  assign mem[794] = 64'b0011111111011101101001100000110001011100111110100001000011011001;
  assign mem[795] = 64'b1011111111101100010110111110111101011001111111101111100001011010;
  assign mem[796] = 64'b0011111111101000100011000110011011100111010010000001101110100001;
  assign mem[797] = 64'b1011111111100100100001110000001100110000011000001001000111111111;
  assign mem[798] = 64'b0011111110110110101111110001101100111110011110011011000100101001;
  assign mem[799] = 64'b1011111111101111110111111001100100100010111101110011001100000111;
  assign mem[800] = 64'b0011111111101111111100100001011000010100111000010011000111101101;
  assign mem[801] = 64'b1011111110101101110101000000011011111001100000001000111011001001;
  assign mem[802] = 64'b0011111111100101010001010100111111110101000101011001110111111100;
  assign mem[803] = 64'b1011111111100111111010000011111110000111101100000011011010000110;
  assign mem[804] = 64'b0011111111101100110011001110111000100000110000101101111010100000;
  assign mem[805] = 64'b1011111111011011111001010001010100010111111111111100000011011001;
  assign mem[806] = 64'b0011111111010101000000010110001111011100000110010111000001001000;
  assign mem[807] = 64'b1011111111101110001110100011001111101100011101011100111010000101;
  assign mem[808] = 64'b0011111111101110111101111101011011100101000111001010001111000000;
  assign mem[809] = 64'b1011111111010000000111110001100000000110101110011111110111010010;
  assign mem[810] = 64'b0011111111100000001100101010111001010101111011011011110110010110;
  assign mem[811] = 64'b1011111111101011100110001111101000011111110110010001010101011110;
  assign mem[812] = 64'b0011111111101001100001101010111011110001010001010111010110010100;
  assign mem[813] = 64'b1011111111100011010011000101001001010010110000010100110111100001;
  assign mem[814] = 64'b0011111111000001100111011000100101000000101111100010010011100111;
  assign mem[815] = 64'b1011111111101111101100100000110111000110100000011101010101001101;
  assign mem[816] = 64'b0011111111101111100110111110110101111100111110111101111000101001;
  assign mem[817] = 64'b1011111111000011111100100010111101010111110110110100100010010011;
  assign mem[818] = 64'b0011111111100010110100110011001111010011010011101001101110111000;
  assign mem[819] = 64'b1011111111101001111000001000001011101101101101000010010001110010;
  assign mem[820] = 64'b0011111111101011010010110111010000001001110111100111100100100101;
  assign mem[821] = 64'b1011111111100000101101000000010110000111100011111000010111101100;
  assign mem[822] = 64'b0011111111001101111101010001011000111111000000010000100110011010;
  assign mem[823] = 64'b1011111111101111000111000111101010111110001010000100011100001000;
  assign mem[824] = 64'b0011111111101110000001110110011011011001001010000000111101010100;
  assign mem[825] = 64'b1011111111010110000111010101100101011100100010001100001000000010;
  assign mem[826] = 64'b0011111111011010110101000111001100010010010111001101110000001001;
  assign mem[827] = 64'b1011111111101101000011010110011100101111010110011101001010111001;
  assign mem[828] = 64'b0011111111100111100000101111101100011011100100001011001101011011;
  assign mem[829] = 64'b1011111111100101101101010000101100100110010011110111010001001000;
  assign mem[830] = 64'b0011111110100100011010100011100101101111111110000110000101111001;
  assign mem[831] = 64'b1011111111101111111110010111110001000010000010001100000000010100;
  assign mem[832] = 64'b0011111111101111111110110101010111100100001001011111110110101110;
  assign mem[833] = 64'b1011111110100001010001101000010111011011010000101100000101111111;
  assign mem[834] = 64'b0011111111100101110110011101111011100111001111100011010001011100;
  assign mem[835] = 64'b1011111111100111011000001100010100101100001100000100011101100100;
  assign mem[836] = 64'b0011111111101101001000100101010111000110111001011010010011100001;
  assign mem[837] = 64'b1011111111011010011110010000110011010011110110111111001100011011;
  assign mem[838] = 64'b0011111111010110011110111001010010011100101011010110001111001011;
  assign mem[839] = 64'b1011111111101101111101011110001101101010100110111010010110011100;
  assign mem[840] = 64'b0011111111101111001010000001011111111100010001100000100111001110;
  assign mem[841] = 64'b1011111111001101001100010111011101001101001011001011110111101110;
  assign mem[842] = 64'b0011111111100000110111101101000010111000010010111100010010110110;
  assign mem[843] = 64'b1011111111101011001100010001010110100101111100110111101111110011;
  assign mem[844] = 64'b0011111111101001111111011111010011110001001100010100100111011110;
  assign mem[845] = 64'b1011111111100010101010100111011011101000011110101110101101011000;
  assign mem[846] = 64'b0011111111000100101110001011000101111111011110011111101010001000;
  assign mem[847] = 64'b1011111111101111100100111111000101001111100001011010110000001000;
  assign mem[848] = 64'b0011111111101111101110001101000110001101011001101010110110110111;
  assign mem[849] = 64'b1011111111000000110101100100110110111100101100100110011110000110;
  assign mem[850] = 64'b0011111111100011011101000101001100011011100000010111111110001101;
  assign mem[851] = 64'b1011111111101001011010000011111101000010101111010111111111100001;
  assign mem[852] = 64'b0011111111101011101100100100100110100000101101101100010000001101;
  assign mem[853] = 64'b1011111111100000000001110100000011001000001010111000001011100001;
  assign mem[854] = 64'b0011111111010000100000000100111000000101111010110110011000011110;
  assign mem[855] = 64'b1011111111101110111010110000011101001100010100001010010101000100;
  assign mem[856] = 64'b0011111111101110010010101000110111111111100000011100111001011110;
  assign mem[857] = 64'b1011111111010100101000100101001111010001000110111000001011110011;
  assign mem[858] = 64'b0011111111011100001111110110110101000111001001100011000100101001;
  assign mem[859] = 64'b1011111111101100101101101110001000001010000000001101101010011001;
  assign mem[860] = 64'b0011111111101000000010011000101101110101011011100101001011111010;
  assign mem[861] = 64'b1011111111100101000111111010100000011100110110011001101010100110;
  assign mem[862] = 64'b0011111110110000011110110110000101001110010001100011000001100100;
  assign mem[863] = 64'b1011111111101111111011110000000100000010100000100110000110010001;
  assign mem[864] = 64'b0011111111101111111000111110100100101011111010011101100010000110;
  assign mem[865] = 64'b1011111110110101001011100111011101001010010011010100110100001010;
  assign mem[866] = 64'b0011111111100100101011010111100101010001011001110010001011110001;
  assign mem[867] = 64'b1011111111101000011011000000101000011101100110101010000110010101;
  assign mem[868] = 64'b0011111111101100011100110001010110001001100111101010101011010111;
  assign mem[869] = 64'b1011111111011101010011001101000000101011101010000110000010011101;
  assign mem[870] = 64'b0011111111010011100000111111010111100011010100111011011010101011;
  assign mem[871] = 64'b1011111111101110011110011101101100101001101001010001011001011010;
  assign mem[872] = 64'b0011111111101110110000101100111101001011000110101111011010110010;
  assign mem[873] = 64'b1011111111010001101000101111011111111011111010001111001001000011;
  assign mem[874] = 64'b0011111111011111000010000001100100000110101111111111011111111110;
  assign mem[875] = 64'b1011111111101011111111001001110100100101101000011011000101000111;
  assign mem[876] = 64'b0011111111101001000010110111100101000011010101110101111011111110;
  assign mem[877] = 64'b1011111111100011111010110011001111101010101111100000011010000000;
  assign mem[878] = 64'b0011111110111100111111110101001100111011001100000111110111000001;
  assign mem[879] = 64'b1011111111101111110010110100011100000011100100010100001101010100;
  assign mem[880] = 64'b0011111111101111011110100010100110011100000110100011001000101010;
  assign mem[881] = 64'b1011111111000111000010101111110110001101000010001100010011111111;
  assign mem[882] = 64'b0011111111100010001011110010110101100110001011000001001111100010;
  assign mem[883] = 64'b1011111111101010010101001100100100010000100100001111010100100011;
  assign mem[884] = 64'b0011111111101010111000000110100011110011010001011110110011101111;
  assign mem[885] = 64'b1011111111100001010111100011011011100100110110111110001010111100;
  assign mem[886] = 64'b0011111111001010111001001111000111010101111100111011100110101011;
  assign mem[887] = 64'b1011111111101111010010010010001000000110101111001010101110110100;
  assign mem[888] = 64'b0011111111101101101111111001111001000011100101010111010110011010;
  assign mem[889] = 64'b1011111111010111100101001111010111100110000100111101111110101110;
  assign mem[890] = 64'b0011111111011001011001010101010110110111101010111001010010001111;
  assign mem[891] = 64'b1011111111101101010111110111000101110010100010001000101001111111;
  assign mem[892] = 64'b0011111111100110111110001100101010011001110010010101101101110101;
  assign mem[893] = 64'b1011111111100110010001110001010101000011011111110101001101011011;
  assign mem[894] = 64'b0011111110001111011010100010100101101010101110011001011111001011;
  assign mem[895] = 64'b1011111111101111111111110000100101000011110001010011101111010001;
  assign mem[896] = 64'b0011111111101111111111100001110001101000011100001100101101110111;
  assign mem[897] = 64'b1011111110010101111111010100110100100001111110101011001000100110;
  assign mem[898] = 64'b0011111111100110001000101110010001001111111011000010001011111111;
  assign mem[899] = 64'b1011111111100111000110111010110010010110000011100100000110111111;
  assign mem[900] = 64'b0011111111101101010010110101101100011011000110000111010100100100;
  assign mem[901] = 64'b1011111111011001110000010111110101000100000011011111100111110010;
  assign mem[902] = 64'b0011111111010111001101110110001111001001001001100001000010010010;
  assign mem[903] = 64'b1011111111101101110100011111111011110011100010101001000101011010;
  assign mem[904] = 64'b0011111111101111001111100110101110111100000110111011110001100101;
  assign mem[905] = 64'b1011111111001011101010010110001100110100111100010101110110101101;
  assign mem[906] = 64'b0011111111100001001100111110100111001111111011100010010101001111;
  assign mem[907] = 64'b1011111111101010111110111000111111011000100111110101011110110110;
  assign mem[908] = 64'b0011111111101010001110000001100001001010010110010011101111000110;
  assign mem[909] = 64'b1011111111100010010110000111001101001100101110110111000100010000;
  assign mem[910] = 64'b0011111111000110010001010001101010000011000111011000001100001101;
  assign mem[911] = 64'b1011111111101111100000110000111101001010010000001100011000001100;
  assign mem[912] = 64'b0011111111101111110001010110111000111011011111011001101011110110;
  assign mem[913] = 64'b1011111110111110100011101011011111111101111001001010101000111111;
  assign mem[914] = 64'b0011111111100011110000111100010001001001100000011100010100011000;
  assign mem[915] = 64'b1011111111101001001010101010010000011111110001011010100000010101;
  assign mem[916] = 64'b0011111111101011111001000001101101100001000100010101010011000001;
  assign mem[917] = 64'b1011111111011111010111111101111011100110010101101100110110100011;
  assign mem[918] = 64'b0011111111010001010000100011111011101111110001101001001101111000;
  assign mem[919] = 64'b1011111111101110110100001000001101011110100110011001000000001001;
  assign mem[920] = 64'b0011111111101110011010100110000111000101010111010101001110100111;
  assign mem[921] = 64'b1011111111010011111000111001101111101001011011101100001001110001;
  assign mem[922] = 64'b0011111111011100111100110100101110101110111000011100110100100001;
  assign mem[923] = 64'b1011111111101100100010011111010110000111000000101001110000010011;
  assign mem[924] = 64'b0011111111101000010010110111000100010001101011111000001111111010;
  assign mem[925] = 64'b1011111111100100110100111011110001101101010110001001111101111111;
  assign mem[926] = 64'b0011111110110011100111011001111100010010110001011010001010011001;
  assign mem[927] = 64'b1011111111101111111001111110101010000101010010000010110101100000;
  assign mem[928] = 64'b0011111111101111111010111001110100100101001100000100000100001111;
  assign mem[929] = 64'b1011111110110010000011001001011001110100111011010100010001001101;
  assign mem[930] = 64'b0011111111100100111110011100110000100101110011001010010010000110;
  assign mem[931] = 64'b1011111111101000001010101001110000010011111101010100010111111111;
  assign mem[932] = 64'b0011111111101100101000001000111100011001101110011100010001001001;
  assign mem[933] = 64'b1011111111011100100110010111111111000011100001100101001110001001;
  assign mem[934] = 64'b0011111111010100010000110001000011011100100010010011011011110000;
  assign mem[935] = 64'b1011111111101110010110101001110101010101000001000110011111010011;
  assign mem[936] = 64'b0011111111101110110111011110101101101010000001111000011001010001;
  assign mem[937] = 64'b1011111111010000111000010101101101001110000101110100100111001110;
  assign mem[938] = 64'b0011111111011111101101110101011101011100001001001101001011011110;
  assign mem[939] = 64'b1011111111101011110010110101010011001011000011010010001100100111;
  assign mem[940] = 64'b0011111111101001010010011001000011100011101011000100101001101100;
  assign mem[941] = 64'b1011111111100011100111000010001111100011110101100011000000101001;
  assign mem[942] = 64'b0011111111000000000011101110100010101101011011111011100001011011;
  assign mem[943] = 64'b1011111111101111101111110100011100001111000010101000110110001000;
  assign mem[944] = 64'b0011111111101111100010111010011100110111110010110100101101111000;
  assign mem[945] = 64'b1011111111000101011111110000000010000110010101001100101111011110;
  assign mem[946] = 64'b0011111111100010100000011000101111101111010011010011110010111010;
  assign mem[947] = 64'b1011111111101010000110110010011011010010110000001010011101011110;
  assign mem[948] = 64'b0011111111101011000101100111010000101010010011001010001011110101;
  assign mem[949] = 64'b1011111111100001000010010111001001001000110100001010100101010111;
  assign mem[950] = 64'b0011111111001100011011011001000001010011010111010111010011011101;
  assign mem[951] = 64'b1011111111101111001100110110100001011010001110101010111011110000;
  assign mem[952] = 64'b0011111111101101111001000001011000001111011011011000110110000001;
  assign mem[953] = 64'b1011111111010110110110011001100001100011100010100000110010110110;
  assign mem[954] = 64'b0011111111011010000111010110010101000011101101010000101011000000;
  assign mem[955] = 64'b1011111111101101001101101111110001111011110010111111101111011100;
  assign mem[956] = 64'b0011111111100111001111100101010110001110000001111001100101000010;
  assign mem[957] = 64'b1011111111100101111111100111110010111101111001010110101000010000;
  assign mem[958] = 64'b0011111110011100010001010100111101001100111001010011101100011101;
  assign mem[959] = 64'b1011111111101111111111001110000010011100111000101010011001111001;
  assign mem[960] = 64'b0011111111101111111101110101001110111011000110111001000101100100;
  assign mem[961] = 64'b1011111110100111100011011011101010100101100001110100011010000110;
  assign mem[962] = 64'b0011111111100101100100000000000111010101111101110010001111011111;
  assign mem[963] = 64'b1011111111100111101001001111011100000111101111111001011111010010;
  assign mem[964] = 64'b0011111111101100111110000011000011101000110011100100011001111011;
  assign mem[965] = 64'b1011111111011011001011111001011100011101101100110001100101110010;
  assign mem[966] = 64'b0011111111010101101111101110011110001011100111011011001110110110;
  assign mem[967] = 64'b1011111111101110000110001010000000101111110111000110011011011001;
  assign mem[968] = 64'b0011111111101111000100001001000010111100100010011000111101011111;
  assign mem[969] = 64'b1011111111001110101110000110101101000110001011011110001101001000;
  assign mem[970] = 64'b0011111111100000100010010001000100100000001100101011000010001100;
  assign mem[971] = 64'b1011111111101011011001011000111100010100111111011011110001000111;
  assign mem[972] = 64'b0011111111101001110000101101000100010000111100000111010111000010;
  assign mem[973] = 64'b1011111111100010111110111100001001001011010001000001000000010101;
  assign mem[974] = 64'b0011111111000011001010110111101111111001010001010001011010100111;
  assign mem[975] = 64'b1011111111101111101000111001101110101100011110100001011110010001;
  assign mem[976] = 64'b0011111111101111101010101111101111001011000011001111110111011100;
  assign mem[977] = 64'b1011111111000010011001001001100101001101111111010011010000001001;
  assign mem[978] = 64'b0011111111100011001001000010000111101100010010011010011000011111;
  assign mem[979] = 64'b1011111111101001101001001101111110100100001010110000011010110010;
  assign mem[980] = 64'b0011111111101011011111110110011010000110111001111001001011101001;
  assign mem[981] = 64'b1011111111100000010111011111001111101100001100011011100010110111;
  assign mem[982] = 64'b0011111111001111011110110111010010000000101111010011100000000010;
  assign mem[983] = 64'b1011111111101111000001000101101000010100110011110111001110001100;
  assign mem[984] = 64'b0011111111101110001010011000111101000100001110010001100101111010;
  assign mem[985] = 64'b1011111111010101011000000100000000010010111101000110011110110100;
  assign mem[986] = 64'b0011111111011011100010100111100000010100111111010101011010010011;
  assign mem[987] = 64'b1011111111101100111000101011001100100111100110011010000001100000;
  assign mem[988] = 64'b0011111111100111110001101011100010011100111000101101001100110011;
  assign mem[989] = 64'b1011111111100101011010101100001101010001100101110110010010011111;
  assign mem[990] = 64'b0011111110101010101100010000000110111101010111111000001100010111;
  assign mem[991] = 64'b1011111111101111111101001101110001010100101100011011111011010011;
  assign mem[992] = 64'b0011111111101111110110101111101001110101000101000101001110001100;
  assign mem[993] = 64'b1011111110111000010011111000011100010010110000010011000010100001;
  assign mem[994] = 64'b0011111111100100011000000101101001101001001010110011001010100010;
  assign mem[995] = 64'b1011111111101000101011001000011100011110110111100001110110001000;
  assign mem[996] = 64'b0011111111101100010001001000001100110001010000011100000000000100;
  assign mem[997] = 64'b1011111111011101111111101111111101100110101010010100000111011110;
  assign mem[998] = 64'b0011111111010010110001000001101001001110100101010100010100100000;
  assign mem[999] = 64'b1011111111101110100101111110110000110110000000010110101100110000;
  assign mem[1000] = 64'b0011111111101110101001101000001110010011111001100101100000000000;
  assign mem[1001] = 64'b1011111111010010011000111110011010011001010101010101010010111010;
  assign mem[1002] = 64'b0011111111011110010101111010100001101101001111001101100000100101;
  assign mem[1003] = 64'b1011111111101100001011001101000101001001001100011110001111110001;
  assign mem[1004] = 64'b0011111111101000110011000110101001110101000110000100011001010101;
  assign mem[1005] = 64'b1011111111100100001110010111111101011011001010100100001110000000;
  assign mem[1006] = 64'b0011111110111001110111111011011011101011001001001010100001011100;
  assign mem[1007] = 64'b1011111111101111110101100000110100101101101001110101110010011110;
  assign mem[1008] = 64'b0011111111101111011001110111010101010110100010000011110011101110;
  assign mem[1009] = 64'b1011111111001000100101100001011100100111110001000001100000000100;
  assign mem[1010] = 64'b0011111111100001110111000001101101100100110111000100100001110010;
  assign mem[1011] = 64'b1011111111101010100011010110011101101110010101000101101011010010;
  assign mem[1012] = 64'b0011111111101010101010010101010001111010001011001011100110001110;
  assign mem[1013] = 64'b1011111111100001101100100101000000010111000100110111001110111111;
  assign mem[1014] = 64'b0011111111001001010110110100100111101001101101100010101011111010;
  assign mem[1015] = 64'b1011111111101111010111011010011011101101010000110110100001011101;
  assign mem[1016] = 64'b0011111111101101100110100000000011011101100010110011110101000110;
  assign mem[1017] = 64'b1011111111011000010011110110101010101010111100111001000000111111;
  assign mem[1018] = 64'b0011111111011000101011000100101110000110110101011110110101000100;
  assign mem[1019] = 64'b1011111111101101100001101100010010000100010001011010010001001111;
  assign mem[1020] = 64'b0011111111100110101100100101110011101101001011111110001010011100;
  assign mem[1021] = 64'b1011111111100110100011101101000111101010101000011001110001110001;
  assign mem[1022] = 64'b0011111101101001001000011111100010111110110011001010010010111010;
  assign mem[1023] = 64'b1011111111101111111111111111011000100001011000100001110100000010;

  always@(*)
  begin
    data_out_t <= mem[addr_f];
  end

  // Build output registers
  wire [63:0] data_out_reg [n_outreg:0];
  generate if (n_outreg > 0)
  begin
    for( i=n_outreg-1; i >= 1; i=i-1)
    begin: data_out_reg_stage
      mgc_generic_reg #(
        .width(64), 
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_data_out_reg (
        .d(data_out_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(data_out_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(64), 
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_data_out_reg_init (
      .d(data_out_t),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(data_out_reg[0])
    );
    assign data_out = data_out_reg[n_outreg-1];
  end
  else
  begin
    assign data_out = data_out_t;
  end
  endgenerate

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Sun Oct  6 01:48:33 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_7_16_10_1024_1024_16_5_gen
// ------------------------------------------------------------------


module stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_7_16_10_1024_1024_16_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [15:0] q;
  output we;
  output [15:0] d;
  output [9:0] adr;
  input [9:0] adr_d;
  input [15:0] d_d;
  input en_d;
  input we_d;
  output [15:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_6_64_10_1024_1024_64_5_gen
// ------------------------------------------------------------------


module stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_6_64_10_1024_1024_64_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [9:0] adr;
  input [9:0] adr_d;
  input [63:0] d_d;
  input en_d;
  input we_d;
  output [63:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_5_16_10_1024_1024_16_5_gen
// ------------------------------------------------------------------


module stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_5_16_10_1024_1024_16_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [15:0] q;
  output we;
  output [15:0] d;
  output [9:0] adr;
  input [9:0] adr_d;
  input [15:0] d_d;
  input en_d;
  input we_d;
  output [15:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_4_64_10_1024_1024_64_5_gen
// ------------------------------------------------------------------


module stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_4_64_10_1024_1024_64_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [9:0] adr;
  input [9:0] adr_d;
  input [63:0] d_d;
  input en_d;
  input we_d;
  output [63:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module stage_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output, for_C_0_tr0, BUTTERFLY_C_15_tr0, BUTTERFLY_C_15_tr1,
      BUTTERFLY_1_C_15_tr0, BUTTERFLY_1_C_15_tr1, for_1_C_2_tr0
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [38:0] fsm_output;
  reg [38:0] fsm_output;
  input for_C_0_tr0;
  input BUTTERFLY_C_15_tr0;
  input BUTTERFLY_C_15_tr1;
  input BUTTERFLY_1_C_15_tr0;
  input BUTTERFLY_1_C_15_tr1;
  input for_1_C_2_tr0;


  // FSM State Type Declaration for stage_run_run_fsm_1
  parameter
    run_rlp_C_0 = 6'd0,
    main_C_0 = 6'd1,
    for_C_0 = 6'd2,
    BUTTERFLY_C_0 = 6'd3,
    BUTTERFLY_C_1 = 6'd4,
    BUTTERFLY_C_2 = 6'd5,
    BUTTERFLY_C_3 = 6'd6,
    BUTTERFLY_C_4 = 6'd7,
    BUTTERFLY_C_5 = 6'd8,
    BUTTERFLY_C_6 = 6'd9,
    BUTTERFLY_C_7 = 6'd10,
    BUTTERFLY_C_8 = 6'd11,
    BUTTERFLY_C_9 = 6'd12,
    BUTTERFLY_C_10 = 6'd13,
    BUTTERFLY_C_11 = 6'd14,
    BUTTERFLY_C_12 = 6'd15,
    BUTTERFLY_C_13 = 6'd16,
    BUTTERFLY_C_14 = 6'd17,
    BUTTERFLY_C_15 = 6'd18,
    BUTTERFLY_1_C_0 = 6'd19,
    BUTTERFLY_1_C_1 = 6'd20,
    BUTTERFLY_1_C_2 = 6'd21,
    BUTTERFLY_1_C_3 = 6'd22,
    BUTTERFLY_1_C_4 = 6'd23,
    BUTTERFLY_1_C_5 = 6'd24,
    BUTTERFLY_1_C_6 = 6'd25,
    BUTTERFLY_1_C_7 = 6'd26,
    BUTTERFLY_1_C_8 = 6'd27,
    BUTTERFLY_1_C_9 = 6'd28,
    BUTTERFLY_1_C_10 = 6'd29,
    BUTTERFLY_1_C_11 = 6'd30,
    BUTTERFLY_1_C_12 = 6'd31,
    BUTTERFLY_1_C_13 = 6'd32,
    BUTTERFLY_1_C_14 = 6'd33,
    BUTTERFLY_1_C_15 = 6'd34,
    for_1_C_0 = 6'd35,
    for_1_C_1 = 6'd36,
    for_1_C_2 = 6'd37,
    main_C_1 = 6'd38;

  reg [5:0] state_var;
  reg [5:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : stage_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 39'b000000000000000000000000000000000000010;
        state_var_NS = for_C_0;
      end
      for_C_0 : begin
        fsm_output = 39'b000000000000000000000000000000000000100;
        if ( for_C_0_tr0 ) begin
          state_var_NS = BUTTERFLY_C_0;
        end
        else begin
          state_var_NS = BUTTERFLY_1_C_0;
        end
      end
      BUTTERFLY_C_0 : begin
        fsm_output = 39'b000000000000000000000000000000000001000;
        state_var_NS = BUTTERFLY_C_1;
      end
      BUTTERFLY_C_1 : begin
        fsm_output = 39'b000000000000000000000000000000000010000;
        state_var_NS = BUTTERFLY_C_2;
      end
      BUTTERFLY_C_2 : begin
        fsm_output = 39'b000000000000000000000000000000000100000;
        state_var_NS = BUTTERFLY_C_3;
      end
      BUTTERFLY_C_3 : begin
        fsm_output = 39'b000000000000000000000000000000001000000;
        state_var_NS = BUTTERFLY_C_4;
      end
      BUTTERFLY_C_4 : begin
        fsm_output = 39'b000000000000000000000000000000010000000;
        state_var_NS = BUTTERFLY_C_5;
      end
      BUTTERFLY_C_5 : begin
        fsm_output = 39'b000000000000000000000000000000100000000;
        state_var_NS = BUTTERFLY_C_6;
      end
      BUTTERFLY_C_6 : begin
        fsm_output = 39'b000000000000000000000000000001000000000;
        state_var_NS = BUTTERFLY_C_7;
      end
      BUTTERFLY_C_7 : begin
        fsm_output = 39'b000000000000000000000000000010000000000;
        state_var_NS = BUTTERFLY_C_8;
      end
      BUTTERFLY_C_8 : begin
        fsm_output = 39'b000000000000000000000000000100000000000;
        state_var_NS = BUTTERFLY_C_9;
      end
      BUTTERFLY_C_9 : begin
        fsm_output = 39'b000000000000000000000000001000000000000;
        state_var_NS = BUTTERFLY_C_10;
      end
      BUTTERFLY_C_10 : begin
        fsm_output = 39'b000000000000000000000000010000000000000;
        state_var_NS = BUTTERFLY_C_11;
      end
      BUTTERFLY_C_11 : begin
        fsm_output = 39'b000000000000000000000000100000000000000;
        state_var_NS = BUTTERFLY_C_12;
      end
      BUTTERFLY_C_12 : begin
        fsm_output = 39'b000000000000000000000001000000000000000;
        state_var_NS = BUTTERFLY_C_13;
      end
      BUTTERFLY_C_13 : begin
        fsm_output = 39'b000000000000000000000010000000000000000;
        state_var_NS = BUTTERFLY_C_14;
      end
      BUTTERFLY_C_14 : begin
        fsm_output = 39'b000000000000000000000100000000000000000;
        state_var_NS = BUTTERFLY_C_15;
      end
      BUTTERFLY_C_15 : begin
        fsm_output = 39'b000000000000000000001000000000000000000;
        if ( BUTTERFLY_C_15_tr0 ) begin
          state_var_NS = for_1_C_0;
        end
        else if ( BUTTERFLY_C_15_tr1 ) begin
          state_var_NS = BUTTERFLY_C_0;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      BUTTERFLY_1_C_0 : begin
        fsm_output = 39'b000000000000000000010000000000000000000;
        state_var_NS = BUTTERFLY_1_C_1;
      end
      BUTTERFLY_1_C_1 : begin
        fsm_output = 39'b000000000000000000100000000000000000000;
        state_var_NS = BUTTERFLY_1_C_2;
      end
      BUTTERFLY_1_C_2 : begin
        fsm_output = 39'b000000000000000001000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_3;
      end
      BUTTERFLY_1_C_3 : begin
        fsm_output = 39'b000000000000000010000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_4;
      end
      BUTTERFLY_1_C_4 : begin
        fsm_output = 39'b000000000000000100000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_5;
      end
      BUTTERFLY_1_C_5 : begin
        fsm_output = 39'b000000000000001000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_6;
      end
      BUTTERFLY_1_C_6 : begin
        fsm_output = 39'b000000000000010000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_7;
      end
      BUTTERFLY_1_C_7 : begin
        fsm_output = 39'b000000000000100000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_8;
      end
      BUTTERFLY_1_C_8 : begin
        fsm_output = 39'b000000000001000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_9;
      end
      BUTTERFLY_1_C_9 : begin
        fsm_output = 39'b000000000010000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_10;
      end
      BUTTERFLY_1_C_10 : begin
        fsm_output = 39'b000000000100000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_11;
      end
      BUTTERFLY_1_C_11 : begin
        fsm_output = 39'b000000001000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_12;
      end
      BUTTERFLY_1_C_12 : begin
        fsm_output = 39'b000000010000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_13;
      end
      BUTTERFLY_1_C_13 : begin
        fsm_output = 39'b000000100000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_14;
      end
      BUTTERFLY_1_C_14 : begin
        fsm_output = 39'b000001000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_15;
      end
      BUTTERFLY_1_C_15 : begin
        fsm_output = 39'b000010000000000000000000000000000000000;
        if ( BUTTERFLY_1_C_15_tr0 ) begin
          state_var_NS = for_1_C_0;
        end
        else if ( BUTTERFLY_1_C_15_tr1 ) begin
          state_var_NS = BUTTERFLY_1_C_0;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      for_1_C_0 : begin
        fsm_output = 39'b000100000000000000000000000000000000000;
        state_var_NS = for_1_C_1;
      end
      for_1_C_1 : begin
        fsm_output = 39'b001000000000000000000000000000000000000;
        state_var_NS = for_1_C_2;
      end
      for_1_C_2 : begin
        fsm_output = 39'b010000000000000000000000000000000000000;
        if ( for_1_C_2_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_1_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 39'b100000000000000000000000000000000000000;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 39'b000000000000000000000000000000000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_staller
// ------------------------------------------------------------------


module stage_run_staller (
  clk, rst, arst_n, run_wen, run_wten, ap_start_rsci_wen_comp, ap_done_rsci_wen_comp,
      out1_rsci_wen_comp
);
  input clk;
  input rst;
  input arst_n;
  output run_wen;
  output run_wten;
  reg run_wten;
  input ap_start_rsci_wen_comp;
  input ap_done_rsci_wen_comp;
  input out1_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = ap_start_rsci_wen_comp & ap_done_rsci_wen_comp & out1_rsci_wen_comp;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten <= 1'b0;
    end
    else if ( rst ) begin
      run_wten <= 1'b0;
    end
    else begin
      run_wten <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_out_u_triosy_obj_out_u_triosy_wait_ctrl
// ------------------------------------------------------------------


module stage_run_out_u_triosy_obj_out_u_triosy_wait_ctrl (
  run_wten, out_u_triosy_obj_iswt0, out_u_triosy_obj_biwt
);
  input run_wten;
  input out_u_triosy_obj_iswt0;
  output out_u_triosy_obj_biwt;



  // Interconnect Declarations for Component Instantiations 
  assign out_u_triosy_obj_biwt = (~ run_wten) & out_u_triosy_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_out_f_d_triosy_obj_out_f_d_triosy_wait_ctrl
// ------------------------------------------------------------------


module stage_run_out_f_d_triosy_obj_out_f_d_triosy_wait_ctrl (
  run_wten, out_f_d_triosy_obj_iswt0, out_f_d_triosy_obj_biwt
);
  input run_wten;
  input out_f_d_triosy_obj_iswt0;
  output out_f_d_triosy_obj_biwt;



  // Interconnect Declarations for Component Instantiations 
  assign out_f_d_triosy_obj_biwt = (~ run_wten) & out_f_d_triosy_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_in_u_triosy_obj_in_u_triosy_wait_ctrl
// ------------------------------------------------------------------


module stage_run_in_u_triosy_obj_in_u_triosy_wait_ctrl (
  run_wten, in_u_triosy_obj_iswt0, in_u_triosy_obj_biwt
);
  input run_wten;
  input in_u_triosy_obj_iswt0;
  output in_u_triosy_obj_biwt;



  // Interconnect Declarations for Component Instantiations 
  assign in_u_triosy_obj_biwt = (~ run_wten) & in_u_triosy_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_in_f_d_triosy_obj_in_f_d_triosy_wait_ctrl
// ------------------------------------------------------------------


module stage_run_in_f_d_triosy_obj_in_f_d_triosy_wait_ctrl (
  run_wten, in_f_d_triosy_obj_iswt0, in_f_d_triosy_obj_biwt
);
  input run_wten;
  input in_f_d_triosy_obj_iswt0;
  output in_f_d_triosy_obj_biwt;



  // Interconnect Declarations for Component Instantiations 
  assign in_f_d_triosy_obj_biwt = (~ run_wten) & in_f_d_triosy_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_mode1_triosy_obj_mode1_triosy_wait_ctrl
// ------------------------------------------------------------------


module stage_run_mode1_triosy_obj_mode1_triosy_wait_ctrl (
  run_wten, mode1_triosy_obj_iswt0, mode1_triosy_obj_biwt
);
  input run_wten;
  input mode1_triosy_obj_iswt0;
  output mode1_triosy_obj_biwt;



  // Interconnect Declarations for Component Instantiations 
  assign mode1_triosy_obj_biwt = (~ run_wten) & mode1_triosy_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_out1_rsci_out1_wait_ctrl
// ------------------------------------------------------------------


module stage_run_out1_rsci_out1_wait_ctrl (
  out1_rsci_iswt0, out1_rsci_biwt, out1_rsci_irdy
);
  input out1_rsci_iswt0;
  output out1_rsci_biwt;
  input out1_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign out1_rsci_biwt = out1_rsci_iswt0 & out1_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_wait_dp
// ------------------------------------------------------------------


module stage_run_wait_dp (
  clk, rst, arst_n, in_f_d_rsci_en_d, in_u_rsci_en_d, out_f_d_rsci_en_d, out_u_rsci_en_d,
      BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en, BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en,
      BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en, BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en,
      r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en, BUTTERFLY_i_div_cmp_z,
      run_wen, in_f_d_rsci_cgo, in_f_d_rsci_cgo_ir_unreg, in_u_rsci_cgo, in_u_rsci_cgo_ir_unreg,
      out_f_d_rsci_cgo, out_f_d_rsci_cgo_ir_unreg, out_u_rsci_cgo, out_u_rsci_cgo_ir_unreg,
      BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo, BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo,
      BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo, BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo,
      r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_cgo, BUTTERFLY_i_div_cmp_z_oreg
);
  input clk;
  input rst;
  input arst_n;
  output in_f_d_rsci_en_d;
  output in_u_rsci_en_d;
  output out_f_d_rsci_en_d;
  output out_u_rsci_en_d;
  output BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en;
  output BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en;
  output BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en;
  output BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en;
  output r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en;
  input [15:0] BUTTERFLY_i_div_cmp_z;
  input run_wen;
  input in_f_d_rsci_cgo;
  input in_f_d_rsci_cgo_ir_unreg;
  input in_u_rsci_cgo;
  input in_u_rsci_cgo_ir_unreg;
  input out_f_d_rsci_cgo;
  input out_f_d_rsci_cgo_ir_unreg;
  input out_u_rsci_cgo;
  input out_u_rsci_cgo_ir_unreg;
  input BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo;
  input BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo;
  input BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo;
  input BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo;
  input r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_cgo;
  output [8:0] BUTTERFLY_i_div_cmp_z_oreg;


  // Interconnect Declarations
  reg [8:0] BUTTERFLY_i_div_cmp_z_oreg_pconst_8_0;


  // Interconnect Declarations for Component Instantiations 
  assign in_f_d_rsci_en_d = run_wen & (in_f_d_rsci_cgo | in_f_d_rsci_cgo_ir_unreg);
  assign in_u_rsci_en_d = run_wen & (in_u_rsci_cgo | in_u_rsci_cgo_ir_unreg);
  assign out_f_d_rsci_en_d = run_wen & (out_f_d_rsci_cgo | out_f_d_rsci_cgo_ir_unreg);
  assign out_u_rsci_en_d = run_wen & (out_u_rsci_cgo | out_u_rsci_cgo_ir_unreg);
  assign BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en = ~(run_wen & BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo);
  assign BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en = ~(run_wen & BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo);
  assign BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en = ~(run_wen & BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo);
  assign BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en = ~(run_wen & BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo);
  assign r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en = ~(run_wen &
      r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_cgo);
  assign BUTTERFLY_i_div_cmp_z_oreg = BUTTERFLY_i_div_cmp_z_oreg_pconst_8_0;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_i_div_cmp_z_oreg_pconst_8_0 <= 9'b000000000;
    end
    else if ( rst ) begin
      BUTTERFLY_i_div_cmp_z_oreg_pconst_8_0 <= 9'b000000000;
    end
    else if ( run_wen ) begin
      BUTTERFLY_i_div_cmp_z_oreg_pconst_8_0 <= BUTTERFLY_i_div_cmp_z[8:0];
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_ap_done_rsci_ap_done_wait_ctrl
// ------------------------------------------------------------------


module stage_run_ap_done_rsci_ap_done_wait_ctrl (
  ap_done_rsci_iswt0, ap_done_rsci_biwt, ap_done_rsci_irdy
);
  input ap_done_rsci_iswt0;
  output ap_done_rsci_biwt;
  input ap_done_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign ap_done_rsci_biwt = ap_done_rsci_iswt0 & ap_done_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_ap_start_rsci_ap_start_wait_ctrl
// ------------------------------------------------------------------


module stage_run_ap_start_rsci_ap_start_wait_ctrl (
  ap_start_rsci_iswt0, ap_start_rsci_biwt, ap_start_rsci_ivld
);
  input ap_start_rsci_iswt0;
  output ap_start_rsci_biwt;
  input ap_start_rsci_ivld;



  // Interconnect Declarations for Component Instantiations 
  assign ap_start_rsci_biwt = ap_start_rsci_iswt0 & ap_start_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_out_u_triosy_obj
// ------------------------------------------------------------------


module stage_run_out_u_triosy_obj (
  out_u_triosy_lz, run_wten, out_u_triosy_obj_iswt0
);
  output out_u_triosy_lz;
  input run_wten;
  input out_u_triosy_obj_iswt0;


  // Interconnect Declarations
  wire out_u_triosy_obj_biwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) out_u_triosy_obj (
      .ld(out_u_triosy_obj_biwt),
      .lz(out_u_triosy_lz)
    );
  stage_run_out_u_triosy_obj_out_u_triosy_wait_ctrl stage_run_out_u_triosy_obj_out_u_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .out_u_triosy_obj_iswt0(out_u_triosy_obj_iswt0),
      .out_u_triosy_obj_biwt(out_u_triosy_obj_biwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_out_f_d_triosy_obj
// ------------------------------------------------------------------


module stage_run_out_f_d_triosy_obj (
  out_f_d_triosy_lz, run_wten, out_f_d_triosy_obj_iswt0
);
  output out_f_d_triosy_lz;
  input run_wten;
  input out_f_d_triosy_obj_iswt0;


  // Interconnect Declarations
  wire out_f_d_triosy_obj_biwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) out_f_d_triosy_obj (
      .ld(out_f_d_triosy_obj_biwt),
      .lz(out_f_d_triosy_lz)
    );
  stage_run_out_f_d_triosy_obj_out_f_d_triosy_wait_ctrl stage_run_out_f_d_triosy_obj_out_f_d_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .out_f_d_triosy_obj_iswt0(out_f_d_triosy_obj_iswt0),
      .out_f_d_triosy_obj_biwt(out_f_d_triosy_obj_biwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_in_u_triosy_obj
// ------------------------------------------------------------------


module stage_run_in_u_triosy_obj (
  in_u_triosy_lz, run_wten, in_u_triosy_obj_iswt0
);
  output in_u_triosy_lz;
  input run_wten;
  input in_u_triosy_obj_iswt0;


  // Interconnect Declarations
  wire in_u_triosy_obj_biwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) in_u_triosy_obj (
      .ld(in_u_triosy_obj_biwt),
      .lz(in_u_triosy_lz)
    );
  stage_run_in_u_triosy_obj_in_u_triosy_wait_ctrl stage_run_in_u_triosy_obj_in_u_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .in_u_triosy_obj_iswt0(in_u_triosy_obj_iswt0),
      .in_u_triosy_obj_biwt(in_u_triosy_obj_biwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_in_f_d_triosy_obj
// ------------------------------------------------------------------


module stage_run_in_f_d_triosy_obj (
  in_f_d_triosy_lz, run_wten, in_f_d_triosy_obj_iswt0
);
  output in_f_d_triosy_lz;
  input run_wten;
  input in_f_d_triosy_obj_iswt0;


  // Interconnect Declarations
  wire in_f_d_triosy_obj_biwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) in_f_d_triosy_obj (
      .ld(in_f_d_triosy_obj_biwt),
      .lz(in_f_d_triosy_lz)
    );
  stage_run_in_f_d_triosy_obj_in_f_d_triosy_wait_ctrl stage_run_in_f_d_triosy_obj_in_f_d_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .in_f_d_triosy_obj_iswt0(in_f_d_triosy_obj_iswt0),
      .in_f_d_triosy_obj_biwt(in_f_d_triosy_obj_biwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_mode1_triosy_obj
// ------------------------------------------------------------------


module stage_run_mode1_triosy_obj (
  mode1_triosy_lz, run_wten, mode1_triosy_obj_iswt0
);
  output mode1_triosy_lz;
  input run_wten;
  input mode1_triosy_obj_iswt0;


  // Interconnect Declarations
  wire mode1_triosy_obj_biwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) mode1_triosy_obj (
      .ld(mode1_triosy_obj_biwt),
      .lz(mode1_triosy_lz)
    );
  stage_run_mode1_triosy_obj_mode1_triosy_wait_ctrl stage_run_mode1_triosy_obj_mode1_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .mode1_triosy_obj_iswt0(mode1_triosy_obj_iswt0),
      .mode1_triosy_obj_biwt(mode1_triosy_obj_biwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_out1_rsci
// ------------------------------------------------------------------


module stage_run_out1_rsci (
  out1_rsc_dat, out1_rsc_vld, out1_rsc_rdy, out1_rsci_oswt, out1_rsci_wen_comp, out1_rsci_idat
);
  output [79:0] out1_rsc_dat;
  output out1_rsc_vld;
  input out1_rsc_rdy;
  input out1_rsci_oswt;
  output out1_rsci_wen_comp;
  input [79:0] out1_rsci_idat;


  // Interconnect Declarations
  wire out1_rsci_biwt;
  wire out1_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd8),
  .width(32'sd80)) out1_rsci (
      .irdy(out1_rsci_irdy),
      .ivld(out1_rsci_oswt),
      .idat(out1_rsci_idat),
      .rdy(out1_rsc_rdy),
      .vld(out1_rsc_vld),
      .dat(out1_rsc_dat)
    );
  stage_run_out1_rsci_out1_wait_ctrl stage_run_out1_rsci_out1_wait_ctrl_inst (
      .out1_rsci_iswt0(out1_rsci_oswt),
      .out1_rsci_biwt(out1_rsci_biwt),
      .out1_rsci_irdy(out1_rsci_irdy)
    );
  assign out1_rsci_wen_comp = (~ out1_rsci_oswt) | out1_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_ap_done_rsci
// ------------------------------------------------------------------


module stage_run_ap_done_rsci (
  ap_done_rsc_dat, ap_done_rsc_vld, ap_done_rsc_rdy, ap_done_rsci_oswt, ap_done_rsci_wen_comp
);
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input ap_done_rsci_oswt;
  output ap_done_rsci_wen_comp;


  // Interconnect Declarations
  wire ap_done_rsci_biwt;
  wire ap_done_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd1)) ap_done_rsci (
      .irdy(ap_done_rsci_irdy),
      .ivld(ap_done_rsci_oswt),
      .idat(1'b1),
      .rdy(ap_done_rsc_rdy),
      .vld(ap_done_rsc_vld),
      .dat(ap_done_rsc_dat)
    );
  stage_run_ap_done_rsci_ap_done_wait_ctrl stage_run_ap_done_rsci_ap_done_wait_ctrl_inst
      (
      .ap_done_rsci_iswt0(ap_done_rsci_oswt),
      .ap_done_rsci_biwt(ap_done_rsci_biwt),
      .ap_done_rsci_irdy(ap_done_rsci_irdy)
    );
  assign ap_done_rsci_wen_comp = (~ ap_done_rsci_oswt) | ap_done_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_ap_start_rsci
// ------------------------------------------------------------------


module stage_run_ap_start_rsci (
  ap_start_rsc_dat, ap_start_rsc_vld, ap_start_rsc_rdy, ap_start_rsci_oswt, ap_start_rsci_wen_comp
);
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  input ap_start_rsci_oswt;
  output ap_start_rsci_wen_comp;


  // Interconnect Declarations
  wire ap_start_rsci_biwt;
  wire ap_start_rsci_ivld;
  wire ap_start_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd1)) ap_start_rsci (
      .rdy(ap_start_rsc_rdy),
      .vld(ap_start_rsc_vld),
      .dat(ap_start_rsc_dat),
      .irdy(ap_start_rsci_oswt),
      .ivld(ap_start_rsci_ivld),
      .idat(ap_start_rsci_idat)
    );
  stage_run_ap_start_rsci_ap_start_wait_ctrl stage_run_ap_start_rsci_ap_start_wait_ctrl_inst
      (
      .ap_start_rsci_iswt0(ap_start_rsci_oswt),
      .ap_start_rsci_biwt(ap_start_rsci_biwt),
      .ap_start_rsci_ivld(ap_start_rsci_ivld)
    );
  assign ap_start_rsci_wen_comp = (~ ap_start_rsci_oswt) | ap_start_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run
// ------------------------------------------------------------------


module stage_run (
  clk, rst, arst_n, ap_start_rsc_dat, ap_start_rsc_vld, ap_start_rsc_rdy, ap_done_rsc_dat,
      ap_done_rsc_vld, ap_done_rsc_rdy, mode1_rsc_dat, mode1_triosy_lz, in_f_d_triosy_lz,
      in_u_triosy_lz, out_f_d_triosy_lz, out_u_triosy_lz, out1_rsc_dat, out1_rsc_vld,
      out1_rsc_rdy, in_f_d_rsci_adr_d, in_f_d_rsci_d_d, in_f_d_rsci_en_d, in_f_d_rsci_q_d,
      in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, in_u_rsci_adr_d, in_u_rsci_d_d,
      in_u_rsci_en_d, in_u_rsci_q_d, in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      out_f_d_rsci_adr_d, out_f_d_rsci_d_d, out_f_d_rsci_en_d, out_f_d_rsci_q_d,
      out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, out_u_rsci_adr_d, out_u_rsci_d_d,
      out_u_rsci_en_d, out_u_rsci_q_d, out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr, BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out,
      BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en, BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out,
      BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en, BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out,
      BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en, BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out,
      BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en, r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out,
      r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en, BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out,
      BUTTERFLY_i_div_cmp_a, BUTTERFLY_i_div_cmp_b, BUTTERFLY_i_div_cmp_z, in_f_d_rsci_we_d_pff,
      in_u_rsci_we_d_pff, out_f_d_rsci_we_d_pff, out_u_rsci_we_d_pff
);
  input clk;
  input rst;
  input arst_n;
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input [15:0] mode1_rsc_dat;
  output mode1_triosy_lz;
  output in_f_d_triosy_lz;
  output in_u_triosy_lz;
  output out_f_d_triosy_lz;
  output out_u_triosy_lz;
  output [79:0] out1_rsc_dat;
  output out1_rsc_vld;
  input out1_rsc_rdy;
  output [9:0] in_f_d_rsci_adr_d;
  output [63:0] in_f_d_rsci_d_d;
  output in_f_d_rsci_en_d;
  input [63:0] in_f_d_rsci_q_d;
  output in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [9:0] in_u_rsci_adr_d;
  output [15:0] in_u_rsci_d_d;
  output in_u_rsci_en_d;
  input [15:0] in_u_rsci_q_d;
  output in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [9:0] out_f_d_rsci_adr_d;
  output [63:0] out_f_d_rsci_d_d;
  output out_f_d_rsci_en_d;
  input [63:0] out_f_d_rsci_q_d;
  output out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [9:0] out_u_rsci_adr_d;
  output [15:0] out_u_rsci_d_d;
  output out_u_rsci_en_d;
  input [15:0] out_u_rsci_q_d;
  output out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [9:0] BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr;
  input [13:0] BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out;
  output BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en;
  input [13:0] BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out;
  output BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en;
  input [13:0] BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out;
  output BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en;
  input [13:0] BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out;
  output BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en;
  input [61:0] r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out;
  output r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en;
  input [63:0] BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out;
  output [15:0] BUTTERFLY_i_div_cmp_a;
  output [15:0] BUTTERFLY_i_div_cmp_b;
  input [15:0] BUTTERFLY_i_div_cmp_z;
  output in_f_d_rsci_we_d_pff;
  output in_u_rsci_we_d_pff;
  output out_f_d_rsci_we_d_pff;
  output out_u_rsci_we_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire ap_start_rsci_wen_comp;
  wire ap_done_rsci_wen_comp;
  wire [15:0] mode1_rsci_idat;
  wire out1_rsci_wen_comp;
  reg BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo;
  reg BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo;
  reg BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo;
  reg BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo;
  wire [8:0] BUTTERFLY_i_div_cmp_z_oreg;
  reg [15:0] out1_rsci_idat_79_64;
  wire [38:0] fsm_output;
  wire return_add_generic_AC_RND_CONV_false_11_if_5_return_add_generic_AC_RND_CONV_false_11_if_5_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_10_if_5_return_add_generic_AC_RND_CONV_false_10_if_5_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_10_else_4_return_add_generic_AC_RND_CONV_false_10_else_4_nand_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_10_e_dif1_acc_1_tmp;
  wire [12:0] nl_return_add_generic_AC_RND_CONV_false_10_e_dif1_acc_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_9_e_dif1_acc_1_tmp;
  wire [12:0] nl_return_add_generic_AC_RND_CONV_false_9_e_dif1_acc_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_9_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_8_if_5_return_add_generic_AC_RND_CONV_false_8_if_5_and_tmp;
  wire return_extract_22_and_1_tmp;
  wire [53:0] return_add_generic_AC_RND_CONV_false_7_res_rounded_acc_tmp;
  wire [54:0] nl_return_add_generic_AC_RND_CONV_false_7_res_rounded_acc_tmp;
  wire [12:0] return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp;
  wire [14:0] nl_return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp;
  wire return_extract_19_return_extract_19_nor_tmp;
  wire return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp;
  wire operator_11_true_19_operator_11_true_19_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_tmp;
  wire [12:0] operator_33_true_12_acc_tmp;
  wire [13:0] nl_operator_33_true_12_acc_tmp;
  wire return_extract_17_and_tmp;
  wire return_extract_16_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp;
  wire return_extract_12_return_extract_12_or_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_2_if_5_return_add_generic_AC_RND_CONV_false_2_if_5_and_1_tmp;
  wire [53:0] return_add_generic_AC_RND_CONV_false_2_res_rounded_acc_tmp;
  wire [54:0] nl_return_add_generic_AC_RND_CONV_false_2_res_rounded_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_2_else_4_return_add_generic_AC_RND_CONV_false_2_else_4_nand_tmp;
  wire [12:0] operator_33_true_4_acc_tmp;
  wire [13:0] nl_operator_33_true_4_acc_tmp;
  wire [53:0] return_add_generic_AC_RND_CONV_false_res_rounded_acc_tmp;
  wire [54:0] nl_return_add_generic_AC_RND_CONV_false_res_rounded_acc_tmp;
  wire [12:0] return_mult_generic_AC_RND_CONV_false_1_exp_acc_tmp;
  wire [14:0] nl_return_mult_generic_AC_RND_CONV_false_1_exp_acc_tmp;
  wire return_extract_17_return_extract_17_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_1_return_add_generic_AC_RND_CONV_false_6_op2_normal_return_extract_13_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_1_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_25_if_5_return_add_generic_AC_RND_CONV_false_25_if_5_and_tmp;
  wire [53:0] return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp;
  wire [54:0] nl_return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_25_else_4_return_add_generic_AC_RND_CONV_false_25_else_4_nand_tmp;
  wire [12:0] operator_33_true_50_acc_tmp;
  wire [13:0] nl_operator_33_true_50_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_24_if_5_return_add_generic_AC_RND_CONV_false_24_if_5_and_tmp;
  wire [53:0] return_add_generic_AC_RND_CONV_false_24_res_rounded_acc_tmp;
  wire [54:0] nl_return_add_generic_AC_RND_CONV_false_24_res_rounded_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_24_else_4_return_add_generic_AC_RND_CONV_false_24_else_4_nand_tmp;
  wire [12:0] operator_33_true_48_acc_tmp;
  wire [13:0] nl_operator_33_true_48_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_23_if_5_return_add_generic_AC_RND_CONV_false_23_if_5_and_tmp;
  wire [53:0] return_add_generic_AC_RND_CONV_false_23_res_rounded_acc_tmp;
  wire [54:0] nl_return_add_generic_AC_RND_CONV_false_23_res_rounded_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_23_else_4_return_add_generic_AC_RND_CONV_false_23_else_4_nand_tmp;
  wire [12:0] operator_33_true_46_acc_tmp;
  wire [13:0] nl_operator_33_true_46_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_22_if_5_return_add_generic_AC_RND_CONV_false_22_if_5_and_1_tmp;
  wire [12:0] operator_33_true_44_acc_tmp;
  wire [13:0] nl_operator_33_true_44_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_23_e_dif1_acc_1_tmp;
  wire [12:0] nl_return_add_generic_AC_RND_CONV_false_23_e_dif1_acc_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_23_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_22_e_dif1_acc_1_tmp;
  wire [12:0] nl_return_add_generic_AC_RND_CONV_false_22_e_dif1_acc_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_22_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_21_if_5_return_add_generic_AC_RND_CONV_false_21_if_5_and_tmp;
  wire [53:0] return_add_generic_AC_RND_CONV_false_21_res_rounded_acc_tmp;
  wire [54:0] nl_return_add_generic_AC_RND_CONV_false_21_res_rounded_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_21_else_4_return_add_generic_AC_RND_CONV_false_21_else_4_nand_tmp;
  wire return_add_generic_AC_RND_CONV_false_20_if_5_return_add_generic_AC_RND_CONV_false_20_if_5_and_1_tmp;
  wire [53:0] return_add_generic_AC_RND_CONV_false_20_res_rounded_acc_tmp;
  wire [54:0] nl_return_add_generic_AC_RND_CONV_false_20_res_rounded_acc_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp;
  wire [12:0] nl_return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp;
  wire return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp;
  wire [12:0] nl_return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp;
  wire return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp;
  wire [12:0] return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp;
  wire [14:0] nl_return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp;
  wire return_extract_51_return_extract_51_nor_tmp;
  wire return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp;
  wire operator_11_true_51_operator_11_true_51_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_19_if_5_return_add_generic_AC_RND_CONV_false_19_if_5_and_tmp;
  wire [53:0] return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp;
  wire [54:0] nl_return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp;
  wire return_mult_generic_AC_RND_CONV_false_3_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_3_exp_ovf_oif_aelse_and_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp;
  wire return_extract_44_return_extract_44_or_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_15_if_5_return_add_generic_AC_RND_CONV_false_15_if_5_and_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_15_else_4_return_add_generic_AC_RND_CONV_false_15_else_4_nand_tmp;
  wire return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp;
  wire return_mult_generic_AC_RND_CONV_false_4_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_4_exp_ovf_oif_aelse_and_tmp;
  wire return_extract_49_return_extract_49_nor_tmp;
  wire return_extract_49_m_zero_return_extract_49_m_zero_nor_tmp;
  wire operator_11_true_49_operator_11_true_49_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_tmp;
  wire [53:0] return_add_generic_AC_RND_CONV_false_18_res_rounded_acc_tmp;
  wire [54:0] nl_return_add_generic_AC_RND_CONV_false_18_res_rounded_acc_tmp;
  wire [53:0] return_add_generic_AC_RND_CONV_false_17_res_rounded_acc_tmp;
  wire [54:0] nl_return_add_generic_AC_RND_CONV_false_17_res_rounded_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_if_1_return_add_generic_AC_RND_CONV_false_17_op2_normal_return_extract_41_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_or_tmp;
  wire [10:0] return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp;
  wire [11:0] nl_return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_17_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_14_e1_eq_e2_equal_tmp;
  wire stage_PE_1_and_1_tmp;
  wire operator_16_false_operator_16_false_nor_tmp;
  wire or_dcpl_3;
  wire nor_tmp;
  wire and_dcpl_1;
  wire or_dcpl_25;
  wire or_dcpl_35;
  wire and_dcpl_35;
  wire and_dcpl_42;
  wire and_dcpl_44;
  wire or_dcpl_60;
  wire and_dcpl_74;
  wire and_dcpl_80;
  wire and_dcpl_83;
  wire or_dcpl_64;
  wire or_dcpl_65;
  wire or_dcpl_69;
  wire or_dcpl_75;
  wire or_dcpl_77;
  wire and_dcpl_85;
  wire and_dcpl_91;
  wire or_dcpl_82;
  wire or_dcpl_83;
  wire or_dcpl_85;
  wire or_dcpl_86;
  wire or_dcpl_87;
  wire or_dcpl_88;
  wire or_dcpl_89;
  wire or_dcpl_92;
  wire or_dcpl_98;
  wire or_dcpl_99;
  wire or_dcpl_101;
  wire or_dcpl_102;
  wire or_dcpl_104;
  wire or_dcpl_106;
  wire or_dcpl_107;
  wire or_dcpl_109;
  wire or_dcpl_111;
  wire and_dcpl_110;
  wire or_dcpl_124;
  wire or_dcpl_125;
  wire or_dcpl_133;
  wire or_dcpl_145;
  wire or_dcpl_147;
  wire or_dcpl_151;
  wire and_dcpl_112;
  wire or_dcpl_152;
  wire or_dcpl_153;
  wire or_dcpl_158;
  wire or_dcpl_159;
  wire and_dcpl_114;
  wire or_dcpl_164;
  wire or_dcpl_167;
  wire or_dcpl_168;
  wire or_dcpl_172;
  wire and_dcpl_118;
  wire and_dcpl_121;
  wire or_dcpl_183;
  wire or_dcpl_190;
  wire and_dcpl_125;
  wire or_dcpl_193;
  wire or_dcpl_198;
  wire and_dcpl_127;
  wire or_dcpl_201;
  wire and_dcpl_129;
  wire or_dcpl_212;
  wire and_dcpl_131;
  wire and_dcpl_132;
  wire or_dcpl_238;
  wire and_dcpl_133;
  wire or_dcpl_245;
  wire and_dcpl_135;
  wire or_dcpl_250;
  wire and_dcpl_136;
  wire and_dcpl_139;
  wire and_dcpl_141;
  wire and_dcpl_143;
  wire and_dcpl_147;
  wire and_dcpl_149;
  wire and_dcpl_150;
  wire and_dcpl_164;
  wire or_dcpl_300;
  wire or_dcpl_305;
  wire and_dcpl_170;
  wire and_dcpl_179;
  wire or_dcpl_316;
  wire or_dcpl_320;
  wire or_dcpl_325;
  wire or_dcpl_326;
  wire or_dcpl_328;
  wire and_dcpl_196;
  wire and_dcpl_197;
  wire or_dcpl_338;
  wire or_dcpl_340;
  wire or_dcpl_343;
  wire or_dcpl_352;
  wire or_dcpl_353;
  wire or_dcpl_354;
  wire or_dcpl_356;
  wire or_dcpl_357;
  wire or_dcpl_358;
  wire or_dcpl_359;
  wire or_dcpl_360;
  wire or_dcpl_361;
  wire or_dcpl_365;
  wire or_dcpl_367;
  wire or_dcpl_377;
  wire or_dcpl_380;
  wire or_dcpl_385;
  wire or_dcpl_387;
  wire or_dcpl_388;
  wire or_dcpl_390;
  wire or_dcpl_396;
  wire and_dcpl_214;
  wire and_dcpl_215;
  wire and_dcpl_216;
  wire and_dcpl_219;
  wire and_dcpl_220;
  wire and_dcpl_224;
  wire or_dcpl_432;
  wire and_dcpl_225;
  wire or_dcpl_436;
  wire or_dcpl_437;
  wire and_dcpl_226;
  wire and_dcpl_227;
  wire or_dcpl_441;
  wire and_dcpl_228;
  wire or_dcpl_442;
  wire or_dcpl_443;
  wire and_dcpl_229;
  wire and_dcpl_231;
  wire or_dcpl_450;
  wire or_dcpl_454;
  wire or_dcpl_456;
  wire and_dcpl_241;
  wire or_dcpl_471;
  wire or_dcpl_474;
  wire or_dcpl_475;
  wire or_dcpl_477;
  wire or_dcpl_480;
  wire or_dcpl_488;
  wire or_dcpl_505;
  wire or_dcpl_511;
  wire or_dcpl_523;
  wire and_dcpl_248;
  wire and_dcpl_249;
  wire and_dcpl_254;
  wire and_dcpl_281;
  wire or_dcpl_551;
  wire or_dcpl_571;
  wire and_dcpl_294;
  wire and_dcpl_300;
  wire or_dcpl_597;
  wire and_dcpl_312;
  wire and_dcpl_314;
  wire and_dcpl_316;
  wire or_dcpl_625;
  wire or_tmp_26;
  wire or_tmp_46;
  wire or_tmp_180;
  wire or_tmp_181;
  wire or_tmp_388;
  wire or_tmp_389;
  wire or_tmp_543;
  wire or_tmp_567;
  wire or_tmp_606;
  wire or_tmp_773;
  wire and_421_cse;
  wire and_450_cse;
  wire and_448_cse;
  wire and_477_cse;
  wire and_475_cse;
  wire and_392_cse;
  wire and_503_cse;
  wire and_539_cse;
  wire and_537_cse;
  wire and_565_cse;
  wire and_569_cse;
  wire and_573_cse;
  wire and_631_cse;
  wire and_1747_cse;
  wire return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_6_lor_lpi_2_dfm_1;
  wire return_extract_3_m_zero_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_6_op1_nan_sva_1;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3;
  wire return_mult_generic_AC_RND_CONV_false_6_e_incr_lpi_2_dfm_2;
  wire return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_or_2;
  wire return_add_generic_AC_RND_CONV_false_12_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  wire return_add_generic_AC_RND_CONV_false_7_if_5_or_3;
  reg operator_11_true_return_13_sva;
  reg return_add_generic_AC_RND_CONV_false_10_op2_inf_sva;
  reg operator_11_true_return_15_sva;
  reg return_add_generic_AC_RND_CONV_false_10_op2_nan_sva;
  reg return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm;
  wire return_add_generic_AC_RND_CONV_false_11_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva;
  reg return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva;
  wire return_add_generic_AC_RND_CONV_false_6_if_5_or_3;
  reg operator_11_true_return_1_sva;
  reg operator_11_true_return_24_sva;
  reg operator_11_true_return_17_sva;
  reg return_add_generic_AC_RND_CONV_false_15_do_sub_sva;
  wire return_add_generic_AC_RND_CONV_false_11_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp;
  wire [5:0] operator_6_false_10_operator_6_false_10_conc_2_6_1;
  wire [6:0] nl_operator_6_false_10_operator_6_false_10_conc_2_6_1;
  wire return_add_generic_AC_RND_CONV_false_10_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_10_op1_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_10_op1_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1;
  reg operator_11_true_return_26_sva;
  reg return_extract_44_m_zero_sva;
  reg [9:0] return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_itm;
  reg return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm;
  wire return_add_generic_AC_RND_CONV_false_9_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_9_op1_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_7_op1_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_9_op1_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_7_op1_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_9_r_inf_lpi_3_dfm_2;
  reg return_extract_1_m_zero_sva;
  wire [11:0] return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm_mx1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_mx0w4;
  wire return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_9_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_8_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_8_if_5_or_3;
  wire return_add_generic_AC_RND_CONV_false_8_op1_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_8_r_inf_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_7_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2;
  reg return_extract_15_m_zero_sva;
  reg return_extract_12_m_zero_sva;
  wire operator_11_true_return_15_sva_mx1;
  wire return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1;
  reg return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm;
  reg drf_qr_lval_14_smx_0_lpi_3_dfm;
  reg [49:0] return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm;
  wire return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_8_e_dif_qr_lpi_3_dfm_mx0;
  reg return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm;
  reg return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm;
  wire return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_7_e_dif_qr_lpi_3_dfm_mx0;
  wire return_mult_generic_AC_RND_CONV_false_2_zero_m_return_mult_generic_AC_RND_CONV_false_2_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_2_r_zero_return_mult_generic_AC_RND_CONV_false_2_r_zero_nor_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_2_lor_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_2_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_2_r_nan_sva_1;
  reg return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1;
  wire [11:0] return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_2_e_incr_lpi_3_dfm_2;
  wire [105:0] return_mult_generic_AC_RND_CONV_false_2_p_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_or_2;
  wire [105:0] return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_2_if_nor_ovfl_sva_1;
  wire return_add_generic_AC_RND_CONV_false_6_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2;
  wire [50:0] return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_3_exp_ovf_lor_lpi_3_dfm_2;
  wire return_mult_generic_AC_RND_CONV_false_zero_m_return_mult_generic_AC_RND_CONV_false_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_r_zero_return_mult_generic_AC_RND_CONV_false_r_zero_nor_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_lor_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_r_nan_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_op1_zero_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_op2_zero_sva_1;
  reg return_extract_15_return_extract_15_nor_cse_sva;
  wire return_add_generic_AC_RND_CONV_false_6_op1_mu_0_lpi_3_dfm_1;
  reg return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50;
  reg return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm;
  reg [49:0] return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0;
  wire return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_1_zero_m_return_mult_generic_AC_RND_CONV_false_1_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_1_r_zero_return_mult_generic_AC_RND_CONV_false_1_r_zero_nor_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_1_lor_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_1_r_nan_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_or_2;
  reg [5:0] return_add_generic_AC_RND_CONV_false_20_ls_sva;
  wire return_add_generic_AC_RND_CONV_false_14_op2_nan_sva_1;
  reg stage_PE_1_tmp_im_d_1_lpi_3_dfm_63;
  wire [50:0] stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0;
  wire return_add_generic_AC_RND_CONV_false_2_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_op1_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_op2_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_op1_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_op2_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_exception_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_1_if_nor_ovfl_sva_1;
  wire return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_4_m_r_51_lpi_3_dfm_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_mx0w2;
  wire [11:0] operator_33_true_10_acc_psp_1_sva_1;
  wire [12:0] nl_operator_33_true_10_acc_psp_1_sva_1;
  wire return_add_generic_AC_RND_CONV_false_do_sub_sva_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_e_dif_qr_lpi_3_dfm_mx0;
  wire stage_PE_tmp_im_d_1_lpi_3_dfm_51_mx0;
  wire [50:0] stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0;
  wire [56:0] return_add_generic_AC_RND_CONV_false_5_res_mant_4_sva_1;
  wire [58:0] nl_return_add_generic_AC_RND_CONV_false_5_res_mant_4_sva_1;
  wire [56:0] return_add_generic_AC_RND_CONV_false_4_res_mant_4_sva_1;
  wire [58:0] nl_return_add_generic_AC_RND_CONV_false_4_res_mant_4_sva_1;
  wire return_add_generic_AC_RND_CONV_false_3_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_14_op1_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_14_op1_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_1_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_1_r_inf_lpi_3_dfm_2;
  reg inverse_lpi_1_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_1_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_25_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_23_op1_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_23_op1_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_25_r_inf_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_24_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_22_op1_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_22_op1_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_24_r_inf_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_23_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_23_r_inf_lpi_3_dfm_2;
  reg return_extract_17_m_zero_sva;
  wire return_add_generic_AC_RND_CONV_false_22_exception_sva_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm_mx2;
  wire [50:0] return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_mx0w6;
  wire return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_21_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_21_op1_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_21_op1_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_20_exception_sva_1;
  wire operator_11_true_return_15_sva_mx2;
  wire return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2;
  wire return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1;
  wire [10:0] drf_qr_lval_26_smx_lpi_3_dfm_mx0;
  reg return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm;
  wire return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_5_zero_m_return_mult_generic_AC_RND_CONV_false_5_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_5_r_zero_return_mult_generic_AC_RND_CONV_false_5_r_zero_nor_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_5_lor_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_5_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_5_r_nan_sva_1;
  wire [105:0] return_mult_generic_AC_RND_CONV_false_5_p_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_or_2;
  wire [105:0] return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_5_if_nor_ovfl_sva_1;
  wire return_add_generic_AC_RND_CONV_false_19_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_19_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp;
  wire BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx3;
  wire [50:0] return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_3_zero_m_return_mult_generic_AC_RND_CONV_false_3_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_3_r_zero_return_mult_generic_AC_RND_CONV_false_3_r_zero_nor_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_3_lor_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_3_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_3_r_nan_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_4_op1_zero_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_3_op2_zero_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1;
  wire return_add_generic_AC_RND_CONV_false_19_op1_mu_0_lpi_3_dfm_1;
  reg return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm;
  wire stage_PE_1_tmp_re_d_1_lpi_3_dfm_63_mx1;
  wire stage_PE_1_tmp_re_d_1_lpi_3_dfm_51_mx1;
  wire [50:0] stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1;
  wire return_add_generic_AC_RND_CONV_false_15_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_13_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx6;
  wire [50:0] return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_4_zero_m_return_mult_generic_AC_RND_CONV_false_4_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_4_r_zero_return_mult_generic_AC_RND_CONV_false_4_r_zero_nor_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_4_lor_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_4_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_4_r_nan_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_4_op2_zero_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_or_2;
  reg return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_cse_sva;
  reg return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_and_1_itm;
  reg return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm;
  wire [50:0] return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_mx0w5;
  wire return_add_generic_AC_RND_CONV_false_13_do_sub_sva_1;
  wire stage_PE_1_tmp_im_d_1_lpi_3_dfm_51_mx1;
  wire [50:0] stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx1;
  wire [11:0] operator_33_true_34_acc_psp_1_sva_1;
  wire [12:0] nl_operator_33_true_34_acc_psp_1_sva_1;
  wire return_add_generic_AC_RND_CONV_false_16_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_14_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_5_do_sub_sva_1;
  wire return_add_generic_AC_RND_CONV_false_4_do_sub_sva_1;
  wire return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1;
  wire operator_16_false_1_operator_16_false_1_and_mdf_sva_1;
  reg operator_16_false_operator_16_false_nor_cse_sva;
  reg BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm;
  reg mode_lpi_1_dfm;
  reg [3:0] for_i_3_0_sva;
  reg [15:0] operator_16_false_io_read_mode1_rsc_cse_sva;
  reg return_add_generic_AC_RND_CONV_false_12_mux_itm;
  reg return_add_generic_AC_RND_CONV_false_12_do_sub_sva;
  reg return_add_generic_AC_RND_CONV_false_10_do_sub_sva;
  reg return_add_generic_AC_RND_CONV_false_21_unequal_tmp;
  reg return_add_generic_AC_RND_CONV_false_13_do_sub_sva;
  wire [11:0] operator_6_false_58_acc_psp_sva_1;
  wire [12:0] nl_operator_6_false_58_acc_psp_sva_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0w1;
  wire [12:0] nl_return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0w1;
  wire [12:0] operator_6_false_16_acc_psp_sva_1;
  wire [13:0] nl_operator_6_false_16_acc_psp_sva_1;
  wire [12:0] operator_6_false_45_acc_psp_sva_1;
  wire [13:0] nl_operator_6_false_45_acc_psp_sva_1;
  wire operator_11_true_return_3_sva_mx1w0;
  reg return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva;
  reg drf_qr_lval_12_smx_0_lpi_3_dfm;
  wire return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm_mx1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_mx0w2;
  wire [9:0] return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1;
  reg [63:0] stage_PE_1_x_im_d_sva;
  reg [63:0] stage_PE_1_x_re_d_sva;
  wire [50:0] return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1;
  reg return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva;
  wire stage_d_mul_return_d_1_63_sva_1;
  wire stage_d_mul_return_d_2_63_sva_1;
  wire stage_d_mul_return_d_63_sva_1;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1;
  reg return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w3;
  reg return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva;
  wire stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx1_50;
  wire [9:0] return_add_generic_AC_RND_CONV_false_4_e_r_qelse_qr_10_1_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_mx1w0;
  wire [9:0] return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1;
  reg return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva;
  wire stage_d_mul_return_d_5_63_sva_1;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_3_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w7;
  reg return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva;
  wire [105:0] return_mult_generic_AC_RND_CONV_false_3_p_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_if_1_aelse_return_mult_generic_AC_RND_CONV_false_if_1_aelse_or_2;
  wire stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx2_50;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_4_exp_1_11_0_lpi_3_dfm_3_10_0_1;
  reg return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva;
  reg return_add_generic_AC_RND_CONV_false_11_mux_itm;
  reg reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd;
  reg [49:0] reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1;
  wire for_1_if_and_ssc;
  reg out1_rsci_idat_63;
  reg [10:0] out1_rsci_idat_62_52;
  reg out1_rsci_idat_51;
  reg [50:0] out1_rsci_idat_50_0;
  wire [11:0] return_add_generic_AC_RND_CONV_false_12_e_dif_qif_acc_1_sdt;
  wire [12:0] nl_return_add_generic_AC_RND_CONV_false_12_e_dif_qif_acc_1_sdt;
  wire [11:0] return_add_generic_AC_RND_CONV_false_11_e_dif_qif_acc_1_sdt;
  wire [12:0] nl_return_add_generic_AC_RND_CONV_false_11_e_dif_qif_acc_1_sdt;
  wire [9:0] stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_1;
  wire stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_2_e_dif_qr_lpi_3_dfm_mx0_10_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt;
  wire [11:0] nl_return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt;
  wire [9:0] return_add_generic_AC_RND_CONV_false_4_e_dif_qif_acc_pmx_lpi_3_dfm_mx0_9_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_3_e_dif_qr_lpi_3_dfm_mx0_10_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_25_e_dif_qr_lpi_3_dfm_mx0_10_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_24_e_dif_qr_lpi_3_dfm_mx0_10_0;
  wire [9:0] stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx1_10_1;
  wire stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx1_0;
  wire [9:0] stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_1;
  wire stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0;
  wire [9:0] stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_1;
  wire stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0;
  reg reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_cgo_cse;
  reg reg_out_u_triosy_obj_iswt0_cse;
  reg reg_out1_rsci_iswt0_cse;
  reg reg_out_u_rsci_cgo_ir_cse;
  reg reg_out_f_d_rsci_cgo_ir_cse;
  reg reg_in_u_rsci_cgo_ir_cse;
  reg reg_in_f_d_rsci_cgo_ir_cse;
  reg reg_ap_start_rsci_iswt0_cse;
  reg [9:0] reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_addr_cse;
  wire [10:0] nl_reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_addr_cse;
  wire operator_16_false_and_cse;
  wire t_in_and_cse;
  wire mode_and_cse;
  wire stage_PE_1_and_2_cse;
  wire return_extract_41_and_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op1_smaller_return_add_generic_AC_RND_CONV_false_11_op1_smaller_or_cse;
  wire return_add_generic_AC_RND_CONV_false_24_op1_smaller_return_add_generic_AC_RND_CONV_false_24_op1_smaller_or_cse;
  wire return_add_generic_AC_RND_CONV_false_25_op1_smaller_return_add_generic_AC_RND_CONV_false_25_op1_smaller_or_cse;
  wire and_336_cse;
  wire and_178_cse;
  wire or_451_cse;
  wire return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse;
  wire return_add_generic_AC_RND_CONV_false_4_op_bigger_mux_3_cse;
  wire [5:0] return_add_generic_AC_RND_CONV_false_4_e_dif_sat_or_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_2_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_6_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_7_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_8_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_9_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_10_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_11_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_12_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_13_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_14_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_15_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_16_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_17_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_18_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_19_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_20_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_21_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_22_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_23_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_24_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_25_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_26_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_27_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_28_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_29_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_30_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_31_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_32_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_33_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_34_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_35_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_36_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_37_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_38_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_39_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_40_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_41_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_42_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_43_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_44_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_45_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_46_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_47_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_48_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_49_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_50_cse;
  wire return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_51_cse;
  wire or_450_cse;
  wire stage_PE_1_and_cse;
  wire nor_8_cse;
  wire return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_and_cse;
  wire and_272_cse;
  wire and_277_cse;
  wire and_275_cse;
  wire and_276_cse;
  wire and_271_cse;
  wire return_add_generic_AC_RND_CONV_false_4_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_4_op1_smaller_oelse_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_11_op1_smaller_oelse_and_cse;
  wire return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_and_cse;
  wire return_add_generic_AC_RND_CONV_false_24_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_24_op1_smaller_oelse_and_cse;
  wire return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_and_cse;
  wire return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_and_cse;
  wire and_344_cse;
  wire and_347_cse;
  wire return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_and_1_cse;
  reg t_in_10_0_lpi_1_dfm_1_10;
  reg t_in_10_0_lpi_1_dfm_1_9;
  reg BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm;
  reg [50:0] return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm;
  reg return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm;
  reg [50:0] return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm;
  wire BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx1;
  wire return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx1;
  wire return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50_mx2;
  wire [49:0] return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0_mx2;
  wire return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1;
  reg return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm;
  reg [50:0] return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm;
  wire return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1;
  wire stage_PE_tmp_re_d_1_lpi_3_dfm_51_mx0;
  wire return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_1_op2_mu_51_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_4_op1_mu_52_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_4_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_4_op2_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1;
  reg stage_PE_1_tmp_re_d_1_lpi_3_dfm_51;
  reg stage_PE_1_tmp_im_d_1_lpi_3_dfm_51;
  reg [50:0] stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0;
  wire return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_4_op1_mu_51_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_4_op2_mu_52_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_4_op2_mu_51_1_lpi_3_dfm_mx0;
  reg [8:0] reg_BUTTERFLY_i_div_cmp_a_reg;
  wire BUTTERFLY_1_i_and_ssc;
  reg reg_BUTTERFLY_1_i_9_0_ftd;
  reg [8:0] reg_BUTTERFLY_1_i_9_0_ftd_1;
  wire [15:0] BUTTERFLY_1_else_3_else_acc_4_sdt;
  wire [16:0] nl_BUTTERFLY_1_else_3_else_acc_4_sdt;
  wire BUTTERFLY_1_else_1_if_and_ssc;
  reg [2:0] reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd;
  wire and_1132_ssc;
  wire and_1141_ssc;
  wire and_1143_ssc;
  wire and_1145_ssc;
  wire and_1149_ssc;
  wire return_add_generic_AC_RND_CONV_false_7_exp_and_ssc;
  reg reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd;
  reg [3:0] reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1;
  reg [5:0] reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2;
  reg operator_6_false_18_acc_psp_sva_11;
  wire BUTTERFLY_and_ssc;
  reg [3:0] BUTTERFLY_mux_5_itm_13_10;
  reg [9:0] BUTTERFLY_mux_5_itm_9_0;
  wire stage_PE_1_tmp_im_d_and_ssc;
  reg [12:0] stage_PE_1_tmp_im_d_1_sva_1_63_51;
  reg [50:0] stage_PE_1_tmp_im_d_1_sva_1_50_0;
  wire BUTTERFLY_else_2_and_ssc;
  reg [5:0] BUTTERFLY_else_2_acc_1_psp_16_0_sva_16_11;
  reg [10:0] BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0;
  wire [11:0] operator_6_false_49_acc_sdt;
  wire [12:0] nl_operator_6_false_49_acc_sdt;
  reg [2:0] operator_6_false_49_acc_psp_sva_11_9;
  reg [8:0] operator_6_false_49_acc_psp_sva_8_0;
  reg [4:0] return_add_generic_AC_RND_CONV_false_17_mux_7_itm_55_51;
  reg [50:0] return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0;
  wire nor_99_ssc;
  reg [4:0] return_add_generic_AC_RND_CONV_false_18_mux_1_itm_55_51;
  reg [50:0] return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0;
  reg [1:0] reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_2_1;
  reg reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0;
  wire BUTTERFLY_if_1_or_3_cse;
  wire BUTTERFLY_if_1_or_1_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  wire return_extract_15_m_zero_mux1h_3_cse;
  wire and_1813_cse;
  wire return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_11_mux_19_cse;
  wire return_add_generic_AC_RND_CONV_false_1_mux_16_cse;
  wire return_add_generic_AC_RND_CONV_false_3_mux_10_cse;
  wire return_add_generic_AC_RND_CONV_false_7_if_5_or_cse;
  wire return_add_generic_AC_RND_CONV_false_9_mux_17_cse;
  wire return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm_mx1;
  wire return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_17_op1_smaller_lor_lpi_3_dfm_2;
  wire [11:0] return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0w0;
  wire [12:0] nl_return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0w0;
  wire [11:0] return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0w0;
  wire [12:0] nl_return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0w0;
  wire drf_qr_lval_10_smx_lpi_3_dfm_mx1_10;
  wire [3:0] drf_qr_lval_10_smx_lpi_3_dfm_mx1_9_6;
  wire [5:0] drf_qr_lval_10_smx_lpi_3_dfm_mx1_5_0;
  wire drf_qr_lval_10_smx_lpi_3_dfm_mx2_10;
  wire [3:0] drf_qr_lval_10_smx_lpi_3_dfm_mx2_9_6;
  wire [5:0] drf_qr_lval_10_smx_lpi_3_dfm_mx2_5_0;
  wire [3:0] return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_mx0w4_9_6;
  wire [5:0] return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_mx0w4_5_0;
  wire return_add_generic_AC_RND_CONV_false_3_op_bigger_mux_1_cse;
  wire [50:0] return_add_generic_AC_RND_CONV_false_3_op_bigger_mux_2_cse;
  wire return_add_generic_AC_RND_CONV_false_op_bigger_mux_1_cse;
  wire [50:0] return_add_generic_AC_RND_CONV_false_op_bigger_mux_2_cse;
  wire return_add_generic_AC_RND_CONV_false_16_op_bigger_mux_1_cse;
  wire [50:0] return_add_generic_AC_RND_CONV_false_16_op_bigger_mux_2_cse;
  wire return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_1_cse;
  wire [50:0] return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_cse;
  wire return_add_generic_AC_RND_CONV_false_9_exp_mux1h_2_cse;
  wire return_add_generic_AC_RND_CONV_false_10_op1_mu_mux1h_3_cse;
  wire and_1808_cse;
  wire or_446_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_mux_cse;
  wire return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_cse;
  wire return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_2_cse;
  wire return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_1_cse;
  wire return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_cse;
  wire [49:0] return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse;
  wire return_add_generic_AC_RND_CONV_false_14_op1_mu_mux_1_cse;
  wire or_452_cse;
  wire or_445_cse;
  wire and_1804_cse;
  wire and_1585_rgt;
  wire and_1587_rgt;
  wire or_673_rmff;
  wire or_672_rmff;
  wire or_671_rmff;
  wire or_670_rmff;
  wire or_709_ssc;
  wire or_710_ssc;
  wire or_683_ssc;
  wire or_685_ssc;
  wire [15:0] BUTTERFLY_1_else_1_if_acc_1_sdt;
  wire [16:0] nl_BUTTERFLY_1_else_1_if_acc_1_sdt;
  reg return_add_generic_AC_RND_CONV_false_10_mux_7_itm;
  reg return_add_generic_AC_RND_CONV_false_17_mux_6_itm;
  wire [9:0] return_add_generic_AC_RND_CONV_false_1_e_r_qelse_qr_10_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_1_mux_32;
  wire return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0;
  reg return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs;
  wire return_add_generic_AC_RND_CONV_false_9_mux_35;
  wire return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs_mx0w0;
  reg return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs;
  wire [51:0] return_add_generic_AC_RND_CONV_false_1_res_rounded_lpi_3_dfm_51_0_1;
  wire return_add_generic_AC_RND_CONV_false_13_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_22_or_1_svs_1;
  wire [9:0] BUTTERFLY_i_9_0_sva_1;
  wire [10:0] nl_BUTTERFLY_i_9_0_sva_1;
  reg [9:0] BUTTERFLY_1_fry_9_0_sva;
  wire out_f_d_rsci_adr_d_mx0c2;
  wire out_f_d_rsci_adr_d_mx0c3;
  wire out_f_d_rsci_adr_d_mx0c5;
  wire [9:0] return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_and_9;
  wire [11:0] return_add_generic_AC_RND_CONV_false_10_exp_plus_1_12_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs_mx0w0;
  wire [9:0] return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_and_9;
  wire [11:0] return_add_generic_AC_RND_CONV_false_11_exp_plus_1_12_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_3_mux_26;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w0;
  reg return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs;
  wire return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_and_11;
  wire return_add_generic_AC_RND_CONV_false_10_exp_plus_1_0_lpi_3_dfm_1;
  reg return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs;
  wire return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_and_11;
  wire return_add_generic_AC_RND_CONV_false_11_exp_plus_1_0_lpi_3_dfm_1;
  reg return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs;
  wire [51:0] return_add_generic_AC_RND_CONV_false_3_res_rounded_lpi_3_dfm_51_0_1;
  wire return_add_generic_AC_RND_CONV_false_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_9_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_10_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_11_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_12_or_1_svs_1;
  wire in_f_d_rsci_adr_d_mx0c2;
  wire [14:0] stage_monty_mul_acc_2_psp_sva_1;
  wire [15:0] nl_stage_monty_mul_acc_2_psp_sva_1;
  wire or_dcpl_629;
  wire or_tmp;
  wire or_tmp_829;
  wire or_tmp_830;
  wire or_tmp_833;
  wire or_tmp_834;
  wire or_tmp_835;
  wire or_1342_ssc;
  wire or_1344_ssc;
  wire BUTTERFLY_if_1_if_and_3_cse;
  wire BUTTERFLY_if_1_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_4_e_r_qelse_and_cse;
  wire return_add_generic_AC_RND_CONV_false_4_e_r_qelse_and_1_cse;
  wire stage_PE_tmp_im_d_and_cse;
  wire stage_PE_tmp_im_d_and_2_cse;
  wire [9:0] return_add_generic_AC_RND_CONV_false_9_e_r_return_add_generic_AC_RND_CONV_false_9_e_r_or_cse;
  wire [11:0] return_add_generic_AC_RND_CONV_false_9_exp_plus_1_12_1_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_7_exp_plus_1_12_1_lpi_3_dfm_1;
  reg return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs;
  wire return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs_mx0w0;
  wire [11:0] return_add_generic_AC_RND_CONV_false_24_exp_plus_1_12_1_lpi_3_dfm_1;
  wire or_1477_tmp;
  wire or_1478_tmp;
  wire nor_113_m1c;
  wire or_1482_tmp;
  wire or_1483_tmp;
  wire BUTTERFLY_if_1_or_9_tmp;
  wire or_1484_tmp;
  wire or_1485_tmp;
  wire and_2106_cse;
  wire and_2105_cse;
  wire and_2108_cse;
  wire and_2107_cse;
  wire and_2114_cse;
  wire [11:0] return_add_generic_AC_RND_CONV_false_23_exp_plus_1_12_1_lpi_3_dfm_1;
  wire [9:0] stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1;
  wire [9:0] stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w4_10_1;
  wire [11:0] return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_1;
  wire stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_0;
  wire stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w4_0;
  wire and_2120_cse;
  wire and_2123_cse;
  wire and_2126_cse;
  wire and_2127_cse;
  wire and_2129_cse;
  wire and_2130_cse;
  wire [5:0] return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_3_itm;
  wire [5:0] return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_5_itm;
  wire [5:0] return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_9_itm;
  wire or_1143_itm;
  wire [15:0] in_u_mux1h_1_itm;
  wire [16:0] nl_in_u_mux1h_1_itm;
  wire or_1285_itm;
  wire [16:0] stage_u_add_3_mux1h_2_itm;
  wire [17:0] nl_stage_u_add_3_mux1h_2_itm;
  wire [13:0] BUTTERFLY_1_if_mux_itm;
  wire [10:0] return_add_generic_AC_RND_CONV_false_7_op_bigger_mux_6_itm;
  wire [56:0] return_add_generic_AC_RND_CONV_false_7_rshift_itm;
  wire [54:0] return_add_generic_AC_RND_CONV_false_7_lshift_itm;
  wire [5:0] return_add_generic_AC_RND_CONV_false_8_mux_8_itm;
  wire [5:0] return_add_generic_AC_RND_CONV_false_18_mux_4_itm;
  wire [56:0] return_add_generic_AC_RND_CONV_false_20_rshift_itm;
  wire [54:0] return_add_generic_AC_RND_CONV_false_20_lshift_itm;
  wire [56:0] return_add_generic_AC_RND_CONV_false_25_rshift_itm;
  wire [54:0] return_add_generic_AC_RND_CONV_false_23_lshift_itm;
  wire [51:0] return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm;
  wire [54:0] return_add_generic_AC_RND_CONV_false_19_lshift_1_itm;
  wire [51:0] z_out;
  wire [52:0] nl_z_out;
  wire [16:0] z_out_1;
  wire [17:0] nl_z_out_1;
  wire [56:0] z_out_5;
  wire [56:0] z_out_6;
  wire [56:0] z_out_7;
  wire [56:0] z_out_8;
  wire [56:0] z_out_9;
  wire [49:0] z_out_10;
  wire [9:0] z_out_12;
  wire [10:0] nl_z_out_12;
  wire [12:0] z_out_13;
  wire [10:0] z_out_14;
  wire [12:0] z_out_15;
  wire [13:0] nl_z_out_15;
  wire [12:0] z_out_16;
  wire [13:0] nl_z_out_16;
  wire [11:0] z_out_17;
  wire [11:0] z_out_18;
  wire or_tmp_900;
  wire [11:0] z_out_19;
  wire [11:0] z_out_21;
  wire [12:0] nl_z_out_21;
  wire [23:0] z_out_22;
  wire [24:0] nl_z_out_22;
  wire [17:0] z_out_23;
  wire [18:0] nl_z_out_23;
  wire [11:0] z_out_24;
  wire [12:0] nl_z_out_24;
  wire [31:0] z_out_25;
  wire signed [32:0] nl_z_out_25;
  wire [105:0] z_out_26;
  wire or_tmp_920;
  wire [9:0] z_out_27;
  wire [10:0] nl_z_out_27;
  wire [16:0] z_out_28;
  wire [56:0] z_out_29;
  wire [56:0] z_out_30;
  wire [56:0] z_out_31;
  wire [56:0] z_out_32;
  wire [56:0] z_out_33;
  wire [56:0] z_out_34;
  wire [53:0] z_out_35;
  wire [56:0] z_out_36;
  wire [56:0] z_out_37;
  wire [56:0] z_out_38;
  wire [56:0] z_out_39;
  wire [56:0] z_out_40;
  wire [56:0] z_out_41;
  wire [54:0] z_out_42;
  wire [54:0] z_out_43;
  wire all_same_out;
  wire [5:0] rtn_out;
  wire all_same_out_1;
  wire [5:0] rtn_out_1;
  wire [9:0] z_out_44;
  wire [12:0] z_out_45;
  wire [53:0] z_out_46;
  wire [54:0] nl_z_out_46;
  wire [53:0] z_out_47;
  wire [54:0] nl_z_out_47;
  wire [14:0] z_out_48;
  wire [15:0] nl_z_out_48;
  wire or_tmp_1003;
  wire [11:0] z_out_49;
  wire [11:0] z_out_50;
  wire [11:0] z_out_51;
  wire [11:0] z_out_52;
  wire [52:0] z_out_53;
  wire [105:0] z_out_54;
  wire [11:0] z_out_55;
  wire [12:0] nl_z_out_55;
  wire [11:0] z_out_56;
  wire [12:0] nl_z_out_56;
  wire [12:0] z_out_57;
  wire [16:0] z_out_58;
  wire [17:0] nl_z_out_58;
  wire [15:0] z_out_59;
  wire [16:0] nl_z_out_59;
  wire [17:0] z_out_60;
  wire [18:0] nl_z_out_60;
  wire [17:0] z_out_61;
  wire or_tmp_1041;
  wire [12:0] z_out_63;
  reg return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm;
  reg stage_PE_1_index_const_15_lpi_2_dfm;
  reg stage_PE_1_index_const_10_lpi_2_dfm;
  reg stage_PE_1_index_const_0_lpi_2_dfm;
  reg stage_PE_1_qr_0_lpi_2_dfm;
  reg stage_PE_1_qr_1_0_lpi_2_dfm;
  reg [61:0] stage_PE_1_gm_im_d_61_0_lpi_3_dfm;
  reg return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs;
  reg [56:0] return_add_generic_AC_RND_CONV_false_15_res_mant_4_sva;
  reg return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs;
  reg return_extract_41_return_extract_41_or_1_cse_sva;
  reg return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_22_unequal_tmp;
  reg return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs;
  reg [31:0] BUTTERFLY_1_else_2_tmp2_1_sva;
  reg return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm;
  reg [50:0] return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm;
  reg return_add_generic_AC_RND_CONV_false_18_mux_itm;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_8;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_7;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_8;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_8;
  reg stage_PE_1_tmp_re_d_1_lpi_3_dfm_63;
  wire out1_rsci_idat_63_0_mx0c1;
  wire out1_rsci_idat_63_0_mx0c2;
  wire out1_rsci_idat_79_64_mx0c1;
  wire return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1;
  wire return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs_mx0w0;
  wire mode_lpi_1_dfm_mx0w0;
  wire stage_PE_asn_13_mx0w0;
  wire stage_PE_index_const_15_lpi_2_dfm_mx0w0;
  wire stage_PE_index_const_10_lpi_2_dfm_mx0w0;
  wire BUTTERFLY_1_i_9_0_sva_mx0c3;
  wire return_add_generic_AC_RND_CONV_false_10_if_2_return_add_generic_AC_RND_CONV_false_10_if_2_and_1_mx3w0;
  wire return_extract_17_m_zero_sva_mx0w3;
  wire return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_svs_1;
  wire return_add_generic_AC_RND_CONV_false_3_do_sub_sva_1;
  wire return_extract_41_return_extract_41_or_1_cse_sva_1;
  wire return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_1_op1_smaller_lor_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_1_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_3_res_mant_3_0_sva_1;
  wire BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c0;
  wire BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c4;
  wire BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c7;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_12_if_2_return_add_generic_AC_RND_CONV_false_12_if_2_nor_mx3w0;
  wire return_add_generic_AC_RND_CONV_false_11_if_2_return_add_generic_AC_RND_CONV_false_11_if_2_nor_mx3w0;
  wire return_add_generic_AC_RND_CONV_false_7_if_2_return_add_generic_AC_RND_CONV_false_7_if_2_and_1_mx1w0;
  wire return_add_generic_AC_RND_CONV_false_8_if_2_return_add_generic_AC_RND_CONV_false_8_if_2_and_1_mx2w0;
  wire return_add_generic_AC_RND_CONV_false_2_do_sub_sva_1;
  wire return_add_generic_AC_RND_CONV_false_16_do_sub_sva_1;
  wire return_add_generic_AC_RND_CONV_false_15_do_sub_sva_1;
  wire [56:0] return_add_generic_AC_RND_CONV_false_6_res_mant_4_sva_1;
  wire [58:0] nl_return_add_generic_AC_RND_CONV_false_6_res_mant_4_sva_1;
  wire [56:0] return_add_generic_AC_RND_CONV_false_8_res_mant_4_sva_1;
  wire [58:0] nl_return_add_generic_AC_RND_CONV_false_8_res_mant_4_sva_1;
  wire [56:0] return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_2;
  wire [58:0] nl_return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_2;
  wire [56:0] return_add_generic_AC_RND_CONV_false_21_res_mant_4_sva_1;
  wire [58:0] nl_return_add_generic_AC_RND_CONV_false_21_res_mant_4_sva_1;
  wire drf_qr_lval_10_smx_lpi_3_dfm_mx0c0;
  wire return_extract_13_return_extract_13_or_1_cse_sva_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_1_exp_plus_1_12_1_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_3_exp_plus_1_12_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_3_exp_plus_1_0_lpi_3_dfm_1;
  wire [56:0] return_add_generic_AC_RND_CONV_false_3_res_rounded_asn_rndc_sva_1;
  wire return_add_generic_AC_RND_CONV_false_1_exp_plus_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_5_res_mant_3_0_sva_1;
  wire in_u_rsc_merge_sva_mx0c2;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_mx0w1;
  wire return_extract_45_return_extract_45_or_1_cse_sva_1;
  wire return_add_generic_AC_RND_CONV_false_6_exp_plus_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_17_e_r_qelse_or_svs_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_6_exp_plus_1_12_1_lpi_3_dfm_1;
  wire return_extract_17_return_extract_17_or_sva_1;
  wire return_add_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_2_res_mant_3_0_sva_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_5_e_r_qelse_qr_10_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1;
  wire [51:0] return_add_generic_AC_RND_CONV_false_5_res_rounded_lpi_3_dfm_51_0_1;
  wire return_add_generic_AC_RND_CONV_false_5_e_r_qelse_or_svs_1;
  wire [51:0] return_add_generic_AC_RND_CONV_false_4_res_rounded_lpi_3_dfm_51_0_1;
  wire return_add_generic_AC_RND_CONV_false_4_e_r_qelse_or_svs_1;
  wire [50:0] stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0w0;
  wire [11:0] return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_1_e_incr_lpi_3_dfm_2;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_tmp_1;
  wire [50:0] stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx0w2;
  wire [51:0] return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_1;
  wire return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_50_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0;
  wire return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_19_op1_smaller_lor_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_6_res_mant_3_0_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_3_e_incr_lpi_3_dfm_2;
  wire [51:0] r_rnd_dummy_1_51_0_sva_1;
  wire [52:0] nl_r_rnd_dummy_1_51_0_sva_1;
  wire [52:0] return_mult_generic_AC_RND_CONV_false_res_bef_rnd_3_53_1_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_if_1_and_1_tmp_1;
  wire [11:0] operator_6_false_13_acc_psp_sva_1;
  wire [12:0] nl_operator_6_false_13_acc_psp_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_19_e_dif_sat_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_2_if_1_and_1_tmp_1;
  wire return_extract_19_return_extract_19_or_sva_1;
  wire return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1;
  wire [51:0] return_add_generic_AC_RND_CONV_false_6_res_rounded_lpi_3_dfm_51_0_1;
  wire [56:0] return_add_generic_AC_RND_CONV_false_6_res_rounded_asn_rndc_sva_1;
  wire return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_7_op1_smaller_lor_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_7_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_8_res_mant_3_0_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1;
  wire [51:0] return_add_generic_AC_RND_CONV_false_7_res_rounded_lpi_3_dfm_51_0_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_8_exp_plus_1_12_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_9_res_mant_3_0_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_9_e_dif_sat_sva_1;
  wire return_add_generic_AC_RND_CONV_false_8_exp_plus_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_7_exp_plus_1_0_lpi_3_dfm_1;
  wire [56:0] return_add_generic_AC_RND_CONV_false_7_res_rounded_asn_rndc_sva_1;
  wire return_add_generic_AC_RND_CONV_false_10_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_9_exp_plus_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_14_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_16_res_mant_3_0_sva_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_18_res_mant_3_0_sva_1;
  wire [51:0] return_add_generic_AC_RND_CONV_false_17_res_rounded_lpi_3_dfm_51_0_1;
  wire [11:0] operator_33_true_36_acc_psp_1_sva_1;
  wire [12:0] nl_operator_33_true_36_acc_psp_1_sva_1;
  wire [10:0] operator_6_false_40_acc_psp_1_sva_1;
  wire [11:0] nl_operator_6_false_40_acc_psp_1_sva_1;
  wire [56:0] return_add_generic_AC_RND_CONV_false_17_res_rounded_asn_rndc_sva_1;
  wire [15:0] operator_32_false_1_mul_atp_sva_1;
  wire [16:0] nl_operator_32_false_1_mul_atp_sva_1;
  wire return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_13_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_15_res_mant_3_0_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_4_e_incr_lpi_3_dfm_2;
  wire [51:0] r_rnd_dummy_4_51_0_sva_1;
  wire [52:0] nl_r_rnd_dummy_4_51_0_sva_1;
  wire [52:0] return_mult_generic_AC_RND_CONV_false_4_res_bef_rnd_3_53_1_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_4_if_1_and_1_tmp_1;
  wire return_extract_49_return_extract_49_or_sva_1;
  wire [17:0] stage_u_add_9_acc_psp_sva_1;
  wire [18:0] nl_stage_u_add_9_acc_psp_sva_1;
  wire return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_50_mx0;
  wire return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_19_res_mant_3_0_sva_1;
  wire [52:0] return_mult_generic_AC_RND_CONV_false_3_res_bef_rnd_3_53_1_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_3_if_1_and_1_tmp_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_5_e_incr_lpi_3_dfm_2;
  wire return_mult_generic_AC_RND_CONV_false_5_if_1_and_1_tmp_1;
  wire return_extract_51_return_extract_51_or_sva_1;
  wire return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_19_exp_plus_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_20_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_21_op1_smaller_lor_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_21_res_mant_3_0_sva_1;
  wire [51:0] return_add_generic_AC_RND_CONV_false_20_res_rounded_lpi_3_dfm_51_0_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_21_exp_plus_1_12_1_lpi_3_dfm_1;
  wire [51:0] return_add_generic_AC_RND_CONV_false_21_res_rounded_lpi_3_dfm_51_0_1;
  wire return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_22_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_23_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_24_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_25_res_mant_3_0_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_25_e_dif_sat_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_24_e_dif_sat_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_23_e_dif_sat_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_22_e_dif_sat_sva_1;
  wire return_add_generic_AC_RND_CONV_false_21_exp_plus_1_0_lpi_3_dfm_1;
  wire [56:0] return_add_generic_AC_RND_CONV_false_20_res_rounded_asn_rndc_sva_1;
  wire [51:0] return_add_generic_AC_RND_CONV_false_23_res_rounded_lpi_3_dfm_51_0_1;
  wire [51:0] return_add_generic_AC_RND_CONV_false_24_res_rounded_lpi_3_dfm_51_0_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_25_exp_plus_1_12_1_lpi_3_dfm_1;
  wire [51:0] return_add_generic_AC_RND_CONV_false_25_res_rounded_lpi_3_dfm_51_0_1;
  wire return_add_generic_AC_RND_CONV_false_25_exp_plus_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_24_exp_plus_1_0_lpi_3_dfm_1;
  wire [11:0] operator_6_false_55_acc_psp_sva_1;
  wire [12:0] nl_operator_6_false_55_acc_psp_sva_1;
  wire return_add_generic_AC_RND_CONV_false_23_exp_plus_1_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1;
  wire [52:0] return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_6_if_1_and_1_tmp_1;
  wire [9:0] operator_32_false_2_mul_atp_sva_1;
  wire [10:0] nl_operator_32_false_2_mul_atp_sva_1;
  wire [11:0] operator_33_true_15_acc_2;
  wire [12:0] nl_operator_33_true_15_acc_2;
  wire return_add_generic_AC_RND_CONV_false_6_r_sign_mux_2;
  wire return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_nor_2;
  wire return_add_generic_AC_RND_CONV_false_7_if_5_return_add_generic_AC_RND_CONV_false_7_if_5_nor_2;
  wire return_mult_generic_AC_RND_CONV_false_mux_15;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_else_2_else_else_mux_2;
  wire return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_and_8;
  wire [9:0] stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w0_10_1;
  wire stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w0_0;
  wire return_mult_generic_AC_RND_CONV_false_1_shift_right_conc_3_5;
  wire return_mult_generic_AC_RND_CONV_false_1_shift_right_conc_3_0;
  wire [9:0] stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w2_10_1;
  wire stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w2_0;
  wire return_mult_generic_AC_RND_CONV_false_2_shift_right_conc_3_5;
  wire [3:0] return_mult_generic_AC_RND_CONV_false_2_shift_right_conc_3_4_1;
  wire return_mult_generic_AC_RND_CONV_false_2_shift_right_conc_3_0;
  wire return_mult_generic_AC_RND_CONV_false_5_shift_right_conc_3_5;
  wire [3:0] return_mult_generic_AC_RND_CONV_false_5_shift_right_conc_3_4_1;
  wire return_mult_generic_AC_RND_CONV_false_5_shift_right_conc_3_0;
  wire [5:0] operator_6_false_6_operator_6_false_6_conc_2_6_1;
  wire [6:0] nl_operator_6_false_6_operator_6_false_6_conc_2_6_1;
  wire [5:0] operator_6_false_2_operator_6_false_2_conc_2_6_1;
  wire [6:0] nl_operator_6_false_2_operator_6_false_2_conc_2_6_1;
  wire return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_50;
  wire [49:0] return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0;
  wire return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_and_10_9;
  wire [8:0] return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_and_10_8_0;
  wire [5:0] leading_sign_53_0_1_out_1;
  wire leading_sign_57_0_1_0_15_out_2;
  wire [5:0] leading_sign_57_0_1_0_15_out_3;
  wire leading_sign_57_0_1_0_2_out_2;
  wire [5:0] leading_sign_57_0_1_0_2_out_3;
  wire leading_sign_57_0_1_0_4_out_2;
  wire [5:0] leading_sign_57_0_1_0_4_out_3;
  wire [5:0] leading_sign_53_0_out_1;
  wire leading_sign_57_0_1_0_6_out_2;
  wire [5:0] leading_sign_57_0_1_0_6_out_3;
  wire [5:0] leading_sign_53_0_2_out_1;
  wire leading_sign_57_0_1_0_8_out_2;
  wire [5:0] leading_sign_57_0_1_0_8_out_3;
  wire leading_sign_57_0_1_0_10_out_2;
  wire [5:0] leading_sign_57_0_1_0_10_out_3;
  wire leading_sign_57_0_1_0_18_out_2;
  wire [5:0] leading_sign_57_0_1_0_18_out_3;
  wire leading_sign_57_0_1_0_17_out_2;
  wire [5:0] leading_sign_57_0_1_0_17_out_3;
  wire [5:0] leading_sign_53_0_4_out_1;
  wire leading_sign_57_0_1_0_19_out_2;
  wire [5:0] leading_sign_57_0_1_0_19_out_3;
  wire [5:0] leading_sign_53_0_5_out_1;
  wire leading_sign_57_0_1_0_21_out_2;
  wire [5:0] leading_sign_57_0_1_0_21_out_3;
  wire leading_sign_57_0_1_0_20_out_2;
  wire [5:0] leading_sign_57_0_1_0_20_out_3;
  wire leading_sign_57_0_1_0_25_out_2;
  wire [5:0] leading_sign_57_0_1_0_25_out_3;
  wire leading_sign_57_0_1_0_24_out_2;
  wire [5:0] leading_sign_57_0_1_0_24_out_3;
  wire [5:0] leading_sign_53_0_6_out_1;
  wire [55:0] return_add_generic_AC_RND_CONV_false_4_res_mant_conc_2_itm_56_1;
  wire [5:0] operator_6_false_8_operator_6_false_8_conc_itm_6_1;
  wire [6:0] nl_operator_6_false_8_operator_6_false_8_conc_itm_6_1;
  wire [4:0] return_add_generic_AC_RND_CONV_false_24_mux_4_itm_5_1;
  reg return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_0;
  reg return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_1;
  reg [3:0] return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2;
  reg [3:0] return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_0;
  reg [1:0] return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_1;
  reg [50:0] return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_2;
  reg [5:0] in_u_rsc_merge_sva_rsp_0;
  wire in_u_and_ssc;
  reg operator_6_false_18_acc_psp_sva_10_0_rsp_0;
  wire operator_6_false_18_and_1_ssc;
  reg [3:0] stage_u_add_3_acc_itm_rsp_0;
  reg [12:0] stage_u_add_3_acc_itm_rsp_1;
  wire stage_u_add_3_and_ssc;
  wire drf_qr_lval_6_smx_lpi_3_dfm_mx0_10;
  wire [9:0] drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_0;
  wire [3:0] return_add_generic_AC_RND_CONV_false_21_mux_8_itm_3_0;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_0;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_14_and_cse;
  wire return_add_generic_AC_RND_CONV_false_17_m_r_and_cse;
  wire return_extract_15_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_14_op1_mu_and_cse;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif_qelse_return_add_generic_AC_RND_CONV_false_1_e_dif_qelse_and_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_return_add_generic_AC_RND_CONV_false_11_sticky_bit_return_add_generic_AC_RND_CONV_false_11_sticky_bit_or_cse;
  wire [11:0] return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_18_res_rounded_and_cse;
  wire return_mult_generic_AC_RND_CONV_false_4_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_4_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_4_else_1_sticky_bit_or_cse;
  wire return_add_generic_AC_RND_CONV_false_15_res_mant_or_1_cse;
  wire BUTTERFLY_1_i_or_3_cse;
  wire or_1367_cse;
  wire or_1556_cse;
  wire or_1531_cse;
  wire stage_PE_tmp_im_d_or_cse;
  wire return_mult_generic_AC_RND_CONV_false_2_else_1_nor_cse;
  wire return_add_generic_AC_RND_CONV_false_5_res_rounded_or_1_cse;
  wire return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_2_cse;
  wire [5:0] return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse;
  wire [5:0] return_add_generic_AC_RND_CONV_false_1_e_dif_sat_or_cse;
  wire [5:0] return_add_generic_AC_RND_CONV_false_2_e_dif_sat_or_cse;
  wire [5:0] return_add_generic_AC_RND_CONV_false_e_dif_sat_or_cse;
  wire return_mult_generic_AC_RND_CONV_false_if_or_3_cse;
  wire [3:0] return_mult_generic_AC_RND_CONV_false_if_nand_1_cse;
  wire return_mult_generic_AC_RND_CONV_false_if_or_cse;
  wire return_mult_generic_AC_RND_CONV_false_4_exp_ovf_oif_aelse_nor_cse;
  wire return_add_generic_AC_RND_CONV_false_10_mux_20_cse;
  wire return_add_generic_AC_RND_CONV_false_15_res_mant_or_cse;
  wire operator_6_false_18_or_cse;
  wire for_or_4_cse;
  wire return_add_generic_AC_RND_CONV_false_1_res_rounded_and_1_cse;
  wire for_or_5_cse;
  wire BUTTERFLY_else_2_mux_1_cse;
  wire BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_1_cse;
  wire [2:0] BUTTERFLY_else_1_if_mux_4_cse;
  wire [1:0] BUTTERFLY_else_1_if_mux_5_cse;
  wire BUTTERFLY_else_1_if_mux_6_cse;
  wire return_add_generic_AC_RND_CONV_false_10_mux_17_cse;
  wire or_1266_cse;
  wire return_add_generic_AC_RND_CONV_false_3_and_20_cse;
  wire return_mult_generic_AC_RND_CONV_false_1_else_1_or_cse;
  wire for_or_10_cse_1;
  wire or_1495_cse_1;
  wire return_add_generic_AC_RND_CONV_false_3_and_cse;
  wire return_add_generic_AC_RND_CONV_false_3_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_3_and_2_cse;
  wire return_add_generic_AC_RND_CONV_false_3_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_3_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_3_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_3_and_6_cse;
  wire return_add_generic_AC_RND_CONV_false_3_and_7_cse;
  wire return_add_generic_AC_RND_CONV_false_3_and_8_cse;
  wire return_add_generic_AC_RND_CONV_false_3_and_9_cse;
  wire return_add_generic_AC_RND_CONV_false_1_and_8_cse;
  wire return_add_generic_AC_RND_CONV_false_1_and_9_cse;
  wire return_add_generic_AC_RND_CONV_false_1_and_14_cse;
  wire return_add_generic_AC_RND_CONV_false_1_and_15_cse;
  wire return_add_generic_AC_RND_CONV_false_1_and_28_cse;
  wire return_add_generic_AC_RND_CONV_false_1_and_30_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_2_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_11_or_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_12_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_11_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_13_cse;
  wire and_1029_cse;
  wire return_add_generic_AC_RND_CONV_false_3_or_4_cse;
  wire return_add_generic_AC_RND_CONV_false_3_or_5_cse;
  wire return_add_generic_AC_RND_CONV_false_3_and_30_cse;
  wire return_add_generic_AC_RND_CONV_false_3_and_32_cse;
  wire return_add_generic_AC_RND_CONV_false_5_or_4_cse;
  wire return_add_generic_AC_RND_CONV_false_5_and_6_cse;
  wire return_add_generic_AC_RND_CONV_false_5_and_8_cse;
  wire return_add_generic_AC_RND_CONV_false_5_and_10_cse;
  wire return_add_generic_AC_RND_CONV_false_5_and_7_cse;
  wire return_add_generic_AC_RND_CONV_false_5_and_9_cse;
  wire and_1014_cse;
  wire and_1032_cse;
  wire return_add_generic_AC_RND_CONV_false_3_or_14_cse;
  wire return_add_generic_AC_RND_CONV_false_3_or_16_cse;
  wire return_add_generic_AC_RND_CONV_false_5_or_6_cse;
  wire or_956_cse;
  wire operator_11_true_return_26_sva_2;
  wire mode_or_cse;
  wire return_add_generic_AC_RND_CONV_false_20_ls_or_cse;
  wire return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse;
  wire return_add_generic_AC_RND_CONV_false_10_res_mant_or_9_cse;
  reg t_in_10_0_lpi_1_dfm_1_8;
  wire [9:0] operator_6_false_18_mux1h_itm_10_1;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_6;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_7;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_7;
  reg reg_BUTTERFLY_i_div_cmp_b_ftd;
  reg reg_BUTTERFLY_i_div_cmp_b_ftd_2;
  reg reg_BUTTERFLY_i_div_cmp_b_ftd_3;
  reg reg_BUTTERFLY_i_div_cmp_b_ftd_4;
  reg reg_BUTTERFLY_i_div_cmp_b_ftd_5;
  reg reg_BUTTERFLY_i_div_cmp_b_ftd_7;
  wire and_255_tmp;
  wire and_258_tmp;
  wire and_261_tmp;
  wire and_264_tmp;
  wire return_add_generic_AC_RND_CONV_false_10_and_3_m1c;
  wire return_add_generic_AC_RND_CONV_false_10_and_5_m1c;
  wire return_add_generic_AC_RND_CONV_false_10_and_7_m1c;
  wire return_add_generic_AC_RND_CONV_false_10_and_9_m1c;
  wire return_add_generic_AC_RND_CONV_false_10_and_11_m1c;
  wire return_add_generic_AC_RND_CONV_false_10_and_13_m1c;
  wire return_add_generic_AC_RND_CONV_false_11_and_26_m1c;
  wire return_add_generic_AC_RND_CONV_false_11_and_28_m1c;
  wire return_add_generic_AC_RND_CONV_false_11_and_32_m1c;
  wire return_add_generic_AC_RND_CONV_false_11_and_34_m1c;
  wire return_add_generic_AC_RND_CONV_false_12_and_6_m1c;
  wire and_342_tmp;
  wire and_352_tmp;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_1;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_0;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_1;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_1;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_0;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_1;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_0;
  wire BUTTERFLY_i_or_4_ssc;
  wire BUTTERFLY_i_or_5_ssc;
  reg reg_BUTTERFLY_i_div_cmp_b_ftd_6_1;
  reg reg_BUTTERFLY_i_div_cmp_b_ftd_6_0;
  wire BUTTERFLY_else_1_if_or_3_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_5_cse;
  wire return_extract_41_and_1_cse;
  wire stage_u_add_3_or_1_cse;
  wire or_954_rgt;
  wire or_955_rgt;
  wire or_959_rgt;
  wire or_960_rgt;
  wire BUTTERFLY_else_2_and_2_rgt;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_2;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_2;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_2;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_2;
  reg reg_BUTTERFLY_i_div_cmp_b_ftd_6_2;
  wire BUTTERFLY_i_or_3_cse;
  wire return_add_generic_AC_RND_CONV_false_14_op1_mu_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_14_op1_mu_and_2_cse;
  wire return_add_generic_AC_RND_CONV_false_17_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_14_op1_mu_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_14_op1_mu_and_6_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse;
  wire return_add_generic_AC_RND_CONV_false_10_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_27_cse;
  wire return_add_generic_AC_RND_CONV_false_10_and_6_cse;
  wire return_add_generic_AC_RND_CONV_false_10_and_12_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_18_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_11_cse;
  wire return_add_generic_AC_RND_CONV_false_18_and_8_cse;
  wire and_1134_cse;
  wire BUTTERFLY_1_fiy_and_4_cse;
  wire BUTTERFLY_1_fiy_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_14_op1_mu_and_13_cse;
  wire return_add_generic_AC_RND_CONV_false_17_and_7_cse;
  wire return_add_generic_AC_RND_CONV_false_17_and_8_cse;
  wire return_add_generic_AC_RND_CONV_false_17_and_9_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_18_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_5_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_24_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse;
  wire return_add_generic_AC_RND_CONV_false_11_exp_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_11_exp_and_2_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_13_cse;
  wire return_add_generic_AC_RND_CONV_false_14_op1_mu_and_8_cse;
  wire return_add_generic_AC_RND_CONV_false_14_op1_mu_and_7_cse;
  wire return_add_generic_AC_RND_CONV_false_14_op1_mu_and_12_cse;
  wire return_add_generic_AC_RND_CONV_false_14_op1_mu_and_11_cse;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_3;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_3;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_3;
  reg reg_BUTTERFLY_i_div_cmp_b_ftd_6_3;
  wire return_add_generic_AC_RND_CONV_false_10_and_16_cse;
  wire return_add_generic_AC_RND_CONV_false_10_and_17_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_37_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_38_cse;
  wire return_add_generic_AC_RND_CONV_false_10_and_18_cse;
  wire return_add_generic_AC_RND_CONV_false_10_and_19_cse;
  wire return_add_generic_AC_RND_CONV_false_10_and_24_cse;
  wire return_add_generic_AC_RND_CONV_false_10_and_25_cse;
  wire stage_PE_1_tmp_im_d_and_6_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_cse;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_4;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_5;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_4;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_4;
  reg reg_BUTTERFLY_i_div_cmp_b_ftd_6_5;
  reg reg_BUTTERFLY_i_div_cmp_b_ftd_6_4;
  reg t_in_10_0_lpi_1_dfm_1_7;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_5;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_6;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_5;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_6;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_5;
  reg t_in_10_0_lpi_1_dfm_1_6;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_6;
  reg t_in_10_0_lpi_1_dfm_1_5;
  reg t_in_10_0_lpi_1_dfm_1_4;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_7;
  reg t_in_10_0_lpi_1_dfm_1_3;
  reg t_in_10_0_lpi_1_dfm_1_2;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_8;
  reg t_in_10_0_lpi_1_dfm_1_1;
  reg t_in_10_0_lpi_1_dfm_1_0;
  reg m_in_15_1_lpi_1_dfm_1_rsp_0_9;
  wire stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_0;
  reg m_in_15_1_lpi_1_dfm_1_rsp_0_10;
  reg stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_1;
  reg reg_BUTTERFLY_i_div_cmp_b_1_ftd_1;
  wire stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_1;
  reg m_in_15_1_lpi_1_dfm_1_rsp_0_11;
  reg stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_1;
  reg reg_BUTTERFLY_i_div_cmp_b_1_ftd_3;
  wire stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_3;
  wire stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_2;
  reg m_in_15_1_lpi_1_dfm_1_rsp_0_13;
  reg m_in_15_1_lpi_1_dfm_1_rsp_0_12;
  reg stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_0_rsp_0;
  reg stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_0_rsp_1;
  reg reg_BUTTERFLY_i_div_cmp_b_1_ftd;
  reg reg_BUTTERFLY_i_div_cmp_b_1_ftd_4;
  wire nor_88_cse;
  wire nor_87_cse;
  wire nor_90_cse;
  wire nor_145_cse;
  wire BUTTERFLY_1_else_1_if_nor_cse;
  wire and_2638_cse;
  wire [49:0] return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1;
  wire return_add_generic_AC_RND_CONV_false_11_and_45_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_46_cse;
  wire nor_155_cse;
  wire return_add_generic_AC_RND_CONV_false_14_or_cse;
  wire stage_PE_qif_qelse_mux_15_itm;
  wire [9:0] and_2143_itm;
  wire or_965_itm;
  wire return_add_generic_AC_RND_CONV_false_1_and_itm;
  wire return_add_generic_AC_RND_CONV_false_1_and_1_itm;
  wire return_add_generic_AC_RND_CONV_false_1_and_2_itm;
  wire return_add_generic_AC_RND_CONV_false_1_and_3_itm;
  wire return_add_generic_AC_RND_CONV_false_5_or_1_itm;
  wire return_add_generic_AC_RND_CONV_false_10_ma1_lt_ma2_acc_1_itm_52;
  wire return_mult_generic_AC_RND_CONV_false_2_if_acc_1_itm_12_1;
  wire return_mult_generic_AC_RND_CONV_false_1_if_acc_1_itm_12_1;
  wire return_mult_generic_AC_RND_CONV_false_5_if_acc_1_itm_12_1;
  wire return_mult_generic_AC_RND_CONV_false_4_if_acc_1_itm_12_1;
  wire return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_19_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_5_acc_2_itm_10_1;
  wire return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1;
  wire return_add_generic_AC_RND_CONV_false_18_acc_2_itm_10;
  wire return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10;
  wire return_add_generic_AC_RND_CONV_false_21_ma1_lt_ma2_acc_1_itm_52;
  wire return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11;
  wire return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11;
  wire return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_2_acc_3_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_22_acc_3_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1;
  wire return_mult_generic_AC_RND_CONV_false_3_if_acc_2_itm_12_1;
  wire return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1;
  wire [4:0] return_add_generic_AC_RND_CONV_false_9_conc_59_itm_5_1;
  reg [8:0] reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0;
  reg reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1;
  wire and_2620_ssc;
  reg [3:0] in_u_rsc_merge_sva_rsp_1_rsp_0;
  reg [5:0] in_u_rsc_merge_sva_rsp_1_rsp_1;
  reg [8:0] operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0;
  reg operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1;
  wire [8:0] return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1_9_1;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1_0;
  wire [8:0] return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1_9_1;
  wire return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1_0;
  wire [3:0] return_add_generic_AC_RND_CONV_false_10_e_dif_sat_conc_4_itm_4_1;
  wire [3:0] return_add_generic_AC_RND_CONV_false_10_exp_conc_5_itm_10_7;
  wire [5:0] return_add_generic_AC_RND_CONV_false_10_exp_conc_5_itm_6_1;
  wire [3:0] return_add_generic_AC_RND_CONV_false_23_mux_11_itm_5_2;
  wire [8:0] return_add_generic_AC_RND_CONV_false_12_e_dif_qr_lpi_3_dfm_mx0_9_1;
  wire [8:0] return_add_generic_AC_RND_CONV_false_11_e_dif_qr_lpi_3_dfm_mx0_9_1;
  wire [8:0] BUTTERFLY_else_1_if_mux_7_cse_9_1;
  wire BUTTERFLY_else_1_if_mux_7_cse_0;
  wire return_add_generic_AC_RND_CONV_false_11_e_dif_sat_or_1_seb;
  wire [4:0] return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1_5_1;
  wire return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1_0;
  wire return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_1_seb;
  wire [4:0] return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1_5_1;
  wire return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1_0;
  wire BUTTERFLY_else_1_if_and_cse;
  wire BUTTERFLY_else_1_if_and_1_cse;
  wire BUTTERFLY_else_1_if_and_5_cse;
  wire BUTTERFLY_1_nor_1_cse;
  wire return_mult_generic_AC_RND_CONV_false_1_else_1_and_1_cse;
  wire return_mult_generic_AC_RND_CONV_false_1_else_1_return_mult_generic_AC_RND_CONV_false_1_else_1_mux_2_cse;
  wire return_add_generic_AC_RND_CONV_false_1_and_54_cse;
  wire return_add_generic_AC_RND_CONV_false_1_and_55_cse;
  wire z_out_2_52;
  wire z_out_3_52;
  wire z_out_20_11;
  wire [15:0] z_out_64_31_16;
  wire return_add_generic_AC_RND_CONV_false_21_res_rounded_and_cse;
  wire return_mult_generic_AC_RND_CONV_false_1_mux1h_8_m1c;
  wire return_mult_generic_AC_RND_CONV_false_1_mux1h_9_m1c;
  wire return_mult_generic_AC_RND_CONV_false_1_mux1h_10_m1c;
  wire return_add_generic_AC_RND_CONV_false_20_op_bigger_mux_7_tmp;

  wire[10:0] return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_or_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_6_else_2_else_return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_6_else_2_else_mux_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_acc_nl;
  wire[11:0] nl_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_acc_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl;
  wire BUTTERFLY_if_1_and_nl;
  wire BUTTERFLY_if_1_and_1_nl;
  wire[50:0] return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_oelse_3_not_1_nl;
  wire stage_PE_index_const_mux_nl;
  wire stage_PE_index_const_mux_3_nl;
  wire stage_PE_index_const_mux_2_nl;
  wire stage_PE_index_const_mux_7_nl;
  wire stage_PE_mux1h_nl;
  wire stage_PE_mux1h_7_nl;
  wire stage_PE_mux1h_1_nl;
  wire stage_PE_mux1h_9_nl;
  wire stage_PE_mux1h_2_nl;
  wire stage_PE_mux1h_11_nl;
  wire BUTTERFLY_i_and_14_nl;
  wire BUTTERFLY_i_or_7_nl;
  wire stage_PE_mux1h_3_nl;
  wire stage_PE_mux1h_13_nl;
  wire[8:0] BUTTERFLY_i_mux_1_nl;
  wire t_in_not_nl;
  wire BUTTERFLY_if_mux_12_nl;
  wire stage_PE_stage_PE_stage_PE_mux_3_nl;
  wire BUTTERFLY_if_mux_13_nl;
  wire BUTTERFLY_if_mux_14_nl;
  wire BUTTERFLY_if_mux_15_nl;
  wire BUTTERFLY_if_mux_16_nl;
  wire BUTTERFLY_if_mux_17_nl;
  wire BUTTERFLY_if_mux_18_nl;
  wire BUTTERFLY_if_mux_19_nl;
  wire BUTTERFLY_if_mux_20_nl;
  wire BUTTERFLY_if_mux_21_nl;
  wire t_in_mux_4_nl;
  wire not_681_nl;
  wire stage_PE_qif_qelse_mux_18_nl;
  wire stage_PE_qif_qelse_mux_5_nl;
  wire stage_PE_qif_qelse_or_nl;
  wire stage_PE_qif_qelse_mux_19_nl;
  wire[9:0] BUTTERFLY_fry_BUTTERFLY_fry_mux_nl;
  wire[8:0] BUTTERFLY_n_and_nl;
  wire[8:0] BUTTERFLY_n_BUTTERFLY_n_mux_nl;
  wire nand_97_nl;
  wire BUTTERFLY_i_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_3_nl;
  wire return_add_generic_AC_RND_CONV_false_25_r_nan_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_14_op1_mu_and_3_nl;
  wire return_add_generic_AC_RND_CONV_false_14_op1_mu_and_4_nl;
  wire return_add_generic_AC_RND_CONV_false_1_if_2_return_add_generic_AC_RND_CONV_false_1_if_2_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_9_if_2_return_add_generic_AC_RND_CONV_false_9_if_2_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_16_if_2_return_add_generic_AC_RND_CONV_false_16_if_2_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_13_if_2_return_add_generic_AC_RND_CONV_false_13_if_2_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_10_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_10_or_5_nl;
  wire return_add_generic_AC_RND_CONV_false_10_and_15_nl;
  wire return_add_generic_AC_RND_CONV_false_10_or_nl;
  wire return_add_generic_AC_RND_CONV_false_10_or_6_nl;
  wire return_add_generic_AC_RND_CONV_false_10_or_7_nl;
  wire return_add_generic_AC_RND_CONV_false_10_and_8_nl;
  wire return_add_generic_AC_RND_CONV_false_10_and_21_nl;
  wire return_add_generic_AC_RND_CONV_false_10_and_10_nl;
  wire return_add_generic_AC_RND_CONV_false_10_and_22_nl;
  wire return_add_generic_AC_RND_CONV_false_10_and_23_nl;
  wire return_extract_17_m_zero_return_extract_17_m_zero_nor_nl;
  wire return_extract_47_m_zero_return_extract_47_m_zero_nor_nl;
  wire return_extract_59_m_zero_return_extract_59_m_zero_nor_nl;
  wire or_916_nl;
  wire return_extract_45_m_zero_return_extract_45_m_zero_nor_nl;
  wire return_extract_44_m_zero_return_extract_44_m_zero_nor_nl;
  wire return_extract_52_m_zero_return_extract_52_m_zero_nor_nl;
  wire return_extract_57_m_zero_return_extract_57_m_zero_nor_nl;
  wire return_extract_17_m_zero_or_1_nl;
  wire operator_11_true_12_operator_11_true_12_and_nl;
  wire operator_11_true_20_operator_11_true_20_and_nl;
  wire operator_11_true_25_operator_11_true_25_and_nl;
  wire operator_11_true_45_operator_11_true_45_and_nl;
  wire operator_11_true_44_operator_11_true_44_and_nl;
  wire operator_11_true_52_operator_11_true_52_and_nl;
  wire operator_11_true_57_operator_11_true_57_and_nl;
  wire or_934_nl;
  wire BUTTERFLY_and_5_nl;
  wire BUTTERFLY_and_6_nl;
  wire return_add_generic_AC_RND_CONV_false_17_or_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_24_return_add_generic_AC_RND_CONV_false_24_and_4_nl;
  wire return_add_generic_AC_RND_CONV_false_24_if_7_return_add_generic_AC_RND_CONV_false_24_if_7_nor_nl;
  wire or_939_nl;
  wire or_940_nl;
  wire and_990_nl;
  wire and_992_nl;
  wire return_add_generic_AC_RND_CONV_false_17_or_4_nl;
  wire return_add_generic_AC_RND_CONV_false_17_or_5_nl;
  wire[9:0] mux1h_3_nl;
  wire[9:0] operator_33_true_37_acc_nl;
  wire[10:0] nl_operator_33_true_37_acc_nl;
  wire and_1161_nl;
  wire and_1163_nl;
  wire and_1169_nl;
  wire and_1171_nl;
  wire not_734_nl;
  wire return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_3_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_nl;
  wire return_add_generic_AC_RND_CONV_false_10_do_sub_return_add_generic_AC_RND_CONV_false_10_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_19_do_sub_return_add_generic_AC_RND_CONV_false_19_do_sub_return_add_generic_AC_RND_CONV_false_19_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_xnor_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_acc_1_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_acc_1_nl;
  wire return_add_generic_AC_RND_CONV_false_4_if_2_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_4_if_2_return_add_generic_AC_RND_CONV_false_4_if_2_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_4_r_sign_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_12_if_2_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_25_r_sign_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_5_if_2_return_add_generic_AC_RND_CONV_false_5_if_2_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_5_r_sign_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_3_if_2_return_add_generic_AC_RND_CONV_false_3_if_2_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_2_if_2_return_add_generic_AC_RND_CONV_false_2_if_2_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_14_if_2_return_add_generic_AC_RND_CONV_false_14_if_2_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_25_nl;
  wire return_add_generic_AC_RND_CONV_false_11_or_4_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_36_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_31_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_42_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_33_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_44_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_10_ma1_lt_ma2_acc_1_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_10_ma1_lt_ma2_acc_1_nl;
  wire return_add_generic_AC_RND_CONV_false_if_2_return_add_generic_AC_RND_CONV_false_if_2_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_7_do_sub_return_add_generic_AC_RND_CONV_false_7_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_15_if_2_return_add_generic_AC_RND_CONV_false_15_if_2_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_20_do_sub_return_add_generic_AC_RND_CONV_false_20_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_5_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_13_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_14_nl;
  wire return_extract_50_and_nl;
  wire return_extract_15_m_zero_return_extract_15_m_zero_nor_nl;
  wire return_extract_27_m_zero_return_extract_27_m_zero_nor_nl;
  wire return_extract_17_m_zero_or_2_nl;
  wire operator_11_true_13_operator_11_true_13_and_nl;
  wire operator_11_true_53_operator_11_true_53_and_nl;
  wire operator_11_true_27_operator_11_true_27_and_nl;
  wire operator_11_true_59_operator_11_true_59_and_nl;
  wire return_add_generic_AC_RND_CONV_false_6_do_sub_return_add_generic_AC_RND_CONV_false_6_do_sub_return_add_generic_AC_RND_CONV_false_6_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_21_do_sub_return_add_generic_AC_RND_CONV_false_21_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_8_do_sub_return_add_generic_AC_RND_CONV_false_8_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_22_do_sub_return_add_generic_AC_RND_CONV_false_22_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_5_e_dif_sat_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_10_e_dif_sat_or_1_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_14_mux1h_8_nl;
  wire nor_157_nl;
  wire[57:0] acc_4_nl;
  wire[58:0] nl_acc_4_nl;
  wire[55:0] return_add_generic_AC_RND_CONV_false_3_mux1h_17_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_18_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_19_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_20_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_21_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_3_mux1h_22_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_23_nl;
  wire return_add_generic_AC_RND_CONV_false_3_or_17_nl;
  wire return_add_generic_AC_RND_CONV_false_15_res_mant_or_4_nl;
  wire return_add_generic_AC_RND_CONV_false_15_res_mant_or_5_nl;
  wire stage_PE_1_x_im_d_and_1_nl;
  wire[3:0] and_2119_nl;
  wire[3:0] mux1h_nl;
  wire not_730_nl;
  wire[5:0] and_2131_nl;
  wire[5:0] mux1h_2_nl;
  wire not_732_nl;
  wire mux_22_nl;
  wire and_2628_nl;
  wire mux_21_nl;
  wire mux_20_nl;
  wire or_1755_nl;
  wire BUTTERFLY_else_2_and_8_nl;
  wire return_add_generic_AC_RND_CONV_false_18_return_add_generic_AC_RND_CONV_false_18_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_18_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_18_and_3_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_25_return_add_generic_AC_RND_CONV_false_25_and_4_nl;
  wire return_add_generic_AC_RND_CONV_false_25_if_7_return_add_generic_AC_RND_CONV_false_25_if_7_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_18_and_15_nl;
  wire and_304_nl;
  wire return_extract_54_m_zero_return_extract_54_m_zero_nor_nl;
  wire[3:0] operator_32_false_acc_nl;
  wire[4:0] nl_operator_32_false_acc_nl;
  wire return_add_generic_AC_RND_CONV_false_19_op2_mu_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_19_op2_mu_and_3_nl;
  wire or_1195_nl;
  wire BUTTERFLY_1_fiy_and_1_nl;
  wire BUTTERFLY_1_fiy_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_1_r_nan_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_14_r_nan_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_23_r_nan_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_9_exp_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_9_exp_or_nl;
  wire return_add_generic_AC_RND_CONV_false_9_exp_and_5_nl;
  wire return_add_generic_AC_RND_CONV_false_9_exp_and_7_nl;
  wire return_add_generic_AC_RND_CONV_false_9_exp_and_9_nl;
  wire return_add_generic_AC_RND_CONV_false_9_exp_and_10_nl;
  wire[9:0] mux_25_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_14_e_r_and_5_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_14_e_r_mux1h_6_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_25_e_r_qelse_return_add_generic_AC_RND_CONV_false_25_e_r_qelse_and_nl;
  wire return_add_generic_AC_RND_CONV_false_25_e_r_qelse_not_2_nl;
  wire return_add_generic_AC_RND_CONV_false_14_e_r_nor_2_nl;
  wire or_1771_nl;
  wire or_1772_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_r_return_add_generic_AC_RND_CONV_false_1_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_5_nl;
  wire return_add_generic_AC_RND_CONV_false_25_e_r_qelse_return_add_generic_AC_RND_CONV_false_25_e_r_qelse_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_25_mux_13_nl;
  wire return_add_generic_AC_RND_CONV_false_25_return_add_generic_AC_RND_CONV_false_25_and_5_nl;
  wire return_add_generic_AC_RND_CONV_false_25_e_r_qelse_mux_1_nl;
  wire or_312_nl;
  wire stage_PE_1_tmp_im_d_and_5_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_3_return_mult_generic_AC_RND_CONV_false_1_if_3_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_if_3_return_mult_generic_AC_RND_CONV_false_2_if_3_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_if_3_return_mult_generic_AC_RND_CONV_false_5_if_3_or_1_nl;
  wire return_extract_13_m_zero_return_extract_13_m_zero_nor_nl;
  wire return_extract_12_m_zero_return_extract_12_m_zero_nor_nl;
  wire return_extract_20_m_zero_return_extract_20_m_zero_nor_nl;
  wire return_extract_25_m_zero_return_extract_25_m_zero_nor_nl;
  wire[9:0] stage_PE_tmp_im_d_mux1h_nl;
  wire not_726_nl;
  wire operator_11_true_17_operator_11_true_17_and_nl;
  wire operator_11_true_22_operator_11_true_22_and_nl;
  wire operator_11_true_54_operator_11_true_54_and_nl;
  wire return_extract_15_return_extract_15_nor_nl;
  wire return_extract_47_return_extract_47_nor_nl;
  wire operator_11_true_15_operator_11_true_15_and_nl;
  wire operator_11_true_47_operator_11_true_47_and_nl;
  wire return_extract_15_return_extract_15_or_1_nl;
  wire return_extract_47_return_extract_47_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_mux_13_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_1_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_1_else_1_sticky_bit_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_mux_13_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_if_1_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_2_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_2_else_1_sticky_bit_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_mux_13_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_if_1_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_5_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_5_else_1_sticky_bit_or_nl;
  wire return_add_generic_AC_RND_CONV_false_10_op2_mu_and_3_nl;
  wire return_add_generic_AC_RND_CONV_false_10_op2_mu_and_4_nl;
  wire return_add_generic_AC_RND_CONV_false_18_return_add_generic_AC_RND_CONV_false_18_and_5_nl;
  wire return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_24_r_nan_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_11_exp_and_3_nl;
  wire return_add_generic_AC_RND_CONV_false_11_exp_and_4_nl;
  wire return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_and_8_nl;
  wire return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_17_mux_19_nl;
  wire return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nand_nl;
  wire return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_23_e_r_return_add_generic_AC_RND_CONV_false_23_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_23_mux_20_nl;
  wire return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_and_4_nl;
  wire return_add_generic_AC_RND_CONV_false_23_e_r_qelse_mux_1_nl;
  wire or_319_nl;
  wire return_add_generic_AC_RND_CONV_false_24_e_r_return_add_generic_AC_RND_CONV_false_24_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_6_if_5_return_add_generic_AC_RND_CONV_false_6_if_5_and_nl;
  wire return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_18_mux_13_nl;
  wire return_add_generic_AC_RND_CONV_false_18_e_r_qelse_nand_nl;
  wire return_add_generic_AC_RND_CONV_false_18_e_r_qelse_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_24_e_r_qelse_return_add_generic_AC_RND_CONV_false_24_e_r_qelse_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_24_mux_13_nl;
  wire return_add_generic_AC_RND_CONV_false_24_return_add_generic_AC_RND_CONV_false_24_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_24_e_r_qelse_mux_1_nl;
  wire or_306_nl;
  wire return_add_generic_AC_RND_CONV_false_25_e_r_return_add_generic_AC_RND_CONV_false_25_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_19_op2_mu_return_add_generic_AC_RND_CONV_false_19_op2_mu_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_19_op2_mu_and_5_nl;
  wire return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_nl;
  wire return_add_generic_AC_RND_CONV_false_9_do_sub_return_add_generic_AC_RND_CONV_false_9_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_23_do_sub_return_add_generic_AC_RND_CONV_false_23_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_2_nl;
  wire[12:0] return_mult_generic_AC_RND_CONV_false_2_if_acc_1_nl;
  wire[13:0] nl_return_mult_generic_AC_RND_CONV_false_2_if_acc_1_nl;
  wire[12:0] return_mult_generic_AC_RND_CONV_false_1_if_acc_1_nl;
  wire[13:0] nl_return_mult_generic_AC_RND_CONV_false_1_if_acc_1_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux_29_nl;
  wire return_add_generic_AC_RND_CONV_false_1_if_5_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux_23_nl;
  wire return_add_generic_AC_RND_CONV_false_3_if_5_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_6_mux_32_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_8_mux_13_nl;
  wire[12:0] return_mult_generic_AC_RND_CONV_false_5_if_acc_1_nl;
  wire[13:0] nl_return_mult_generic_AC_RND_CONV_false_5_if_acc_1_nl;
  wire[12:0] return_mult_generic_AC_RND_CONV_false_4_if_acc_1_nl;
  wire[13:0] nl_return_mult_generic_AC_RND_CONV_false_4_if_acc_1_nl;
  wire return_add_generic_AC_RND_CONV_false_20_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_21_mux_13_nl;
  wire[11:0] return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl;
  wire[12:0] nl_return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl;
  wire return_add_generic_AC_RND_CONV_false_9_mux_32_nl;
  wire return_add_generic_AC_RND_CONV_false_9_if_5_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_10_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_11_mux_9_nl;
  wire return_add_generic_AC_RND_CONV_false_24_mux_9_nl;
  wire return_add_generic_AC_RND_CONV_false_24_if_5_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_25_mux_9_nl;
  wire return_add_generic_AC_RND_CONV_false_25_if_5_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_23_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_23_if_5_or_1_nl;
  wire stage_PE_qif_qelse_mux_11_nl;
  wire return_add_generic_AC_RND_CONV_false_18_mux_9_nl;
  wire return_add_generic_AC_RND_CONV_false_18_if_5_or_1_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_1_else_2_else_return_mult_generic_AC_RND_CONV_false_1_else_2_else_and_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_1_else_2_else_else_mux_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_3_else_2_else_return_mult_generic_AC_RND_CONV_false_3_else_2_else_and_nl;
  wire return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif_sat_or_1_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_18_ma1_lt_ma2_acc_2_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_18_ma1_lt_ma2_acc_2_nl;
  wire and_287_nl;
  wire and_292_nl;
  wire return_add_generic_AC_RND_CONV_false_7_r_sign_mux_1_nl;
  wire nand_84_nl;
  wire return_add_generic_AC_RND_CONV_false_20_r_sign_mux_1_nl;
  wire nand_85_nl;
  wire return_add_generic_AC_RND_CONV_false_5_if_7_not_7_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_oelse_3_return_mult_generic_AC_RND_CONV_false_3_if_3_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_4_if_7_not_6_nl;
  wire return_add_generic_AC_RND_CONV_false_8_if_7_return_add_generic_AC_RND_CONV_false_8_if_7_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_5_if_7_not_5_nl;
  wire return_add_generic_AC_RND_CONV_false_21_if_7_return_add_generic_AC_RND_CONV_false_21_if_7_nor_nl;
  wire[55:0] return_add_generic_AC_RND_CONV_false_5_mux_20_nl;
  wire return_add_generic_AC_RND_CONV_false_5_mux_19_nl;
  wire[55:0] return_add_generic_AC_RND_CONV_false_6_mux_31_nl;
  wire return_add_generic_AC_RND_CONV_false_6_mux_30_nl;
  wire return_add_generic_AC_RND_CONV_false_6_op_bigger_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_6_op_bigger_mux_2_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_6_op_bigger_mux_9_nl;
  wire return_add_generic_AC_RND_CONV_false_6_op_bigger_mux_3_nl;
  wire[55:0] return_add_generic_AC_RND_CONV_false_8_mux_25_nl;
  wire return_add_generic_AC_RND_CONV_false_8_mux_24_nl;
  wire return_add_generic_AC_RND_CONV_false_8_op_bigger_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_8_op_bigger_mux_2_nl;
  wire return_add_generic_AC_RND_CONV_false_8_op_bigger_mux_4_nl;
  wire return_add_generic_AC_RND_CONV_false_5_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_10_mux_26_nl;
  wire return_add_generic_AC_RND_CONV_false_10_op_bigger_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_10_op_bigger_mux_1_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_10_op_bigger_mux_2_nl;
  wire return_add_generic_AC_RND_CONV_false_10_op_bigger_mux_3_nl;
  wire[55:0] return_add_generic_AC_RND_CONV_false_21_mux_23_nl;
  wire return_add_generic_AC_RND_CONV_false_21_mux_22_nl;
  wire return_add_generic_AC_RND_CONV_false_21_op_bigger_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_21_op_bigger_mux_2_nl;
  wire return_add_generic_AC_RND_CONV_false_21_op_bigger_mux_4_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_else_2_else_return_mult_generic_AC_RND_CONV_false_else_2_else_and_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_4_else_2_else_return_mult_generic_AC_RND_CONV_false_4_else_2_else_and_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_4_else_2_else_else_mux_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_8_ma1_lt_ma2_acc_1_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_8_ma1_lt_ma2_acc_1_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_20_ma1_lt_ma2_acc_1_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_20_ma1_lt_ma2_acc_1_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl;
  wire return_add_generic_AC_RND_CONV_false_3_r_nan_or_1_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_3_return_add_generic_AC_RND_CONV_false_3_and_4_nl;
  wire return_add_generic_AC_RND_CONV_false_3_if_7_return_add_generic_AC_RND_CONV_false_3_if_7_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_1_nl;
  wire[9:0] mux_16_nl;
  wire and_2152_nl;
  wire not_736_nl;
  wire return_add_generic_AC_RND_CONV_false_1_not_6_nl;
  wire[9:0] mux_17_nl;
  wire and_2154_nl;
  wire not_738_nl;
  wire[11:0] operator_33_true_7_acc_1_nl;
  wire[12:0] nl_operator_33_true_7_acc_1_nl;
  wire return_add_generic_AC_RND_CONV_false_3_res_rounded_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_3_not_6_nl;
  wire return_add_generic_AC_RND_CONV_false_3_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_1_if_5_or_nl;
  wire and_328_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_7_e_r_qelse_return_add_generic_AC_RND_CONV_false_7_e_r_qelse_and_nl;
  wire return_add_generic_AC_RND_CONV_false_7_e_r_qelse_not_2_nl;
  wire return_add_generic_AC_RND_CONV_false_21_e_r_qelse_return_add_generic_AC_RND_CONV_false_21_e_r_qelse_and_nl;
  wire return_add_generic_AC_RND_CONV_false_21_mux_16_nl;
  wire[8:0] return_add_generic_AC_RND_CONV_false_21_e_r_qelse_return_add_generic_AC_RND_CONV_false_21_e_r_qelse_and_2_nl;
  wire[8:0] return_add_generic_AC_RND_CONV_false_21_mux_24_nl;
  wire return_add_generic_AC_RND_CONV_false_21_e_r_qelse_not_3_nl;
  wire return_add_generic_AC_RND_CONV_false_8_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_8_e_r_qelse_mux_1_nl;
  wire or_230_nl;
  wire return_add_generic_AC_RND_CONV_false_21_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_21_e_r_qelse_mux_1_nl;
  wire or_249_nl;
  wire return_add_generic_AC_RND_CONV_false_6_mux_6_nl;
  wire return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_and_nl;
  wire return_add_generic_AC_RND_CONV_false_19_mux_6_nl;
  wire return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_and_nl;
  wire return_add_generic_AC_RND_CONV_false_16_r_nan_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_5_nl;
  wire return_add_generic_AC_RND_CONV_false_25_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_25_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_17_mux_15_nl;
  wire return_add_generic_AC_RND_CONV_false_17_if_5_or_1_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_6_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_6_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_11_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_11_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_19_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_19_acc_2_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_16_return_add_generic_AC_RND_CONV_false_16_and_4_nl;
  wire return_add_generic_AC_RND_CONV_false_16_if_7_return_add_generic_AC_RND_CONV_false_16_if_7_nor_nl;
  wire[11:0] operator_33_true_13_acc_nl;
  wire[12:0] nl_operator_33_true_13_acc_nl;
  wire[11:0] return_mult_generic_AC_RND_CONV_false_1_exp_acc_1_nl;
  wire[12:0] nl_return_mult_generic_AC_RND_CONV_false_1_exp_acc_1_nl;
  wire return_add_generic_AC_RND_CONV_false_5_if_7_not_6_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_4_mux_18_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_1_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux_19_nl;
  wire return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_2_nl;
  wire return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_8_r_sign_mux_1_nl;
  wire nand_87_nl;
  wire return_add_generic_AC_RND_CONV_false_21_r_sign_mux_1_nl;
  wire nand_88_nl;
  wire return_add_generic_AC_RND_CONV_false_2_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif_sat_or_1_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_5_mux_12_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_1_nl;
  wire[9:0] operator_33_true_11_acc_nl;
  wire[10:0] nl_operator_33_true_11_acc_nl;
  wire return_add_generic_AC_RND_CONV_false_5_mux_13_nl;
  wire return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_2_nl;
  wire return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_5_not_3_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_5_acc_2_nl;
  wire[11:0] nl_return_add_generic_AC_RND_CONV_false_5_acc_2_nl;
  wire return_add_generic_AC_RND_CONV_false_5_mux_9_nl;
  wire return_add_generic_AC_RND_CONV_false_5_if_5_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_4_not_3_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_4_acc_2_nl;
  wire[11:0] nl_return_add_generic_AC_RND_CONV_false_4_acc_2_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux_15_nl;
  wire return_add_generic_AC_RND_CONV_false_4_if_5_or_1_nl;
  wire return_extract_27_return_extract_27_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_8_r_nan_or_1_nl;
  wire and_357_nl;
  wire return_add_generic_AC_RND_CONV_false_21_r_nan_or_1_nl;
  wire and_359_nl;
  wire return_add_generic_AC_RND_CONV_false_8_e_r_qelse_return_add_generic_AC_RND_CONV_false_8_e_r_qelse_and_nl;
  wire return_add_generic_AC_RND_CONV_false_8_mux_16_nl;
  wire[8:0] return_add_generic_AC_RND_CONV_false_8_e_r_qelse_return_add_generic_AC_RND_CONV_false_8_e_r_qelse_and_2_nl;
  wire[8:0] return_add_generic_AC_RND_CONV_false_8_mux_28_nl;
  wire return_add_generic_AC_RND_CONV_false_8_e_r_qelse_not_3_nl;
  wire return_extract_13_return_extract_13_return_extract_13_m_zero_not_6_nl;
  wire return_extract_13_return_extract_13_return_extract_13_m_zero_not_5_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_21_nl;
  wire return_add_generic_AC_RND_CONV_false_7_e_r_qelse_mux_1_nl;
  wire or_222_nl;
  wire[5:0] operator_6_false_12_acc_nl;
  wire[6:0] nl_operator_6_false_12_acc_nl;
  wire return_add_generic_AC_RND_CONV_false_2_r_nan_or_1_nl;
  wire and_362_nl;
  wire and_365_nl;
  wire return_add_generic_AC_RND_CONV_false_2_if_7_return_add_generic_AC_RND_CONV_false_2_if_7_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_3_nl;
  wire or_206_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_if_not_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_15_r_nan_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_7_nl;
  wire return_add_generic_AC_RND_CONV_false_24_mux_14_nl;
  wire return_add_generic_AC_RND_CONV_false_24_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_15_if_7_return_add_generic_AC_RND_CONV_false_15_if_7_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_18_not_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_oelse_3_return_mult_generic_AC_RND_CONV_false_if_3_nor_nl;
  wire[8:0] return_mult_generic_AC_RND_CONV_false_2_exp_mux_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_exp_mux_2_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_19_ma1_lt_ma2_acc_2_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_19_ma1_lt_ma2_acc_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_if_not_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_return_mult_generic_AC_RND_CONV_false_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_dif_sat_or_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_if_not_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_oelse_3_return_mult_generic_AC_RND_CONV_false_4_if_3_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_6_res_rounded_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_if_if_not_nl;
  wire[11:0] return_mult_generic_AC_RND_CONV_false_2_exp_acc_1_nl;
  wire[12:0] nl_return_mult_generic_AC_RND_CONV_false_2_exp_acc_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_6_r_nan_or_1_nl;
  wire and_369_nl;
  wire return_add_generic_AC_RND_CONV_false_6_if_7_return_add_generic_AC_RND_CONV_false_6_if_7_nor_nl;
  wire[8:0] return_add_generic_AC_RND_CONV_false_6_e_r_qelse_return_add_generic_AC_RND_CONV_false_6_e_r_qelse_and_nl;
  wire[8:0] return_add_generic_AC_RND_CONV_false_6_mux_18_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_not_6_nl;
  wire return_add_generic_AC_RND_CONV_false_6_mux_35_nl;
  wire return_add_generic_AC_RND_CONV_false_6_mux_19_nl;
  wire return_add_generic_AC_RND_CONV_false_19_e_r_qelse_mux_nl;
  wire or_214_nl;
  wire return_add_generic_AC_RND_CONV_false_6_not_4_nl;
  wire return_add_generic_AC_RND_CONV_false_6_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_6_if_5_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_if_not_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_7_e_dif_qif_acc_1_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_7_e_dif_qif_acc_1_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_7_ma1_lt_ma2_acc_1_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_7_ma1_lt_ma2_acc_1_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_8_e_dif_qif_acc_1_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_8_e_dif_qif_acc_1_nl;
  wire return_add_generic_AC_RND_CONV_false_8_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_7_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_7_res_rounded_and_nl;
  wire return_add_generic_AC_RND_CONV_false_7_r_nan_or_1_nl;
  wire and_373_nl;
  wire return_add_generic_AC_RND_CONV_false_7_not_3_nl;
  wire[11:0] operator_33_true_17_acc_nl;
  wire[12:0] nl_operator_33_true_17_acc_nl;
  wire return_add_generic_AC_RND_CONV_false_7_if_7_return_add_generic_AC_RND_CONV_false_7_if_7_nor_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_9_e_dif_qif_acc_1_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_9_e_dif_qif_acc_1_nl;
  wire return_extract_25_return_extract_25_or_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_10_e_dif_qif_acc_1_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_10_e_dif_qif_acc_1_nl;
  wire return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_8_mux_14_nl;
  wire return_add_generic_AC_RND_CONV_false_8_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_18_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_dif_qelse_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_dif_qelse_mux_2_nl;
  wire return_add_generic_AC_RND_CONV_false_9_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_10_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_dif_qelse_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_dif_qelse_mux_2_nl;
  wire return_add_generic_AC_RND_CONV_false_11_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_11_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_17_not_3_nl;
  wire[5:0] operator_6_false_39_acc_nl;
  wire[6:0] nl_operator_6_false_39_acc_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_18_acc_2_nl;
  wire[11:0] nl_return_add_generic_AC_RND_CONV_false_18_acc_2_nl;
  wire[5:0] operator_6_false_37_acc_nl;
  wire[6:0] nl_operator_6_false_37_acc_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_17_acc_2_nl;
  wire[11:0] nl_return_add_generic_AC_RND_CONV_false_17_acc_2_nl;
  wire return_add_generic_AC_RND_CONV_false_17_res_rounded_and_nl;
  wire[3:0] operator_32_false_1_acc_nl;
  wire[4:0] nl_operator_32_false_1_acc_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_mux_13_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_if_1_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_return_mult_generic_AC_RND_CONV_false_4_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_4_if_7_not_7_nl;
  wire return_extract_2_return_extract_2_return_extract_2_m_zero_not_7_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_return_mult_generic_AC_RND_CONV_false_3_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_if_if_not_nl;
  wire[11:0] return_mult_generic_AC_RND_CONV_false_5_exp_acc_1_nl;
  wire[12:0] nl_return_mult_generic_AC_RND_CONV_false_5_exp_acc_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_19_r_nan_or_1_nl;
  wire and_376_nl;
  wire return_add_generic_AC_RND_CONV_false_19_if_7_return_add_generic_AC_RND_CONV_false_19_if_7_nor_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_19_e_r_qelse_return_add_generic_AC_RND_CONV_false_19_e_r_qelse_and_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_19_mux_18_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_not_3_nl;
  wire return_add_generic_AC_RND_CONV_false_19_mux_19_nl;
  wire return_add_generic_AC_RND_CONV_false_19_e_r_qelse_mux_2_nl;
  wire or_241_nl;
  wire return_add_generic_AC_RND_CONV_false_19_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_19_if_5_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_if_not_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_21_ma1_lt_ma2_acc_1_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_21_ma1_lt_ma2_acc_1_nl;
  wire return_add_generic_AC_RND_CONV_false_20_res_rounded_and_nl;
  wire return_add_generic_AC_RND_CONV_false_20_r_nan_or_1_nl;
  wire and_378_nl;
  wire return_add_generic_AC_RND_CONV_false_20_not_3_nl;
  wire[11:0] operator_33_true_43_acc_nl;
  wire[12:0] nl_operator_33_true_43_acc_nl;
  wire return_add_generic_AC_RND_CONV_false_21_not_3_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_20_e_r_qelse_return_add_generic_AC_RND_CONV_false_20_e_r_qelse_and_nl;
  wire return_add_generic_AC_RND_CONV_false_20_e_r_qelse_not_2_nl;
  wire return_add_generic_AC_RND_CONV_false_20_mux_21_nl;
  wire return_add_generic_AC_RND_CONV_false_20_e_r_qelse_mux_1_nl;
  wire or_245_nl;
  wire return_add_generic_AC_RND_CONV_false_20_if_7_return_add_generic_AC_RND_CONV_false_20_if_7_nor_nl;
  wire return_extract_57_return_extract_57_or_2_nl;
  wire return_extract_59_return_extract_59_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_25_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_24_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_23_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_22_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_21_mux_14_nl;
  wire return_add_generic_AC_RND_CONV_false_21_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_20_mux_18_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_23_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_23_acc_2_nl;
  wire[11:0] operator_33_true_47_acc_nl;
  wire[12:0] nl_operator_33_true_47_acc_nl;
  wire return_add_generic_AC_RND_CONV_false_23_res_rounded_and_nl;
  wire return_add_generic_AC_RND_CONV_false_23_not_3_nl;
  wire[5:0] operator_6_false_54_acc_nl;
  wire[6:0] nl_operator_6_false_54_acc_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_24_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_24_acc_2_nl;
  wire[11:0] operator_33_true_49_acc_nl;
  wire[12:0] nl_operator_33_true_49_acc_nl;
  wire return_add_generic_AC_RND_CONV_false_24_not_3_nl;
  wire[5:0] operator_6_false_56_acc_nl;
  wire[6:0] nl_operator_6_false_56_acc_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_25_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_25_acc_2_nl;
  wire[11:0] operator_33_true_51_acc_nl;
  wire[12:0] nl_operator_33_true_51_acc_nl;
  wire return_add_generic_AC_RND_CONV_false_25_res_rounded_and_nl;
  wire return_add_generic_AC_RND_CONV_false_25_not_3_nl;
  wire return_add_generic_AC_RND_CONV_false_23_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_23_if_5_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_if_if_not_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_mux_1_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_15_acc_3_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_15_acc_3_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_2_acc_3_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_2_acc_3_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_22_acc_3_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_22_acc_3_nl;
  wire return_add_generic_AC_RND_CONV_false_3_return_add_generic_AC_RND_CONV_false_3_and_8_nl;
  wire return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_10_nl;
  wire return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_and_10_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_10_acc_3_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_10_acc_3_nl;
  wire[12:0] return_mult_generic_AC_RND_CONV_false_3_if_acc_2_nl;
  wire[13:0] nl_return_mult_generic_AC_RND_CONV_false_3_if_acc_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_1_or_1_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_21_acc_3_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_21_acc_3_nl;
  wire[3:0] for_acc_nl;
  wire[4:0] nl_for_acc_nl;
  wire BUTTERFLY_1_i_mux1h_2_nl;
  wire or_723_nl;
  wire or_726_nl;
  wire[8:0] mux1h_4_nl;
  wire nor_129_nl;
  wire BUTTERFLY_if_1_if_mux1h_nl;
  wire BUTTERFLY_if_1_if_or_nl;
  wire BUTTERFLY_if_1_if_or_1_nl;
  wire[9:0] or_1488_nl;
  wire[9:0] and_2164_nl;
  wire[9:0] mux1h_1_nl;
  wire and_2157_nl;
  wire and_2158_nl;
  wire and_2159_nl;
  wire and_2160_nl;
  wire and_2161_nl;
  wire or_1732_nl;
  wire BUTTERFLY_if_1_if_and_10_nl;
  wire BUTTERFLY_if_1_if_and_11_nl;
  wire not_741_nl;
  wire BUTTERFLY_if_1_if_mux1h_2_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_return_add_generic_AC_RND_CONV_false_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_3_nl;
  wire or_202_nl;
  wire return_add_generic_AC_RND_CONV_false_9_e_r_return_add_generic_AC_RND_CONV_false_9_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_22_e_r_qelse_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_10_e_r_return_add_generic_AC_RND_CONV_false_10_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_10_e_r_qelse_mux_1_nl;
  wire or_281_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_return_add_generic_AC_RND_CONV_false_11_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_11_mux_13_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_1_nl;
  wire or_292_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_r_return_add_generic_AC_RND_CONV_false_12_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_1_nl;
  wire or_300_nl;
  wire BUTTERFLY_if_1_if_or_2_nl;
  wire BUTTERFLY_if_1_if_mux1h_3_nl;
  wire return_add_generic_AC_RND_CONV_false_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_9_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_10_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_11_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_12_r_nan_or_nl;
  wire BUTTERFLY_if_1_if_and_nl;
  wire BUTTERFLY_if_1_if_and_2_nl;
  wire BUTTERFLY_if_1_if_or_3_nl;
  wire[50:0] and_2165_nl;
  wire[50:0] mux1h_5_nl;
  wire and_2166_nl;
  wire and_2167_nl;
  wire and_2168_nl;
  wire and_2169_nl;
  wire and_2170_nl;
  wire or_1733_nl;
  wire not_742_nl;
  wire BUTTERFLY_1_i_mux1h_1_nl;
  wire[8:0] BUTTERFLY_1_i_mux1h_7_nl;
  wire BUTTERFLY_else_1_if_or_nl;
  wire BUTTERFLY_if_1_mux1h_2_nl;
  wire[8:0] mux1h_6_nl;
  wire nor_130_nl;
  wire BUTTERFLY_if_1_mux1h_1_nl;
  wire BUTTERFLY_if_1_or_nl;
  wire[9:0] or_1489_nl;
  wire[9:0] mux1h_7_nl;
  wire and_2176_nl;
  wire or_1491_nl;
  wire and_2179_nl;
  wire BUTTERFLY_if_1_mux1h_7_nl;
  wire return_add_generic_AC_RND_CONV_false_13_e_r_return_add_generic_AC_RND_CONV_false_13_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_7_nl;
  wire return_add_generic_AC_RND_CONV_false_22_e_r_return_add_generic_AC_RND_CONV_false_22_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_22_e_r_qelse_mux_3_nl;
  wire BUTTERFLY_if_1_or_4_nl;
  wire BUTTERFLY_if_1_mux1h_8_nl;
  wire return_add_generic_AC_RND_CONV_false_13_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_22_r_nan_or_nl;
  wire BUTTERFLY_if_1_and_2_nl;
  wire BUTTERFLY_if_1_and_4_nl;
  wire[50:0] and_2181_nl;
  wire[50:0] mux1h_8_nl;
  wire and_2182_nl;
  wire or_1492_nl;
  wire and_2186_nl;
  wire not_746_nl;
  wire BUTTERFLY_1_i_mux1h_nl;
  wire[8:0] BUTTERFLY_1_i_mux1h_8_nl;
  wire[2:0] BUTTERFLY_else_1_if_mux1h_1_nl;
  wire[1:0] BUTTERFLY_else_1_if_mux1h_7_nl;
  wire BUTTERFLY_else_1_if_mux1h_8_nl;
  wire[9:0] BUTTERFLY_else_1_if_mux1h_9_nl;
  wire[9:0] mux_18_nl;
  wire and_2189_nl;
  wire not_748_nl;
  wire[3:0] return_mult_generic_AC_RND_CONV_false_1_if_nand_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_not_nl;
  wire return_add_generic_AC_RND_CONV_false_11_mux_23_nl;
  wire stage_u_add_3_and_1_nl;
  wire stage_u_add_3_and_3_nl;
  wire operator_14_false_1_or_nl;
  wire stage_PE_qif_qelse_mux_12_nl;
  wire stage_PE_qif_qelse_mux_16_nl;
  wire stage_PE_qif_qelse_mux_1_nl;
  wire stage_PE_qif_qelse_mux_17_nl;
  wire mux_19_nl;
  wire and_2619_nl;
  wire mux_nl;
  wire or_1746_nl;
  wire or_1743_nl;
  wire[3:0] or_1486_nl;
  wire[3:0] and_2115_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_4_e_r_qelse_mux1h_nl;
  wire not_724_nl;
  wire[5:0] or_1487_nl;
  wire[5:0] and_2116_nl;
  wire[5:0] return_add_generic_AC_RND_CONV_false_4_e_r_qelse_mux1h_1_nl;
  wire not_725_nl;
  wire and_2118_nl;
  wire stage_PE_tmp_im_d_mux1h_1_nl;
  wire[51:0] return_mult_generic_AC_RND_CONV_false_mux1h_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_mux1h_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_mux_12_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_if_1_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_or_1_nl;
  wire[3:0] operator_32_false_operator_32_false_or_3_nl;
  wire[5:0] operator_32_false_mux_7_nl;
  wire[3:0] operator_32_false_mux_8_nl;
  wire[5:0] operator_32_false_mux_9_nl;
  wire[53:0] acc_2_nl;
  wire[54:0] nl_acc_2_nl;
  wire return_add_generic_AC_RND_CONV_false_9_ma1_lt_ma2_mux_4_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_9_ma1_lt_ma2_mux_5_nl;
  wire[53:0] acc_3_nl;
  wire[54:0] nl_acc_3_nl;
  wire[51:0] return_add_generic_AC_RND_CONV_false_3_ma1_lt_ma2_mux_3_nl;
  wire[57:0] acc_5_nl;
  wire[58:0] nl_acc_5_nl;
  wire[4:0] return_add_generic_AC_RND_CONV_false_17_mux_32_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_17_mux_33_nl;
  wire return_add_generic_AC_RND_CONV_false_17_mux_34_nl;
  wire return_add_generic_AC_RND_CONV_false_17_mux_35_nl;
  wire return_add_generic_AC_RND_CONV_false_17_mux_36_nl;
  wire return_add_generic_AC_RND_CONV_false_17_mux_37_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_17_mux_38_nl;
  wire return_add_generic_AC_RND_CONV_false_17_mux_39_nl;
  wire[57:0] acc_6_nl;
  wire[58:0] nl_acc_6_nl;
  wire[4:0] return_add_generic_AC_RND_CONV_false_18_mux_23_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_18_mux_24_nl;
  wire return_add_generic_AC_RND_CONV_false_18_mux_25_nl;
  wire return_add_generic_AC_RND_CONV_false_18_mux_26_nl;
  wire return_add_generic_AC_RND_CONV_false_18_mux_27_nl;
  wire return_add_generic_AC_RND_CONV_false_18_mux_28_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_18_mux_29_nl;
  wire return_add_generic_AC_RND_CONV_false_18_mux_30_nl;
  wire[57:0] acc_7_nl;
  wire[58:0] nl_acc_7_nl;
  wire[55:0] return_add_generic_AC_RND_CONV_false_1_mux1h_20_nl;
  wire return_add_generic_AC_RND_CONV_false_1_or_13_nl;
  wire return_add_generic_AC_RND_CONV_false_1_or_14_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_21_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_22_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_23_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_24_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_1_mux1h_25_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_26_nl;
  wire return_add_generic_AC_RND_CONV_false_1_or_15_nl;
  wire return_add_generic_AC_RND_CONV_false_1_or_16_nl;
  wire[57:0] acc_8_nl;
  wire[58:0] nl_acc_8_nl;
  wire[55:0] return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_mux1h_1_nl;
  wire return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_7_and_4_nl;
  wire return_add_generic_AC_RND_CONV_false_7_and_5_nl;
  wire return_add_generic_AC_RND_CONV_false_7_and_6_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_40_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_41_nl;
  wire return_add_generic_AC_RND_CONV_false_12_mux_23_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_42_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_43_nl;
  wire return_add_generic_AC_RND_CONV_false_7_op_bigger_mux_13_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_44_nl;
  wire return_add_generic_AC_RND_CONV_false_7_op_bigger_mux_14_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_7_mux_45_nl;
  wire return_add_generic_AC_RND_CONV_false_7_and_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_46_nl;
  wire return_add_generic_AC_RND_CONV_false_7_op_bigger_mux_15_nl;
  wire[57:0] acc_9_nl;
  wire[58:0] nl_acc_9_nl;
  wire[55:0] return_add_generic_AC_RND_CONV_false_11_mux1h_17_nl;
  wire return_add_generic_AC_RND_CONV_false_11_or_7_nl;
  wire return_add_generic_AC_RND_CONV_false_11_or_8_nl;
  wire return_add_generic_AC_RND_CONV_false_11_mux1h_18_nl;
  wire return_add_generic_AC_RND_CONV_false_11_mux1h_19_nl;
  wire return_add_generic_AC_RND_CONV_false_11_mux1h_20_nl;
  wire return_add_generic_AC_RND_CONV_false_11_mux1h_21_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_11_mux1h_22_nl;
  wire return_add_generic_AC_RND_CONV_false_11_or_9_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_48_nl;
  wire return_add_generic_AC_RND_CONV_false_11_mux1h_23_nl;
  wire[13:0] acc_11_nl;
  wire[14:0] nl_acc_11_nl;
  wire for_and_4_nl;
  wire for_mux1h_11_nl;
  wire[2:0] for_and_5_nl;
  wire[2:0] for_mux1h_12_nl;
  wire not_889_nl;
  wire[4:0] for_and_6_nl;
  wire[4:0] for_mux1h_13_nl;
  wire not_890_nl;
  wire for_and_7_nl;
  wire for_mux1h_14_nl;
  wire for_or_14_nl;
  wire for_mux1h_15_nl;
  wire for_or_15_nl;
  wire for_for_or_1_nl;
  wire for_mux_1_nl;
  wire for_mux1h_16_nl;
  wire for_mux1h_17_nl;
  wire for_mux1h_18_nl;
  wire[1:0] for_mux1h_19_nl;
  wire for_mux1h_20_nl;
  wire[11:0] acc_12_nl;
  wire[12:0] nl_acc_12_nl;
  wire operator_6_false_9_mux_6_nl;
  wire operator_6_false_9_mux_7_nl;
  wire[3:0] operator_6_false_9_mux_8_nl;
  wire operator_6_false_19_mux_5_nl;
  wire[3:0] operator_6_false_19_mux_6_nl;
  wire[5:0] operator_6_false_19_mux_7_nl;
  wire[5:0] operator_6_false_19_mux_8_nl;
  wire[5:0] operator_6_false_19_acc_1_nl;
  wire[6:0] nl_operator_6_false_19_acc_1_nl;
  wire[5:0] operator_6_false_48_acc_1_nl;
  wire[6:0] nl_operator_6_false_48_acc_1_nl;
  wire operator_6_false_19_mux_9_nl;
  wire operator_6_false_17_mux1h_7_nl;
  wire[2:0] operator_6_false_17_mux1h_8_nl;
  wire operator_6_false_17_mux1h_9_nl;
  wire[4:0] operator_6_false_17_mux1h_10_nl;
  wire operator_6_false_17_mux1h_11_nl;
  wire[5:0] operator_6_false_17_mux1h_12_nl;
  wire[5:0] operator_6_false_17_acc_1_nl;
  wire[6:0] nl_operator_6_false_17_acc_1_nl;
  wire[5:0] operator_6_false_23_acc_1_nl;
  wire[6:0] nl_operator_6_false_23_acc_1_nl;
  wire[5:0] operator_6_false_27_acc_1_nl;
  wire[6:0] nl_operator_6_false_27_acc_1_nl;
  wire[5:0] operator_6_false_46_acc_1_nl;
  wire[6:0] nl_operator_6_false_46_acc_1_nl;
  wire[5:0] operator_6_false_41_acc_1_nl;
  wire[6:0] nl_operator_6_false_41_acc_1_nl;
  wire operator_6_false_17_mux1h_13_nl;
  wire[12:0] acc_15_nl;
  wire[13:0] nl_acc_15_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_1_e_dif_qif_return_add_generic_AC_RND_CONV_false_1_e_dif_qif_mux_2_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_1_e_dif_qif_return_add_generic_AC_RND_CONV_false_1_e_dif_qif_mux_3_nl;
  wire[12:0] acc_16_nl;
  wire[13:0] nl_acc_16_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_1_e_dif1_return_add_generic_AC_RND_CONV_false_1_e_dif1_mux_2_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_1_e_dif1_return_add_generic_AC_RND_CONV_false_1_e_dif1_mux_3_nl;
  wire[12:0] acc_17_nl;
  wire[13:0] nl_acc_17_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_8_nl;
  wire[8:0] return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_9_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_11_nl;
  wire[8:0] return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_12_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_13_nl;
  wire[12:0] acc_18_nl;
  wire[13:0] nl_acc_18_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_4_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_5_nl;
  wire[5:0] operator_32_false_operator_32_false_and_2_nl;
  wire operator_32_false_nor_2_nl;
  wire[1:0] operator_32_false_operator_32_false_and_3_nl;
  wire[1:0] operator_32_false_mux_10_nl;
  wire operator_32_false_nor_3_nl;
  wire[1:0] operator_32_false_mux1h_11_nl;
  wire operator_32_false_and_5_nl;
  wire operator_32_false_mux1h_12_nl;
  wire operator_32_false_and_6_nl;
  wire operator_32_false_mux1h_13_nl;
  wire operator_32_false_and_7_nl;
  wire operator_32_false_mux1h_14_nl;
  wire operator_32_false_and_8_nl;
  wire operator_32_false_mux1h_15_nl;
  wire[1:0] operator_32_false_mux1h_16_nl;
  wire[5:0] operator_32_false_mux1h_17_nl;
  wire operator_32_false_and_9_nl;
  wire operator_32_false_mux1h_18_nl;
  wire operator_32_false_or_3_nl;
  wire operator_32_false_mux1h_19_nl;
  wire[6:0] operator_32_false_operator_32_false_or_4_nl;
  wire operator_32_false_or_4_nl;
  wire[3:0] operator_32_false_mux1h_20_nl;
  wire[11:0] operator_32_false_operator_32_false_or_5_nl;
  wire[11:0] operator_32_false_mux_11_nl;
  wire[11:0] return_mult_generic_AC_RND_CONV_false_2_exp_plus_1_mux_1_nl;
  wire[3:0] BUTTERFLY_1_else_2_mux_5_nl;
  wire[9:0] BUTTERFLY_1_else_2_mux_6_nl;
  wire[1:0] BUTTERFLY_1_else_1_BUTTERFLY_1_else_1_and_1_nl;
  wire[5:0] BUTTERFLY_1_else_1_mux_9_nl;
  wire[3:0] BUTTERFLY_1_else_1_mux_10_nl;
  wire[5:0] BUTTERFLY_1_else_1_mux_11_nl;
  wire BUTTERFLY_i_and_16_nl;
  wire BUTTERFLY_i_and_17_nl;
  wire BUTTERFLY_i_BUTTERFLY_i_mux_3_nl;
  wire[41:0] BUTTERFLY_i_BUTTERFLY_i_and_1_nl;
  wire[41:0] BUTTERFLY_i_mux_12_nl;
  wire not_898_nl;
  wire[8:0] BUTTERFLY_i_mux1h_22_nl;
  wire BUTTERFLY_i_or_8_nl;
  wire BUTTERFLY_i_and_18_nl;
  wire BUTTERFLY_i_mux1h_23_nl;
  wire BUTTERFLY_i_and_19_nl;
  wire BUTTERFLY_i_BUTTERFLY_i_mux_4_nl;
  wire BUTTERFLY_i_and_20_nl;
  wire BUTTERFLY_i_mux1h_24_nl;
  wire[39:0] BUTTERFLY_i_and_21_nl;
  wire[39:0] BUTTERFLY_i_mux1h_25_nl;
  wire not_902_nl;
  wire BUTTERFLY_i_mux1h_26_nl;
  wire BUTTERFLY_i_mux1h_27_nl;
  wire BUTTERFLY_i_mux1h_28_nl;
  wire BUTTERFLY_i_mux1h_29_nl;
  wire BUTTERFLY_i_mux1h_30_nl;
  wire BUTTERFLY_i_mux1h_31_nl;
  wire BUTTERFLY_i_mux1h_32_nl;
  wire BUTTERFLY_i_mux1h_33_nl;
  wire BUTTERFLY_i_mux1h_34_nl;
  wire BUTTERFLY_i_mux1h_35_nl;
  wire BUTTERFLY_fry_mux_10_nl;
  wire BUTTERFLY_fry_mux_11_nl;
  wire BUTTERFLY_fry_mux_12_nl;
  wire BUTTERFLY_fry_mux_13_nl;
  wire BUTTERFLY_fry_mux_14_nl;
  wire BUTTERFLY_fry_mux_15_nl;
  wire BUTTERFLY_fry_mux_16_nl;
  wire BUTTERFLY_fry_mux_17_nl;
  wire BUTTERFLY_fry_mux_18_nl;
  wire BUTTERFLY_fry_mux_19_nl;
  wire[17:0] acc_24_nl;
  wire[18:0] nl_acc_24_nl;
  wire[13:0] acc_25_nl;
  wire[14:0] nl_acc_25_nl;
  wire[11:0] return_mult_generic_AC_RND_CONV_false_3_exp_mux_5_nl;
  wire[11:0] return_mult_generic_AC_RND_CONV_false_exp_acc_4_nl;
  wire[12:0] nl_return_mult_generic_AC_RND_CONV_false_exp_acc_4_nl;
  wire[11:0] return_mult_generic_AC_RND_CONV_false_4_exp_acc_2_nl;
  wire[12:0] nl_return_mult_generic_AC_RND_CONV_false_4_exp_acc_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_exp_mux_6_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_exp_mux_7_nl;
  wire[8:0] return_mult_generic_AC_RND_CONV_false_3_exp_mux_8_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_exp_mux_9_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_5_res_rounded_return_add_generic_AC_RND_CONV_false_5_res_rounded_mux_2_nl;
  wire return_add_generic_AC_RND_CONV_false_5_res_rounded_return_add_generic_AC_RND_CONV_false_5_res_rounded_mux_3_nl;
  wire return_add_generic_AC_RND_CONV_false_5_res_rounded_and_1_nl;
  wire[13:0] operator_6_false_25_mux_5_nl;
  wire operator_6_false_25_operator_6_false_25_or_1_nl;
  wire[2:0] operator_6_false_25_operator_6_false_25_and_1_nl;
  wire[8:0] operator_6_false_25_mux_6_nl;
  wire operator_6_false_25_mux_7_nl;
  wire operator_6_false_25_mux_8_nl;
  wire[12:0] acc_29_nl;
  wire[13:0] nl_acc_29_nl;
  wire BUTTERFLY_1_BUTTERFLY_1_and_3_nl;
  wire BUTTERFLY_1_BUTTERFLY_1_and_4_nl;
  wire BUTTERFLY_1_mux_1548_nl;
  wire[2:0] BUTTERFLY_1_mux1h_7_nl;
  wire[5:0] BUTTERFLY_1_mux1h_8_nl;
  wire BUTTERFLY_1_or_1_nl;
  wire BUTTERFLY_1_BUTTERFLY_1_or_2_nl;
  wire[4:0] BUTTERFLY_1_BUTTERFLY_1_and_5_nl;
  wire[4:0] BUTTERFLY_1_mux_1549_nl;
  wire not_905_nl;
  wire BUTTERFLY_1_BUTTERFLY_1_or_3_nl;
  wire BUTTERFLY_1_mux_1550_nl;
  wire[12:0] acc_30_nl;
  wire[13:0] nl_acc_30_nl;
  wire operator_6_false_18_mux1h_22_nl;
  wire[3:0] operator_6_false_18_mux1h_23_nl;
  wire[5:0] operator_6_false_18_mux1h_24_nl;
  wire[5:0] operator_6_false_18_mux1h_25_nl;
  wire[12:0] acc_31_nl;
  wire[13:0] nl_acc_31_nl;
  wire[3:0] operator_6_false_3_mux1h_6_nl;
  wire[5:0] operator_6_false_3_mux1h_7_nl;
  wire operator_6_false_3_mux1h_8_nl;
  wire[4:0] operator_6_false_3_mux1h_9_nl;
  wire operator_6_false_3_mux1h_10_nl;
  wire[12:0] acc_32_nl;
  wire[13:0] nl_acc_32_nl;
  wire[3:0] operator_6_false_7_mux_5_nl;
  wire[5:0] operator_6_false_7_mux_6_nl;
  wire operator_6_false_7_mux_7_nl;
  wire[5:0] operator_6_false_7_mux_8_nl;
  wire[1:0] return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_and_1_nl;
  wire[1:0] return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_mux_1_nl;
  wire not_906_nl;
  wire[9:0] return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_mux1h_2_nl;
  wire[13:0] acc_35_nl;
  wire[14:0] nl_acc_35_nl;
  wire[1:0] operator_6_false_15_operator_6_false_15_and_1_nl;
  wire operator_6_false_15_not_1_nl;
  wire[10:0] operator_6_false_15_mux_3_nl;
  wire[10:0] operator_32_false_2_acc_7_nl;
  wire[11:0] nl_operator_32_false_2_acc_7_nl;
  wire operator_6_false_15_or_1_nl;
  wire[5:0] operator_6_false_15_mux_4_nl;
  wire[3:0] BUTTERFLY_else_2_mux_5_nl;
  wire[12:0] BUTTERFLY_else_2_mux_6_nl;
  wire[15:0] BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_3_nl;
  wire[5:0] stage_u_add_3_mux_2_nl;
  wire[10:0] stage_u_add_3_mux_3_nl;
  wire[18:0] acc_39_nl;
  wire[19:0] nl_acc_39_nl;
  wire[3:0] stage_u_add_mux_5_nl;
  wire[1:0] stage_u_add_mux_6_nl;
  wire[10:0] stage_u_add_mux_7_nl;
  wire stage_u_add_or_5_nl;
  wire[13:0] acc_41_nl;
  wire[14:0] nl_acc_41_nl;
  wire[5:0] operator_6_false_43_mux_3_nl;
  wire[31:0] operator_32_false_1_acc_nl_1;
  wire[32:0] nl_operator_32_false_1_acc_nl_1;
  wire[17:0] operator_32_false_1_mux_4_nl;
  wire[17:0] operator_32_false_1_acc_7_nl;
  wire[18:0] nl_operator_32_false_1_acc_7_nl;
  wire[15:0] operator_32_false_1_acc_8_nl;
  wire[16:0] nl_operator_32_false_1_acc_8_nl;
  wire[1:0] operator_32_false_1_mux_5_nl;
  wire[3:0] operator_32_false_1_mux_6_nl;
  wire[5:0] operator_32_false_1_mux_7_nl;
  wire return_add_generic_AC_RND_CONV_false_8_op_bigger_mux_6_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_47_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_return_mult_generic_AC_RND_CONV_false_1_nor_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_return_mult_generic_AC_RND_CONV_false_2_nor_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_return_mult_generic_AC_RND_CONV_false_5_nor_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_and_5_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_and_6_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_and_7_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_and_8_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_and_9_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_and_10_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_and_11_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_and_12_nl;

  // Interconnect Declarations for Component Instantiations 
  wire return_mult_generic_AC_RND_CONV_false_1_if_return_mult_generic_AC_RND_CONV_false_1_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_mux_1_nl;
  wire[50:0] return_mult_generic_AC_RND_CONV_false_1_if_mux_2_nl;
  wire [52:0] nl_leading_sign_53_0_1_rg_mantissa;
  assign return_mult_generic_AC_RND_CONV_false_1_if_return_mult_generic_AC_RND_CONV_false_1_if_and_nl
      = return_extract_17_return_extract_17_or_sva_1 & BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm;
  assign return_mult_generic_AC_RND_CONV_false_1_if_mux_1_nl = MUX_s_1_2_2(stage_PE_1_tmp_im_d_1_lpi_3_dfm_51,
      return_add_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_1, BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm);
  assign return_mult_generic_AC_RND_CONV_false_1_if_mux_2_nl = MUX_v_51_2_2(stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0,
      return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1, BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm);
  assign nl_leading_sign_53_0_1_rg_mantissa = {return_mult_generic_AC_RND_CONV_false_1_if_return_mult_generic_AC_RND_CONV_false_1_if_and_nl
      , return_mult_generic_AC_RND_CONV_false_1_if_mux_1_nl , return_mult_generic_AC_RND_CONV_false_1_if_mux_2_nl};
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_3_lshift_1_rg_s;
  assign nl_return_add_generic_AC_RND_CONV_false_3_lshift_1_rg_s = MUX_v_6_2_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[5:0]),
      leading_sign_57_0_1_0_15_out_3, return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1);
  wire [56:0] nl_leading_sign_57_0_1_0_2_rg_mantissa;
  assign nl_leading_sign_57_0_1_0_2_rg_mantissa = {return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_0
      , return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_1 , return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_2};
  wire [5:0] nl_return_mult_generic_AC_RND_CONV_false_3_if_1_lshift_rg_s;
  assign nl_return_mult_generic_AC_RND_CONV_false_3_if_1_lshift_rg_s = MUX_v_6_2_2(leading_sign_53_0_out_1,
      (z_out_45[5:0]), z_out_63[12]);
  wire return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_2_nl;
  wire [52:0] nl_leading_sign_53_0_rg_mantissa;
  assign return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_2_nl
      = return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm & BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm;
  assign nl_leading_sign_53_0_rg_mantissa = {return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_2_nl
      , return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm , return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm};
  wire [5:0] nl_return_mult_generic_AC_RND_CONV_false_2_if_1_lshift_rg_s;
  assign nl_return_mult_generic_AC_RND_CONV_false_2_if_1_lshift_rg_s = MUX_v_6_2_2(leading_sign_53_0_2_out_1,
      (return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp[5:0]), operator_6_false_16_acc_psp_sva_1[12]);
  wire return_mult_generic_AC_RND_CONV_false_2_if_return_mult_generic_AC_RND_CONV_false_2_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_if_mux_1_nl;
  wire[50:0] return_mult_generic_AC_RND_CONV_false_2_if_mux_2_nl;
  wire [52:0] nl_leading_sign_53_0_2_rg_mantissa;
  assign return_mult_generic_AC_RND_CONV_false_2_if_return_mult_generic_AC_RND_CONV_false_2_if_and_nl
      = return_extract_19_return_extract_19_or_sva_1 & return_extract_41_return_extract_41_or_1_cse_sva;
  assign return_mult_generic_AC_RND_CONV_false_2_if_mux_1_nl = MUX_s_1_2_2((stage_PE_1_gm_im_d_61_0_lpi_3_dfm[51]),
      return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0, return_extract_41_return_extract_41_or_1_cse_sva);
  assign return_mult_generic_AC_RND_CONV_false_2_if_mux_2_nl = MUX_v_51_2_2((stage_PE_1_gm_im_d_61_0_lpi_3_dfm[50:0]),
      return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1, return_extract_41_return_extract_41_or_1_cse_sva);
  assign nl_leading_sign_53_0_2_rg_mantissa = {return_mult_generic_AC_RND_CONV_false_2_if_return_mult_generic_AC_RND_CONV_false_2_if_and_nl
      , return_mult_generic_AC_RND_CONV_false_2_if_mux_1_nl , return_mult_generic_AC_RND_CONV_false_2_if_mux_2_nl};
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_6_lshift_1_rg_s;
  assign nl_return_add_generic_AC_RND_CONV_false_6_lshift_1_rg_s = {return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_0
      , return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_1 , return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2};
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_7_rshift_rg_a;
  assign nl_return_add_generic_AC_RND_CONV_false_7_rshift_rg_a = {1'b0 , return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_52_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_0_lpi_3_dfm_mx0 , 3'b000};
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_7_lshift_1_rg_a;
  assign nl_return_add_generic_AC_RND_CONV_false_7_lshift_1_rg_a = {return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_0
      , return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_1 , return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_2};
  wire return_add_generic_AC_RND_CONV_false_7_mux_12_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_38_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_7_mux_39_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_7_lshift_1_rg_s;
  assign return_add_generic_AC_RND_CONV_false_7_mux_12_nl = MUX_s_1_2_2((reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[5]),
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_0, return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_7_mux_38_nl = MUX_s_1_2_2((reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[4]),
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_1, return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_7_mux_39_nl = MUX_v_4_2_2((reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[3:0]),
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2, return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1);
  assign nl_return_add_generic_AC_RND_CONV_false_7_lshift_1_rg_s = {return_add_generic_AC_RND_CONV_false_7_mux_12_nl
      , return_add_generic_AC_RND_CONV_false_7_mux_38_nl , return_add_generic_AC_RND_CONV_false_7_mux_39_nl};
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_17_lshift_3_rg_s;
  assign nl_return_add_generic_AC_RND_CONV_false_17_lshift_3_rg_s = MUX_v_6_2_2(reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2,
      leading_sign_57_0_1_0_17_out_3, return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10);
  wire return_mult_generic_AC_RND_CONV_false_4_if_return_mult_generic_AC_RND_CONV_false_4_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_if_mux_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_if_mux_2_nl;
  wire[49:0] return_mult_generic_AC_RND_CONV_false_4_if_mux_4_nl;
  wire [52:0] nl_leading_sign_53_0_4_rg_mantissa;
  assign return_mult_generic_AC_RND_CONV_false_4_if_return_mult_generic_AC_RND_CONV_false_4_if_and_nl
      = return_extract_49_return_extract_49_or_sva_1 & BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm;
  assign return_mult_generic_AC_RND_CONV_false_4_if_mux_1_nl = MUX_s_1_2_2(stage_PE_1_tmp_im_d_1_lpi_3_dfm_51,
      drf_qr_lval_14_smx_0_lpi_3_dfm, BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm);
  assign return_mult_generic_AC_RND_CONV_false_4_if_mux_2_nl = MUX_s_1_2_2((stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0[50]),
      return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_50, BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm);
  assign return_mult_generic_AC_RND_CONV_false_4_if_mux_4_nl = MUX_v_50_2_2((stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0[49:0]),
      return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0, BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm);
  assign nl_leading_sign_53_0_4_rg_mantissa = {return_mult_generic_AC_RND_CONV_false_4_if_return_mult_generic_AC_RND_CONV_false_4_if_and_nl
      , return_mult_generic_AC_RND_CONV_false_4_if_mux_1_nl , return_mult_generic_AC_RND_CONV_false_4_if_mux_2_nl
      , return_mult_generic_AC_RND_CONV_false_4_if_mux_4_nl};
  wire [5:0] nl_return_mult_generic_AC_RND_CONV_false_5_if_1_lshift_rg_s;
  assign nl_return_mult_generic_AC_RND_CONV_false_5_if_1_lshift_rg_s = MUX_v_6_2_2(leading_sign_53_0_5_out_1,
      (return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp[5:0]), operator_6_false_45_acc_psp_sva_1[12]);
  wire return_mult_generic_AC_RND_CONV_false_5_if_return_mult_generic_AC_RND_CONV_false_5_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_if_mux_1_nl;
  wire[50:0] return_mult_generic_AC_RND_CONV_false_5_if_mux_2_nl;
  wire [52:0] nl_leading_sign_53_0_5_rg_mantissa;
  assign return_mult_generic_AC_RND_CONV_false_5_if_return_mult_generic_AC_RND_CONV_false_5_if_and_nl
      = return_extract_51_return_extract_51_or_sva_1 & return_extract_41_return_extract_41_or_1_cse_sva;
  assign return_mult_generic_AC_RND_CONV_false_5_if_mux_1_nl = MUX_s_1_2_2((stage_PE_1_gm_im_d_61_0_lpi_3_dfm[51]),
      return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0, return_extract_41_return_extract_41_or_1_cse_sva);
  assign return_mult_generic_AC_RND_CONV_false_5_if_mux_2_nl = MUX_v_51_2_2((stage_PE_1_gm_im_d_61_0_lpi_3_dfm[50:0]),
      return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1, return_extract_41_return_extract_41_or_1_cse_sva);
  assign nl_leading_sign_53_0_5_rg_mantissa = {return_mult_generic_AC_RND_CONV_false_5_if_return_mult_generic_AC_RND_CONV_false_5_if_and_nl
      , return_mult_generic_AC_RND_CONV_false_5_if_mux_1_nl , return_mult_generic_AC_RND_CONV_false_5_if_mux_2_nl};
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_20_rshift_rg_a;
  assign nl_return_add_generic_AC_RND_CONV_false_20_rshift_rg_a = {1'b0 , return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_52_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_51_lpi_3_dfm_mx0 ,
      return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0 ,
      return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_0_lpi_3_dfm_mx0 , 3'b000};
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_25_rshift_rg_a;
  assign nl_return_add_generic_AC_RND_CONV_false_25_rshift_rg_a = {1'b0 , return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_52_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_51_lpi_3_dfm_mx0 ,
      return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0 ,
      return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_0_lpi_3_dfm_mx0 , 3'b000};
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_20_lshift_1_rg_s;
  assign nl_return_add_generic_AC_RND_CONV_false_20_lshift_1_rg_s = MUX_v_6_2_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[5:0]),
      return_add_generic_AC_RND_CONV_false_20_ls_sva, return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1);
  wire [3:0] nl_return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_rg_s;
  assign nl_return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_rg_s = ~ (z_out_51[3:0]);
  wire[51:0] return_mult_generic_AC_RND_CONV_false_6_if_return_mult_generic_AC_RND_CONV_false_6_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_op1_normal_not_5_nl;
  wire [52:0] nl_leading_sign_53_0_6_rg_mantissa;
  assign return_mult_generic_AC_RND_CONV_false_6_op1_normal_not_5_nl = ~ return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp;
  assign return_mult_generic_AC_RND_CONV_false_6_if_return_mult_generic_AC_RND_CONV_false_6_if_and_nl
      = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000, (out_f_d_rsci_q_d[51:0]),
      return_mult_generic_AC_RND_CONV_false_6_op1_normal_not_5_nl);
  assign nl_leading_sign_53_0_6_rg_mantissa = {return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp
      , return_mult_generic_AC_RND_CONV_false_6_if_return_mult_generic_AC_RND_CONV_false_6_if_and_nl};
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_3_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_13_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_1_mux1h_15_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_14_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_13_rshift_rg_a;
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_3_nl = MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_op_smaller_qr_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_52_lpi_3_dfm_mx0,
      {(fsm_output[6]) , (fsm_output[8]) , (fsm_output[22]) , (fsm_output[24]) ,
      (fsm_output[29])});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_13_nl = MUX1HOT_s_1_5_2((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      (return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_51_lpi_3_dfm_mx0, {(fsm_output[6])
      , (fsm_output[8]) , (fsm_output[22]) , (fsm_output[24]) , (fsm_output[29])});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_15_nl = MUX1HOT_v_50_5_2((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      (return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0, {(fsm_output[6])
      , (fsm_output[8]) , (fsm_output[22]) , (fsm_output[24]) , (fsm_output[29])});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_14_nl = MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_op_smaller_qr_0_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_0_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_0_lpi_3_dfm_mx0,
      {(fsm_output[6]) , (fsm_output[8]) , (fsm_output[22]) , (fsm_output[24]) ,
      (fsm_output[29])});
  assign nl_return_add_generic_AC_RND_CONV_false_13_rshift_rg_a = {1'b0 , return_add_generic_AC_RND_CONV_false_1_mux1h_3_nl
      , return_add_generic_AC_RND_CONV_false_1_mux1h_13_nl , return_add_generic_AC_RND_CONV_false_1_mux1h_15_nl
      , return_add_generic_AC_RND_CONV_false_1_mux1h_14_nl , 3'b000};
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_13_rshift_rg_s;
  assign nl_return_add_generic_AC_RND_CONV_false_13_rshift_rg_s = MUX1HOT_v_6_4_2(return_add_generic_AC_RND_CONV_false_1_e_dif_sat_or_cse,
      return_add_generic_AC_RND_CONV_false_2_e_dif_sat_or_cse, return_add_generic_AC_RND_CONV_false_e_dif_sat_or_cse,
      return_add_generic_AC_RND_CONV_false_23_e_dif_sat_sva_1, {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , (fsm_output[8]) , (fsm_output[24]) , (fsm_output[29])});
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_3_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_14_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_3_mux1h_16_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_15_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_15_rshift_rg_a;
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_3_nl = MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_op_smaller_qr_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_11_op_smaller_mux_cse,
      return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_52_lpi_3_dfm_mx0, {(fsm_output[6])
      , (fsm_output[8]) , (fsm_output[13]) , (fsm_output[22]) , (fsm_output[24])
      , (fsm_output[29])});
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_14_nl = MUX1HOT_s_1_6_2((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      (return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_cse, (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_51_lpi_3_dfm_mx0, {(fsm_output[6])
      , (fsm_output[8]) , (fsm_output[13]) , (fsm_output[22]) , (fsm_output[24])
      , (fsm_output[29])});
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_16_nl = MUX1HOT_v_50_6_2((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      (return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1, (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0, {(fsm_output[6])
      , (fsm_output[8]) , (fsm_output[13]) , (fsm_output[22]) , (fsm_output[24])
      , (fsm_output[29])});
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_15_nl = MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_op_smaller_qr_0_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_2_cse,
      return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_0_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_0_lpi_3_dfm_mx0, {(fsm_output[6])
      , (fsm_output[8]) , (fsm_output[13]) , (fsm_output[22]) , (fsm_output[24])
      , (fsm_output[29])});
  assign nl_return_add_generic_AC_RND_CONV_false_15_rshift_rg_a = {1'b0 , return_add_generic_AC_RND_CONV_false_3_mux1h_3_nl
      , return_add_generic_AC_RND_CONV_false_3_mux1h_14_nl , return_add_generic_AC_RND_CONV_false_3_mux1h_16_nl
      , return_add_generic_AC_RND_CONV_false_3_mux1h_15_nl , 3'b000};
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_15_rshift_rg_s;
  assign nl_return_add_generic_AC_RND_CONV_false_15_rshift_rg_s = MUX1HOT_v_6_5_2(return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse,
      return_add_generic_AC_RND_CONV_false_e_dif_sat_or_cse, return_add_generic_AC_RND_CONV_false_9_e_dif_sat_sva_1,
      return_add_generic_AC_RND_CONV_false_2_e_dif_sat_or_cse, return_add_generic_AC_RND_CONV_false_22_e_dif_sat_sva_1,
      {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , (fsm_output[8])
      , (fsm_output[13]) , (fsm_output[24]) , (fsm_output[29])});
  wire return_add_generic_AC_RND_CONV_false_5_mux_21_nl;
  wire return_add_generic_AC_RND_CONV_false_5_mux_22_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_5_mux_23_nl;
  wire return_add_generic_AC_RND_CONV_false_5_mux_24_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_a;
  assign return_add_generic_AC_RND_CONV_false_5_mux_21_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_1_cse, fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_5_mux_22_nl = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[50]),
      return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_cse, fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_5_mux_23_nl = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[49:0]),
      return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse, fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_5_mux_24_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_14_op1_mu_mux_1_cse, fsm_output[14]);
  assign nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_a = {1'b0 , return_add_generic_AC_RND_CONV_false_5_mux_21_nl
      , return_add_generic_AC_RND_CONV_false_5_mux_22_nl , return_add_generic_AC_RND_CONV_false_5_mux_23_nl
      , return_add_generic_AC_RND_CONV_false_5_mux_24_nl , 3'b000};
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_s;
  assign nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_s = {return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_0
      , return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_1 , return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2};
  wire return_add_generic_AC_RND_CONV_false_6_mux1h_2_nl;
  wire return_add_generic_AC_RND_CONV_false_6_mux1h_3_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_6_mux1h_5_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_11_rshift_rg_a;
  assign return_add_generic_AC_RND_CONV_false_6_mux1h_2_nl = MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_52_lpi_3_dfm_mx0,
      {(fsm_output[10]) , or_dcpl_104 , (fsm_output[26])});
  assign return_add_generic_AC_RND_CONV_false_6_mux1h_3_nl = MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_50_mx0,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_50_mx0,
      {(fsm_output[10]) , or_dcpl_104 , (fsm_output[26])});
  assign return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_mux_nl
      = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm, or_dcpl_104);
  assign return_add_generic_AC_RND_CONV_false_6_mux1h_5_nl = MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_0_lpi_3_dfm_mx0,
      {(fsm_output[10]) , or_dcpl_104 , (fsm_output[26])});
  assign nl_return_add_generic_AC_RND_CONV_false_11_rshift_rg_a = {1'b0 , return_add_generic_AC_RND_CONV_false_6_mux1h_2_nl
      , return_add_generic_AC_RND_CONV_false_6_mux1h_3_nl , return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_mux_nl
      , return_add_generic_AC_RND_CONV_false_6_mux1h_5_nl , 3'b000};
  wire[4:0] return_add_generic_AC_RND_CONV_false_6_mux1h_1_nl;
  wire return_add_generic_AC_RND_CONV_false_6_mux1h_6_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_11_rshift_rg_s;
  assign return_add_generic_AC_RND_CONV_false_6_mux1h_1_nl = MUX1HOT_v_5_3_2((return_add_generic_AC_RND_CONV_false_19_e_dif_sat_sva_1[5:1]),
      return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1_5_1, return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1_5_1,
      {or_1556_cse , (fsm_output[14]) , (fsm_output[16])});
  assign return_add_generic_AC_RND_CONV_false_6_mux1h_6_nl = MUX1HOT_s_1_3_2((return_add_generic_AC_RND_CONV_false_19_e_dif_sat_sva_1[0]),
      return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1_0, return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1_0,
      {or_1556_cse , (fsm_output[14]) , (fsm_output[16])});
  assign nl_return_add_generic_AC_RND_CONV_false_11_rshift_rg_s = {return_add_generic_AC_RND_CONV_false_6_mux1h_1_nl
      , return_add_generic_AC_RND_CONV_false_6_mux1h_6_nl};
  wire return_add_generic_AC_RND_CONV_false_8_mux_27_nl;
  wire return_add_generic_AC_RND_CONV_false_8_mux_29_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_8_mux_30_nl;
  wire return_add_generic_AC_RND_CONV_false_8_mux_31_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_21_rshift_rg_a;
  assign return_add_generic_AC_RND_CONV_false_8_mux_27_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_52_lpi_3_dfm_mx0, fsm_output[28]);
  assign return_add_generic_AC_RND_CONV_false_8_mux_29_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_51_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_51_lpi_3_dfm_mx0, fsm_output[28]);
  assign return_add_generic_AC_RND_CONV_false_8_mux_30_nl = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0, fsm_output[28]);
  assign return_add_generic_AC_RND_CONV_false_8_mux_31_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_0_lpi_3_dfm_mx0, fsm_output[28]);
  assign nl_return_add_generic_AC_RND_CONV_false_21_rshift_rg_a = {1'b0 , return_add_generic_AC_RND_CONV_false_8_mux_27_nl
      , return_add_generic_AC_RND_CONV_false_8_mux_29_nl , return_add_generic_AC_RND_CONV_false_8_mux_30_nl
      , return_add_generic_AC_RND_CONV_false_8_mux_31_nl , 3'b000};
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_21_rshift_rg_s;
  assign nl_return_add_generic_AC_RND_CONV_false_21_rshift_rg_s = MUX_v_6_2_2(return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1,
      return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1, fsm_output[28]);
  wire return_mult_generic_AC_RND_CONV_false_2_else_1_return_mult_generic_AC_RND_CONV_false_2_else_1_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_else_1_mux_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_else_1_return_mult_generic_AC_RND_CONV_false_2_else_1_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_else_1_mux_1_nl;
  wire[49:0] return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_4_nl;
  wire[1:0] return_mult_generic_AC_RND_CONV_false_2_else_1_return_mult_generic_AC_RND_CONV_false_2_else_1_and_2_nl;
  wire[1:0] return_mult_generic_AC_RND_CONV_false_2_else_1_mux_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_else_1_nor_2_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_17_rshift_1_rg_a;
  assign return_mult_generic_AC_RND_CONV_false_2_else_1_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_4_op_bigger_mux_3_cse,
      return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_52_lpi_3_dfm_mx0, fsm_output[29]);
  assign return_mult_generic_AC_RND_CONV_false_2_else_1_return_mult_generic_AC_RND_CONV_false_2_else_1_and_nl
      = return_mult_generic_AC_RND_CONV_false_2_else_1_mux_nl & return_mult_generic_AC_RND_CONV_false_2_else_1_nor_cse;
  assign return_mult_generic_AC_RND_CONV_false_2_else_1_mux_1_nl = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_51_lpi_3_dfm_mx0, fsm_output[29]);
  assign return_mult_generic_AC_RND_CONV_false_2_else_1_return_mult_generic_AC_RND_CONV_false_2_else_1_and_1_nl
      = return_mult_generic_AC_RND_CONV_false_2_else_1_mux_1_nl & return_mult_generic_AC_RND_CONV_false_2_else_1_nor_cse;
  assign return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_nl = MUX1HOT_v_50_4_2((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[105:56]),
      (return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[105:56]), (return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0, {(fsm_output[11])
      , (fsm_output[27]) , (fsm_output[22]) , (fsm_output[29])});
  assign return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_4_nl = MUX1HOT_s_1_4_2((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[55]),
      (return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[55]), return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_0_lpi_3_dfm_mx0, {(fsm_output[11])
      , (fsm_output[27]) , (fsm_output[22]) , (fsm_output[29])});
  assign return_mult_generic_AC_RND_CONV_false_2_else_1_mux_2_nl = MUX_v_2_2_2((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[54:53]),
      (return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[54:53]), fsm_output[27]);
  assign return_mult_generic_AC_RND_CONV_false_2_else_1_nor_2_nl = ~((fsm_output[22])
      | (fsm_output[29]));
  assign return_mult_generic_AC_RND_CONV_false_2_else_1_return_mult_generic_AC_RND_CONV_false_2_else_1_and_2_nl
      = MUX_v_2_2_2(2'b00, return_mult_generic_AC_RND_CONV_false_2_else_1_mux_2_nl,
      return_mult_generic_AC_RND_CONV_false_2_else_1_nor_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_17_rshift_1_rg_a = {1'b0 , return_mult_generic_AC_RND_CONV_false_2_else_1_return_mult_generic_AC_RND_CONV_false_2_else_1_and_nl
      , return_mult_generic_AC_RND_CONV_false_2_else_1_return_mult_generic_AC_RND_CONV_false_2_else_1_and_1_nl
      , return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_nl , return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_4_nl
      , return_mult_generic_AC_RND_CONV_false_2_else_1_return_mult_generic_AC_RND_CONV_false_2_else_1_and_2_nl
      , 1'b0};
  wire return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_1_nl;
  wire[3:0] return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_3_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_17_rshift_1_rg_s;
  assign return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_1_nl = MUX1HOT_s_1_4_2(return_mult_generic_AC_RND_CONV_false_2_shift_right_conc_3_5,
      return_mult_generic_AC_RND_CONV_false_5_shift_right_conc_3_5, (return_add_generic_AC_RND_CONV_false_4_e_dif_sat_or_cse[5]),
      (return_add_generic_AC_RND_CONV_false_24_e_dif_sat_sva_1[5]), {(fsm_output[11])
      , (fsm_output[27]) , (fsm_output[22]) , (fsm_output[29])});
  assign return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_2_nl = MUX1HOT_v_4_4_2(return_mult_generic_AC_RND_CONV_false_2_shift_right_conc_3_4_1,
      return_mult_generic_AC_RND_CONV_false_5_shift_right_conc_3_4_1, (return_add_generic_AC_RND_CONV_false_4_e_dif_sat_or_cse[4:1]),
      (return_add_generic_AC_RND_CONV_false_24_e_dif_sat_sva_1[4:1]), {(fsm_output[11])
      , (fsm_output[27]) , (fsm_output[22]) , (fsm_output[29])});
  assign return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_3_nl = MUX1HOT_s_1_4_2(return_mult_generic_AC_RND_CONV_false_2_shift_right_conc_3_0,
      return_mult_generic_AC_RND_CONV_false_5_shift_right_conc_3_0, (return_add_generic_AC_RND_CONV_false_4_e_dif_sat_or_cse[0]),
      (return_add_generic_AC_RND_CONV_false_24_e_dif_sat_sva_1[0]), {(fsm_output[11])
      , (fsm_output[27]) , (fsm_output[22]) , (fsm_output[29])});
  assign nl_return_add_generic_AC_RND_CONV_false_17_rshift_1_rg_s = {return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_1_nl
      , return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_2_nl , return_mult_generic_AC_RND_CONV_false_2_else_1_mux1h_3_nl};
  wire[50:0] return_mult_generic_AC_RND_CONV_false_1_else_1_return_mult_generic_AC_RND_CONV_false_1_else_1_mux_1_nl;
  wire [53:0] nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_a;
  assign return_mult_generic_AC_RND_CONV_false_1_else_1_return_mult_generic_AC_RND_CONV_false_1_else_1_mux_1_nl
      = MUX_v_51_2_2((z_out_26[103:53]), (out_f_d_rsci_q_d[51:1]), fsm_output[36]);
  assign nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_a = {return_mult_generic_AC_RND_CONV_false_1_else_1_and_1_cse
      , return_mult_generic_AC_RND_CONV_false_1_else_1_return_mult_generic_AC_RND_CONV_false_1_else_1_mux_2_cse
      , return_mult_generic_AC_RND_CONV_false_1_else_1_return_mult_generic_AC_RND_CONV_false_1_else_1_mux_1_nl
      , 1'b0};
  wire return_mult_generic_AC_RND_CONV_false_1_else_1_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_else_1_return_mult_generic_AC_RND_CONV_false_1_else_1_mux_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_else_1_return_mult_generic_AC_RND_CONV_false_1_else_1_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_else_1_mux_nl;
  wire[2:0] return_mult_generic_AC_RND_CONV_false_1_else_1_mux1h_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_else_1_mux1h_4_nl;
  wire [5:0] nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_s;
  assign return_mult_generic_AC_RND_CONV_false_1_else_1_return_mult_generic_AC_RND_CONV_false_1_else_1_mux_nl
      = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_1_shift_right_conc_3_5,
      return_mult_generic_AC_RND_CONV_false_if_or_3_cse, return_mult_generic_AC_RND_CONV_false_1_else_1_or_cse);
  assign return_mult_generic_AC_RND_CONV_false_1_else_1_and_nl = return_mult_generic_AC_RND_CONV_false_1_else_1_return_mult_generic_AC_RND_CONV_false_1_else_1_mux_nl
      & (~ (fsm_output[36]));
  assign return_mult_generic_AC_RND_CONV_false_1_else_1_mux_nl = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2[3]),
      (return_mult_generic_AC_RND_CONV_false_if_nand_1_cse[3]), return_mult_generic_AC_RND_CONV_false_1_else_1_or_cse);
  assign return_mult_generic_AC_RND_CONV_false_1_else_1_return_mult_generic_AC_RND_CONV_false_1_else_1_and_nl
      = return_mult_generic_AC_RND_CONV_false_1_else_1_mux_nl & (~ (fsm_output[36]));
  assign return_mult_generic_AC_RND_CONV_false_1_else_1_mux1h_3_nl = MUX1HOT_v_3_3_2((return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2[2:0]),
      (return_mult_generic_AC_RND_CONV_false_if_nand_1_cse[2:0]), (~ (z_out_51[3:1])),
      {(fsm_output[9]) , return_mult_generic_AC_RND_CONV_false_1_else_1_or_cse ,
      (fsm_output[36])});
  assign return_mult_generic_AC_RND_CONV_false_1_else_1_mux1h_4_nl = MUX1HOT_s_1_3_2(return_mult_generic_AC_RND_CONV_false_1_shift_right_conc_3_0,
      return_mult_generic_AC_RND_CONV_false_if_or_cse, (~ (z_out_51[0])), {(fsm_output[9])
      , return_mult_generic_AC_RND_CONV_false_1_else_1_or_cse , (fsm_output[36])});
  assign nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_s = {return_mult_generic_AC_RND_CONV_false_1_else_1_and_nl
      , return_mult_generic_AC_RND_CONV_false_1_else_1_return_mult_generic_AC_RND_CONV_false_1_else_1_and_nl
      , return_mult_generic_AC_RND_CONV_false_1_else_1_mux1h_3_nl , return_mult_generic_AC_RND_CONV_false_1_else_1_mux1h_4_nl};
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_1_lshift_1_rg_a;
  assign nl_return_add_generic_AC_RND_CONV_false_1_lshift_1_rg_a = {return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_0
      , return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_1 , return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_2};
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_5_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_16_nl;
  wire[2:0] return_add_generic_AC_RND_CONV_false_1_mux1h_17_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_18_nl;
  wire return_add_generic_AC_RND_CONV_false_1_or_nl;
  wire return_add_generic_AC_RND_CONV_false_1_and_52_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_1_lshift_1_rg_s;
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_5_nl = MUX1HOT_s_1_5_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[5]),
      (leading_sign_57_0_1_0_2_out_3[5]), (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[5]),
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_0, (return_add_generic_AC_RND_CONV_false_9_conc_59_itm_5_1[4]),
      {return_add_generic_AC_RND_CONV_false_1_and_itm , return_add_generic_AC_RND_CONV_false_1_and_1_itm
      , return_add_generic_AC_RND_CONV_false_1_and_2_itm , return_add_generic_AC_RND_CONV_false_1_and_3_itm
      , or_tmp_567});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_16_nl = MUX1HOT_s_1_5_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[4]),
      (leading_sign_57_0_1_0_2_out_3[4]), (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[4]),
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_1, (return_add_generic_AC_RND_CONV_false_9_conc_59_itm_5_1[3]),
      {return_add_generic_AC_RND_CONV_false_1_and_itm , return_add_generic_AC_RND_CONV_false_1_and_1_itm
      , return_add_generic_AC_RND_CONV_false_1_and_2_itm , return_add_generic_AC_RND_CONV_false_1_and_3_itm
      , or_tmp_567});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_17_nl = MUX1HOT_v_3_5_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[3:1]),
      (leading_sign_57_0_1_0_2_out_3[3:1]), (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[3:1]),
      (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2[3:1]), (return_add_generic_AC_RND_CONV_false_9_conc_59_itm_5_1[2:0]),
      {return_add_generic_AC_RND_CONV_false_1_and_itm , return_add_generic_AC_RND_CONV_false_1_and_1_itm
      , return_add_generic_AC_RND_CONV_false_1_and_2_itm , return_add_generic_AC_RND_CONV_false_1_and_3_itm
      , or_tmp_567});
  assign return_add_generic_AC_RND_CONV_false_1_or_nl = return_add_generic_AC_RND_CONV_false_1_and_1_itm
      | (return_add_generic_AC_RND_CONV_false_22_acc_3_itm_11_1 & or_tmp_567);
  assign return_add_generic_AC_RND_CONV_false_1_and_52_nl = (~ return_add_generic_AC_RND_CONV_false_22_acc_3_itm_11_1)
      & or_tmp_567;
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_18_nl = MUX1HOT_s_1_5_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[0]),
      (leading_sign_57_0_1_0_2_out_3[0]), (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[0]),
      (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2[0]), drf_qr_lval_12_smx_0_lpi_3_dfm,
      {return_add_generic_AC_RND_CONV_false_1_and_itm , return_add_generic_AC_RND_CONV_false_1_or_nl
      , return_add_generic_AC_RND_CONV_false_1_and_2_itm , return_add_generic_AC_RND_CONV_false_1_and_3_itm
      , return_add_generic_AC_RND_CONV_false_1_and_52_nl});
  assign nl_return_add_generic_AC_RND_CONV_false_1_lshift_1_rg_s = {return_add_generic_AC_RND_CONV_false_1_mux1h_5_nl
      , return_add_generic_AC_RND_CONV_false_1_mux1h_16_nl , return_add_generic_AC_RND_CONV_false_1_mux1h_17_nl
      , return_add_generic_AC_RND_CONV_false_1_mux1h_18_nl};
  wire return_add_generic_AC_RND_CONV_false_5_or_2_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_21_lshift_rg_a;
  assign return_add_generic_AC_RND_CONV_false_5_or_2_nl = (fsm_output[12]) | (fsm_output[28]);
  assign nl_return_add_generic_AC_RND_CONV_false_21_lshift_rg_a = MUX_v_57_2_2(return_add_generic_AC_RND_CONV_false_15_res_mant_4_sva,
      57'b001111111111111111111111111111111111111111111111111111111, return_add_generic_AC_RND_CONV_false_5_or_2_nl);
  wire return_add_generic_AC_RND_CONV_false_5_and_nl;
  wire return_add_generic_AC_RND_CONV_false_5_and_1_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_21_lshift_rg_s;
  assign return_add_generic_AC_RND_CONV_false_5_and_nl = (~ return_add_generic_AC_RND_CONV_false_5_acc_2_itm_10_1)
      & (fsm_output[8]);
  assign return_add_generic_AC_RND_CONV_false_5_and_1_nl = return_add_generic_AC_RND_CONV_false_5_acc_2_itm_10_1
      & (fsm_output[8]);
  assign nl_return_add_generic_AC_RND_CONV_false_21_lshift_rg_s = MUX1HOT_v_6_4_2(({(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0[4:0])
      , reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1}), return_add_generic_AC_RND_CONV_false_20_ls_sva,
      return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1, return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1,
      {return_add_generic_AC_RND_CONV_false_5_and_nl , return_add_generic_AC_RND_CONV_false_5_and_1_nl
      , (fsm_output[12]) , (fsm_output[28])});
  wire return_add_generic_AC_RND_CONV_false_3_or_nl;
  wire return_add_generic_AC_RND_CONV_false_3_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_3_or_3_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_15_lshift_rg_a;
  assign return_add_generic_AC_RND_CONV_false_3_or_nl = (fsm_output[6]) | (fsm_output[8])
      | (fsm_output[22]) | (fsm_output[24]) | (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_3_or_2_nl = (fsm_output[9]) | (fsm_output[11])
      | (fsm_output[27]);
  assign return_add_generic_AC_RND_CONV_false_3_or_3_nl = (fsm_output[23]) | (fsm_output[30]);
  assign nl_return_add_generic_AC_RND_CONV_false_15_lshift_rg_a = MUX1HOT_v_57_3_2(57'b001111111111111111111111111111111111111111111111111111111,
      57'b000011111111111111111111111111111111111111111111111111111, z_out_6, {return_add_generic_AC_RND_CONV_false_3_or_nl
      , return_add_generic_AC_RND_CONV_false_3_or_2_nl , return_add_generic_AC_RND_CONV_false_3_or_3_nl});
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_6_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_3_mux1h_12_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_13_nl;
  wire return_add_generic_AC_RND_CONV_false_3_and_28_nl;
  wire return_add_generic_AC_RND_CONV_false_3_and_29_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_15_lshift_rg_s;
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_6_nl = MUX1HOT_s_1_8_2((return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse[5]),
      (return_add_generic_AC_RND_CONV_false_2_e_dif_sat_or_cse[5]), return_mult_generic_AC_RND_CONV_false_1_shift_right_conc_3_5,
      return_mult_generic_AC_RND_CONV_false_2_shift_right_conc_3_5, (return_add_generic_AC_RND_CONV_false_18_mux_4_itm[5]),
      return_mult_generic_AC_RND_CONV_false_5_shift_right_conc_3_5, (return_add_generic_AC_RND_CONV_false_24_e_dif_sat_sva_1[5]),
      (return_add_generic_AC_RND_CONV_false_24_mux_4_itm_5_1[4]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , or_1495_cse_1 , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[23]) , (fsm_output[27])
      , (fsm_output[29]) , (fsm_output[30])});
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_12_nl = MUX1HOT_v_4_8_2((return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse[4:1]),
      (return_add_generic_AC_RND_CONV_false_2_e_dif_sat_or_cse[4:1]), return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2,
      return_mult_generic_AC_RND_CONV_false_2_shift_right_conc_3_4_1, (return_add_generic_AC_RND_CONV_false_18_mux_4_itm[4:1]),
      return_mult_generic_AC_RND_CONV_false_5_shift_right_conc_3_4_1, (return_add_generic_AC_RND_CONV_false_24_e_dif_sat_sva_1[4:1]),
      (return_add_generic_AC_RND_CONV_false_24_mux_4_itm_5_1[3:0]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , or_1495_cse_1 , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[23]) , (fsm_output[27])
      , (fsm_output[29]) , (fsm_output[30])});
  assign return_add_generic_AC_RND_CONV_false_3_and_28_nl = (~ return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11)
      & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_3_and_29_nl = return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11
      & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_13_nl = MUX1HOT_s_1_9_2((return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse[0]),
      (return_add_generic_AC_RND_CONV_false_2_e_dif_sat_or_cse[0]), return_mult_generic_AC_RND_CONV_false_1_shift_right_conc_3_0,
      return_mult_generic_AC_RND_CONV_false_2_shift_right_conc_3_0, (return_add_generic_AC_RND_CONV_false_18_mux_4_itm[0]),
      return_mult_generic_AC_RND_CONV_false_5_shift_right_conc_3_0, (return_add_generic_AC_RND_CONV_false_24_e_dif_sat_sva_1[0]),
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm, (leading_sign_57_0_1_0_24_out_3[0]),
      {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , or_1495_cse_1
      , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[23]) , (fsm_output[27])
      , (fsm_output[29]) , return_add_generic_AC_RND_CONV_false_3_and_28_nl , return_add_generic_AC_RND_CONV_false_3_and_29_nl});
  assign nl_return_add_generic_AC_RND_CONV_false_15_lshift_rg_s = {return_add_generic_AC_RND_CONV_false_3_mux1h_6_nl
      , return_add_generic_AC_RND_CONV_false_3_mux1h_12_nl , return_add_generic_AC_RND_CONV_false_3_mux1h_13_nl};
  wire[3:0] return_add_generic_AC_RND_CONV_false_5_mux1h_2_nl;
  wire[1:0] return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_or_nl;
  wire[1:0] return_add_generic_AC_RND_CONV_false_5_mux_25_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_or_1_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_5_mux_26_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_a;
  assign return_add_generic_AC_RND_CONV_false_5_mux1h_2_nl = MUX1HOT_v_4_3_2(4'b0011,
      (return_add_generic_AC_RND_CONV_false_15_res_mant_4_sva[56:53]), return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_0,
      {return_add_generic_AC_RND_CONV_false_20_ls_or_cse , or_dcpl_147 , return_add_generic_AC_RND_CONV_false_5_or_1_itm});
  assign return_add_generic_AC_RND_CONV_false_5_mux_25_nl = MUX_v_2_2_2((return_add_generic_AC_RND_CONV_false_15_res_mant_4_sva[52:51]),
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_1, return_add_generic_AC_RND_CONV_false_5_or_1_itm);
  assign return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_or_nl
      = MUX_v_2_2_2(return_add_generic_AC_RND_CONV_false_5_mux_25_nl, 2'b11, return_add_generic_AC_RND_CONV_false_20_ls_or_cse);
  assign return_add_generic_AC_RND_CONV_false_5_mux_26_nl = MUX_v_51_2_2((return_add_generic_AC_RND_CONV_false_15_res_mant_4_sva[50:0]),
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_2, return_add_generic_AC_RND_CONV_false_5_or_1_itm);
  assign return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_or_1_nl
      = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_5_mux_26_nl, 51'b111111111111111111111111111111111111111111111111111,
      return_add_generic_AC_RND_CONV_false_20_ls_or_cse);
  assign nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_a = {return_add_generic_AC_RND_CONV_false_5_mux1h_2_nl
      , return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_or_nl
      , return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_or_1_nl};
  wire return_add_generic_AC_RND_CONV_false_5_mux1h_3_nl;
  wire return_add_generic_AC_RND_CONV_false_5_mux1h_5_nl;
  wire[2:0] return_add_generic_AC_RND_CONV_false_5_mux1h_6_nl;
  wire return_add_generic_AC_RND_CONV_false_5_mux1h_4_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_s;
  assign return_add_generic_AC_RND_CONV_false_5_mux1h_3_nl = MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_0,
      (return_add_generic_AC_RND_CONV_false_8_mux_8_itm[5]), (in_u_rsc_merge_sva_rsp_1_rsp_1[4]),
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_1, (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[4]),
      (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[5]), {return_add_generic_AC_RND_CONV_false_5_or_4_cse
      , (fsm_output[13]) , return_add_generic_AC_RND_CONV_false_5_and_6_cse , (fsm_output[16])
      , return_add_generic_AC_RND_CONV_false_5_and_8_cse , return_add_generic_AC_RND_CONV_false_5_and_10_cse});
  assign return_add_generic_AC_RND_CONV_false_5_mux1h_5_nl = MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_1,
      (return_add_generic_AC_RND_CONV_false_8_mux_8_itm[4]), (in_u_rsc_merge_sva_rsp_1_rsp_1[3]),
      (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2[3]), (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[3]),
      (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[4]), {return_add_generic_AC_RND_CONV_false_5_or_4_cse
      , (fsm_output[13]) , return_add_generic_AC_RND_CONV_false_5_and_6_cse , (fsm_output[16])
      , return_add_generic_AC_RND_CONV_false_5_and_8_cse , return_add_generic_AC_RND_CONV_false_5_and_10_cse});
  assign return_add_generic_AC_RND_CONV_false_5_mux1h_6_nl = MUX1HOT_v_3_6_2((return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2[3:1]),
      (return_add_generic_AC_RND_CONV_false_8_mux_8_itm[3:1]), (in_u_rsc_merge_sva_rsp_1_rsp_1[2:0]),
      (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2[2:0]), (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[2:0]),
      (return_add_generic_AC_RND_CONV_false_21_mux_8_itm_3_0[3:1]), {return_add_generic_AC_RND_CONV_false_5_or_6_cse
      , (fsm_output[13]) , return_add_generic_AC_RND_CONV_false_5_and_6_cse , (fsm_output[16])
      , return_add_generic_AC_RND_CONV_false_5_and_8_cse , (fsm_output[29])});
  assign return_add_generic_AC_RND_CONV_false_5_mux1h_4_nl = MUX1HOT_s_1_6_2((return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2[0]),
      (return_add_generic_AC_RND_CONV_false_8_mux_8_itm[0]), return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm,
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm, drf_qr_lval_12_smx_0_lpi_3_dfm,
      (return_add_generic_AC_RND_CONV_false_21_mux_8_itm_3_0[0]), {return_add_generic_AC_RND_CONV_false_5_or_6_cse
      , (fsm_output[13]) , return_add_generic_AC_RND_CONV_false_5_and_6_cse , (fsm_output[16])
      , return_add_generic_AC_RND_CONV_false_5_and_8_cse , (fsm_output[29])});
  assign nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_s = {return_add_generic_AC_RND_CONV_false_5_mux1h_3_nl
      , return_add_generic_AC_RND_CONV_false_5_mux1h_5_nl , return_add_generic_AC_RND_CONV_false_5_mux1h_6_nl
      , return_add_generic_AC_RND_CONV_false_5_mux1h_4_nl};
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_13_lshift_rg_a;
  assign nl_return_add_generic_AC_RND_CONV_false_13_lshift_rg_a = MUX_v_57_2_2(57'b001111111111111111111111111111111111111111111111111111111,
      z_out_5, fsm_output[30]);
  wire[4:0] return_add_generic_AC_RND_CONV_false_1_mux1h_7_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_19_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_13_lshift_rg_s;
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_7_nl = MUX1HOT_v_5_6_2((return_add_generic_AC_RND_CONV_false_1_e_dif_sat_or_cse[5:1]),
      (return_add_generic_AC_RND_CONV_false_e_dif_sat_or_cse[5:1]), (return_add_generic_AC_RND_CONV_false_9_e_dif_sat_sva_1[5:1]),
      (return_add_generic_AC_RND_CONV_false_22_e_dif_sat_sva_1[5:1]), (in_u_rsc_merge_sva_rsp_1_rsp_1[4:0]),
      (leading_sign_57_0_1_0_25_out_3[5:1]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , or_1495_cse_1 , (fsm_output[13]) , (fsm_output[29]) , return_add_generic_AC_RND_CONV_false_1_and_54_cse
      , return_add_generic_AC_RND_CONV_false_1_and_55_cse});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_19_nl = MUX1HOT_s_1_6_2((return_add_generic_AC_RND_CONV_false_1_e_dif_sat_or_cse[0]),
      (return_add_generic_AC_RND_CONV_false_e_dif_sat_or_cse[0]), (return_add_generic_AC_RND_CONV_false_9_e_dif_sat_sva_1[0]),
      (return_add_generic_AC_RND_CONV_false_22_e_dif_sat_sva_1[0]), return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm,
      (leading_sign_57_0_1_0_25_out_3[0]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , or_1495_cse_1 , (fsm_output[13]) , (fsm_output[29]) , return_add_generic_AC_RND_CONV_false_1_and_54_cse
      , return_add_generic_AC_RND_CONV_false_1_and_55_cse});
  assign nl_return_add_generic_AC_RND_CONV_false_13_lshift_rg_s = {return_add_generic_AC_RND_CONV_false_1_mux1h_7_nl
      , return_add_generic_AC_RND_CONV_false_1_mux1h_19_nl};
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_23_lshift_1_rg_a;
  assign nl_return_add_generic_AC_RND_CONV_false_23_lshift_1_rg_a = MUX_v_57_2_2(57'b000011111111111111111111111111111111111111111111111111111,
      return_add_generic_AC_RND_CONV_false_15_res_mant_4_sva, fsm_output[30]);
  wire return_mult_generic_AC_RND_CONV_false_4_else_1_return_mult_generic_AC_RND_CONV_false_4_else_1_mux_1_nl;
  wire[2:0] return_mult_generic_AC_RND_CONV_false_4_else_1_return_mult_generic_AC_RND_CONV_false_4_else_1_mux_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_else_1_return_mult_generic_AC_RND_CONV_false_4_else_1_mux_3_nl;
  wire return_add_generic_AC_RND_CONV_false_23_mux_29_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_else_1_mux1h_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_else_1_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_else_1_and_1_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_23_lshift_1_rg_s;
  assign return_mult_generic_AC_RND_CONV_false_4_else_1_return_mult_generic_AC_RND_CONV_false_4_else_1_mux_1_nl
      = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_if_or_3_cse, (return_add_generic_AC_RND_CONV_false_23_mux_11_itm_5_2[3]),
      fsm_output[30]);
  assign return_mult_generic_AC_RND_CONV_false_4_else_1_return_mult_generic_AC_RND_CONV_false_4_else_1_mux_2_nl
      = MUX_v_3_2_2((return_mult_generic_AC_RND_CONV_false_if_nand_1_cse[3:1]), (return_add_generic_AC_RND_CONV_false_23_mux_11_itm_5_2[2:0]),
      fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_23_mux_29_nl = MUX_s_1_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1,
      (leading_sign_57_0_1_0_15_out_3[1]), return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1);
  assign return_mult_generic_AC_RND_CONV_false_4_else_1_return_mult_generic_AC_RND_CONV_false_4_else_1_mux_3_nl
      = MUX_s_1_2_2((return_mult_generic_AC_RND_CONV_false_if_nand_1_cse[0]), return_add_generic_AC_RND_CONV_false_23_mux_29_nl,
      fsm_output[30]);
  assign return_mult_generic_AC_RND_CONV_false_4_else_1_and_nl = (~ return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1)
      & (fsm_output[30]);
  assign return_mult_generic_AC_RND_CONV_false_4_else_1_and_1_nl = return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1
      & (fsm_output[30]);
  assign return_mult_generic_AC_RND_CONV_false_4_else_1_mux1h_3_nl = MUX1HOT_s_1_3_2(return_mult_generic_AC_RND_CONV_false_if_or_cse,
      drf_qr_lval_14_smx_0_lpi_3_dfm, (leading_sign_57_0_1_0_15_out_3[0]), {return_mult_generic_AC_RND_CONV_false_1_else_1_or_cse
      , return_mult_generic_AC_RND_CONV_false_4_else_1_and_nl , return_mult_generic_AC_RND_CONV_false_4_else_1_and_1_nl});
  assign nl_return_add_generic_AC_RND_CONV_false_23_lshift_1_rg_s = {return_mult_generic_AC_RND_CONV_false_4_else_1_return_mult_generic_AC_RND_CONV_false_4_else_1_mux_1_nl
      , return_mult_generic_AC_RND_CONV_false_4_else_1_return_mult_generic_AC_RND_CONV_false_4_else_1_mux_2_nl
      , return_mult_generic_AC_RND_CONV_false_4_else_1_return_mult_generic_AC_RND_CONV_false_4_else_1_mux_3_nl
      , return_mult_generic_AC_RND_CONV_false_4_else_1_mux1h_3_nl};
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_17_lshift_1_rg_s;
  assign nl_return_add_generic_AC_RND_CONV_false_17_lshift_1_rg_s = MUX_v_6_2_2(return_add_generic_AC_RND_CONV_false_4_e_dif_sat_or_cse,
      return_add_generic_AC_RND_CONV_false_25_e_dif_sat_sva_1, fsm_output[29]);
  wire[4:0] return_add_generic_AC_RND_CONV_false_11_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_11_mux_24_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_11_lshift_rg_s;
  assign return_add_generic_AC_RND_CONV_false_11_mux_nl = MUX_v_5_2_2(return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1_5_1,
      return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1_5_1, fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_11_mux_24_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1_0,
      return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1_0, fsm_output[16]);
  assign nl_return_add_generic_AC_RND_CONV_false_11_lshift_rg_s = {return_add_generic_AC_RND_CONV_false_11_mux_nl
      , return_add_generic_AC_RND_CONV_false_11_mux_24_nl};
  wire [56:0] nl_leading_sign_57_0_1_0_11_rg_mantissa;
  assign nl_leading_sign_57_0_1_0_11_rg_mantissa = MUX_v_57_2_2(return_add_generic_AC_RND_CONV_false_5_res_mant_4_sva_1,
      z_out_9, fsm_output[14]);
  wire[51:0] return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_mux_2_nl;
  wire[51:0] return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_not_1_nl;
  wire [105:0] nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_a;
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_mux_2_nl
      = MUX_v_52_2_2((z_out_26[103:52]), (out_f_d_rsci_q_d[51:0]), fsm_output[36]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_not_1_nl = ~ (fsm_output[36]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_nl
      = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000, (z_out_26[51:0]),
      return_mult_generic_AC_RND_CONV_false_1_if_1_not_1_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_a = {return_mult_generic_AC_RND_CONV_false_1_else_1_and_1_cse
      , return_mult_generic_AC_RND_CONV_false_1_else_1_return_mult_generic_AC_RND_CONV_false_1_else_1_mux_2_cse
      , return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_mux_2_nl
      , return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_nl};
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_and_4_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_and_5_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_and_6_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_and_7_nl;
  wire [5:0] nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_s;
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_and_2_nl = (~ (z_out_57[12]))
      & (fsm_output[9]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_and_3_nl = (z_out_57[12]) &
      (fsm_output[9]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_and_4_nl = (~ (z_out_63[12]))
      & (fsm_output[24]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_and_5_nl = (z_out_63[12]) &
      (fsm_output[24]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_and_6_nl = (~ (operator_6_false_58_acc_psp_sva_1[11]))
      & (fsm_output[36]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_and_7_nl = (operator_6_false_58_acc_psp_sva_1[11])
      & (fsm_output[36]);
  assign nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_s = MUX1HOT_v_6_6_2(return_add_generic_AC_RND_CONV_false_20_ls_sva,
      (stage_u_add_3_acc_itm_rsp_1[5:0]), leading_sign_53_0_4_out_1, (z_out_45[5:0]),
      leading_sign_53_0_6_out_1, (z_out_51[5:0]), {return_mult_generic_AC_RND_CONV_false_1_if_1_and_2_nl
      , return_mult_generic_AC_RND_CONV_false_1_if_1_and_3_nl , return_mult_generic_AC_RND_CONV_false_1_if_1_and_4_nl
      , return_mult_generic_AC_RND_CONV_false_1_if_1_and_5_nl , return_mult_generic_AC_RND_CONV_false_1_if_1_and_6_nl
      , return_mult_generic_AC_RND_CONV_false_1_if_1_and_7_nl});
  wire [79:0] nl_stage_run_out1_rsci_inst_out1_rsci_idat;
  assign nl_stage_run_out1_rsci_inst_out1_rsci_idat = {out1_rsci_idat_79_64 , out1_rsci_idat_63
      , out1_rsci_idat_62_52 , out1_rsci_idat_51 , out1_rsci_idat_50_0};
  wire  nl_stage_run_run_fsm_inst_for_C_0_tr0;
  assign nl_stage_run_run_fsm_inst_for_C_0_tr0 = for_i_3_0_sva[0];
  wire  nl_stage_run_run_fsm_inst_BUTTERFLY_C_15_tr0;
  assign nl_stage_run_run_fsm_inst_BUTTERFLY_C_15_tr0 = (nor_tmp | (z_out_49[9]))
      & or_dcpl_60;
  wire  nl_stage_run_run_fsm_inst_BUTTERFLY_1_C_15_tr0;
  assign nl_stage_run_run_fsm_inst_BUTTERFLY_1_C_15_tr0 = (nor_tmp | (BUTTERFLY_mux_5_itm_9_0[9]))
      & or_dcpl_60;
  wire  nl_stage_run_run_fsm_inst_for_1_C_2_tr0;
  assign nl_stage_run_run_fsm_inst_for_1_C_2_tr0 = z_out_55[10];
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd16)) mode1_rsci (
      .dat(mode1_rsc_dat),
      .idat(mode1_rsci_idat)
    );
  leading_sign_53_0  leading_sign_53_0_1_rg (
      .mantissa(nl_leading_sign_53_0_1_rg_mantissa[52:0]),
      .rtn(leading_sign_53_0_1_out_1)
    );
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_3_lshift_1_rg (
      .a(return_add_generic_AC_RND_CONV_false_15_res_mant_4_sva),
      .s(nl_return_add_generic_AC_RND_CONV_false_3_lshift_1_rg_s[5:0]),
      .z(return_add_generic_AC_RND_CONV_false_3_res_rounded_asn_rndc_sva_1)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_15_rg (
      .mantissa(return_add_generic_AC_RND_CONV_false_15_res_mant_4_sva),
      .all_same(leading_sign_57_0_1_0_15_out_2),
      .rtn(leading_sign_57_0_1_0_15_out_3)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_2_rg (
      .mantissa(nl_leading_sign_57_0_1_0_2_rg_mantissa[56:0]),
      .all_same(leading_sign_57_0_1_0_2_out_2),
      .rtn(leading_sign_57_0_1_0_2_out_3)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_4_rg (
      .mantissa(return_add_generic_AC_RND_CONV_false_4_res_mant_4_sva_1),
      .all_same(leading_sign_57_0_1_0_4_out_2),
      .rtn(leading_sign_57_0_1_0_4_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd106),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd106)) return_mult_generic_AC_RND_CONV_false_3_if_1_lshift_rg (
      .a(z_out_26),
      .s(nl_return_mult_generic_AC_RND_CONV_false_3_if_1_lshift_rg_s[5:0]),
      .z(return_mult_generic_AC_RND_CONV_false_3_p_sva_1)
    );
  leading_sign_53_0  leading_sign_53_0_rg (
      .mantissa(nl_leading_sign_53_0_rg_mantissa[52:0]),
      .rtn(leading_sign_53_0_out_1)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_6_rg (
      .mantissa(return_add_generic_AC_RND_CONV_false_6_res_mant_4_sva_1),
      .all_same(leading_sign_57_0_1_0_6_out_2),
      .rtn(leading_sign_57_0_1_0_6_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd106),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd106)) return_mult_generic_AC_RND_CONV_false_2_if_1_lshift_rg (
      .a(return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1),
      .s(nl_return_mult_generic_AC_RND_CONV_false_2_if_1_lshift_rg_s[5:0]),
      .z(return_mult_generic_AC_RND_CONV_false_2_p_sva_1)
    );
  leading_sign_53_0  leading_sign_53_0_2_rg (
      .mantissa(nl_leading_sign_53_0_2_rg_mantissa[52:0]),
      .rtn(leading_sign_53_0_2_out_1)
    );
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_6_lshift_1_rg (
      .a(return_add_generic_AC_RND_CONV_false_15_res_mant_4_sva),
      .s(nl_return_add_generic_AC_RND_CONV_false_6_lshift_1_rg_s[5:0]),
      .z(return_add_generic_AC_RND_CONV_false_6_res_rounded_asn_rndc_sva_1)
    );
  mgc_shift_r_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_7_rshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_7_rshift_rg_a[56:0]),
      .s(return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1),
      .z(return_add_generic_AC_RND_CONV_false_7_rshift_itm)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_8_rg (
      .mantissa(return_add_generic_AC_RND_CONV_false_8_res_mant_4_sva_1),
      .all_same(leading_sign_57_0_1_0_8_out_2),
      .rtn(leading_sign_57_0_1_0_8_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd55),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd55)) return_add_generic_AC_RND_CONV_false_7_lshift_rg (
      .a(55'b1111111111111111111111111111111111111111111111111111111),
      .s(return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1),
      .z(return_add_generic_AC_RND_CONV_false_7_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_7_lshift_1_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_7_lshift_1_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_7_lshift_1_rg_s[5:0]),
      .z(return_add_generic_AC_RND_CONV_false_7_res_rounded_asn_rndc_sva_1)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_10_rg (
      .mantissa(return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_2),
      .all_same(leading_sign_57_0_1_0_10_out_2),
      .rtn(leading_sign_57_0_1_0_10_out_3)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_18_rg (
      .mantissa(z_out_6),
      .all_same(leading_sign_57_0_1_0_18_out_2),
      .rtn(leading_sign_57_0_1_0_18_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_17_lshift_3_rg (
      .a(z_out_5),
      .s(nl_return_add_generic_AC_RND_CONV_false_17_lshift_3_rg_s[5:0]),
      .z(return_add_generic_AC_RND_CONV_false_17_res_rounded_asn_rndc_sva_1)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_17_rg (
      .mantissa(z_out_5),
      .all_same(leading_sign_57_0_1_0_17_out_2),
      .rtn(leading_sign_57_0_1_0_17_out_3)
    );
  leading_sign_53_0  leading_sign_53_0_4_rg (
      .mantissa(nl_leading_sign_53_0_4_rg_mantissa[52:0]),
      .rtn(leading_sign_53_0_4_out_1)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_19_rg (
      .mantissa(z_out_9),
      .all_same(leading_sign_57_0_1_0_19_out_2),
      .rtn(leading_sign_57_0_1_0_19_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd106),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd106)) return_mult_generic_AC_RND_CONV_false_5_if_1_lshift_rg (
      .a(return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1),
      .s(nl_return_mult_generic_AC_RND_CONV_false_5_if_1_lshift_rg_s[5:0]),
      .z(return_mult_generic_AC_RND_CONV_false_5_p_sva_1)
    );
  leading_sign_53_0  leading_sign_53_0_5_rg (
      .mantissa(nl_leading_sign_53_0_5_rg_mantissa[52:0]),
      .rtn(leading_sign_53_0_5_out_1)
    );
  mgc_shift_r_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_20_rshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_20_rshift_rg_a[56:0]),
      .s(return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1),
      .z(return_add_generic_AC_RND_CONV_false_20_rshift_itm)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_21_rg (
      .mantissa(return_add_generic_AC_RND_CONV_false_21_res_mant_4_sva_1),
      .all_same(leading_sign_57_0_1_0_21_out_2),
      .rtn(leading_sign_57_0_1_0_21_out_3)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_20_rg (
      .mantissa(z_out_9),
      .all_same(leading_sign_57_0_1_0_20_out_2),
      .rtn(leading_sign_57_0_1_0_20_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd55),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd55)) return_add_generic_AC_RND_CONV_false_20_lshift_rg (
      .a(55'b1111111111111111111111111111111111111111111111111111111),
      .s(return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1),
      .z(return_add_generic_AC_RND_CONV_false_20_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_25_rshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_25_rshift_rg_a[56:0]),
      .s(return_add_generic_AC_RND_CONV_false_25_e_dif_sat_sva_1),
      .z(return_add_generic_AC_RND_CONV_false_25_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd55),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd55)) return_add_generic_AC_RND_CONV_false_23_lshift_rg (
      .a(55'b1111111111111111111111111111111111111111111111111111111),
      .s(return_add_generic_AC_RND_CONV_false_23_e_dif_sat_sva_1),
      .z(return_add_generic_AC_RND_CONV_false_23_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_20_lshift_1_rg (
      .a(return_add_generic_AC_RND_CONV_false_15_res_mant_4_sva),
      .s(nl_return_add_generic_AC_RND_CONV_false_20_lshift_1_rg_s[5:0]),
      .z(return_add_generic_AC_RND_CONV_false_20_res_rounded_asn_rndc_sva_1)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_25_rg (
      .mantissa(z_out_5),
      .all_same(leading_sign_57_0_1_0_25_out_2),
      .rtn(leading_sign_57_0_1_0_25_out_3)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_24_rg (
      .mantissa(z_out_6),
      .all_same(leading_sign_57_0_1_0_24_out_2),
      .rtn(leading_sign_57_0_1_0_24_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd52),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd52)) return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_rg (
      .a(52'b1111111111111111111111111111111111111111111111111111),
      .s(nl_return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_rg_s[3:0]),
      .z(return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm)
    );
  leading_sign_53_0  leading_sign_53_0_6_rg (
      .mantissa(nl_leading_sign_53_0_6_rg_mantissa[52:0]),
      .rtn(leading_sign_53_0_6_out_1)
    );
  mgc_shift_l_v5 #(.width_a(32'sd55),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd55)) return_add_generic_AC_RND_CONV_false_19_lshift_1_rg (
      .a(55'b1111111111111111111111111111111111111111111111111111111),
      .s(return_add_generic_AC_RND_CONV_false_19_e_dif_sat_sva_1),
      .z(return_add_generic_AC_RND_CONV_false_19_lshift_1_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_13_rshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_13_rshift_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_13_rshift_rg_s[5:0]),
      .z(z_out_29)
    );
  mgc_shift_r_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_15_rshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_15_rshift_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_15_rshift_rg_s[5:0]),
      .z(z_out_30)
    );
  mgc_shift_r_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_10_rshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_s[5:0]),
      .z(z_out_31)
    );
  mgc_shift_r_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_11_rshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_11_rshift_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_11_rshift_rg_s[5:0]),
      .z(z_out_32)
    );
  mgc_shift_r_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_21_rshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_21_rshift_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_21_rshift_rg_s[5:0]),
      .z(z_out_33)
    );
  mgc_shift_r_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_17_rshift_1_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_17_rshift_1_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_17_rshift_1_rg_s[5:0]),
      .z(z_out_34)
    );
  mgc_shift_r_v5 #(.width_a(32'sd54),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd54)) return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg (
      .a(nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_a[53:0]),
      .s(nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_s[5:0]),
      .z(z_out_35)
    );
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_1_lshift_1_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_1_lshift_1_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_1_lshift_1_rg_s[5:0]),
      .z(z_out_36)
    );
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_21_lshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_21_lshift_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_21_lshift_rg_s[5:0]),
      .z(z_out_37)
    );
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_15_lshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_15_lshift_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_15_lshift_rg_s[5:0]),
      .z(z_out_38)
    );
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_10_lshift_1_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_s[5:0]),
      .z(z_out_39)
    );
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_13_lshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_13_lshift_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_13_lshift_rg_s[5:0]),
      .z(z_out_40)
    );
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_23_lshift_1_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_23_lshift_1_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_23_lshift_1_rg_s[5:0]),
      .z(z_out_41)
    );
  mgc_shift_l_v5 #(.width_a(32'sd55),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd55)) return_add_generic_AC_RND_CONV_false_17_lshift_1_rg (
      .a(55'b1111111111111111111111111111111111111111111111111111111),
      .s(nl_return_add_generic_AC_RND_CONV_false_17_lshift_1_rg_s[5:0]),
      .z(z_out_42)
    );
  mgc_shift_l_v5 #(.width_a(32'sd55),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd55)) return_add_generic_AC_RND_CONV_false_11_lshift_rg (
      .a(55'b1111111111111111111111111111111111111111111111111111111),
      .s(nl_return_add_generic_AC_RND_CONV_false_11_lshift_rg_s[5:0]),
      .z(z_out_43)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_11_rg (
      .mantissa(nl_leading_sign_57_0_1_0_11_rg_mantissa[56:0]),
      .all_same(all_same_out),
      .rtn(rtn_out)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_12_rg (
      .mantissa(z_out_8),
      .all_same(all_same_out_1),
      .rtn(rtn_out_1)
    );
  mgc_shift_l_v5 #(.width_a(32'sd106),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd106)) return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg (
      .a(nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_a[105:0]),
      .s(nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_s[5:0]),
      .z(z_out_54)
    );
  stage_run_ap_start_rsci stage_run_ap_start_rsci_inst (
      .ap_start_rsc_dat(ap_start_rsc_dat),
      .ap_start_rsc_vld(ap_start_rsc_vld),
      .ap_start_rsc_rdy(ap_start_rsc_rdy),
      .ap_start_rsci_oswt(reg_ap_start_rsci_iswt0_cse),
      .ap_start_rsci_wen_comp(ap_start_rsci_wen_comp)
    );
  stage_run_ap_done_rsci stage_run_ap_done_rsci_inst (
      .ap_done_rsc_dat(ap_done_rsc_dat),
      .ap_done_rsc_vld(ap_done_rsc_vld),
      .ap_done_rsc_rdy(ap_done_rsc_rdy),
      .ap_done_rsci_oswt(reg_out_u_triosy_obj_iswt0_cse),
      .ap_done_rsci_wen_comp(ap_done_rsci_wen_comp)
    );
  stage_run_wait_dp stage_run_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .in_f_d_rsci_en_d(in_f_d_rsci_en_d),
      .in_u_rsci_en_d(in_u_rsci_en_d),
      .out_f_d_rsci_en_d(out_f_d_rsci_en_d),
      .out_u_rsci_en_d(out_u_rsci_en_d),
      .BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en),
      .BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en(BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en),
      .BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en),
      .BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en(BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en),
      .r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en),
      .BUTTERFLY_i_div_cmp_z(BUTTERFLY_i_div_cmp_z),
      .run_wen(run_wen),
      .in_f_d_rsci_cgo(reg_in_f_d_rsci_cgo_ir_cse),
      .in_f_d_rsci_cgo_ir_unreg(or_673_rmff),
      .in_u_rsci_cgo(reg_in_u_rsci_cgo_ir_cse),
      .in_u_rsci_cgo_ir_unreg(or_672_rmff),
      .out_f_d_rsci_cgo(reg_out_f_d_rsci_cgo_ir_cse),
      .out_f_d_rsci_cgo_ir_unreg(or_671_rmff),
      .out_u_rsci_cgo(reg_out_u_rsci_cgo_ir_cse),
      .out_u_rsci_cgo_ir_unreg(or_670_rmff),
      .BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo),
      .BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo(BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo),
      .BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo),
      .BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo(BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo),
      .r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_cgo(reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_cgo_cse),
      .BUTTERFLY_i_div_cmp_z_oreg(BUTTERFLY_i_div_cmp_z_oreg)
    );
  stage_run_out1_rsci stage_run_out1_rsci_inst (
      .out1_rsc_dat(out1_rsc_dat),
      .out1_rsc_vld(out1_rsc_vld),
      .out1_rsc_rdy(out1_rsc_rdy),
      .out1_rsci_oswt(reg_out1_rsci_iswt0_cse),
      .out1_rsci_wen_comp(out1_rsci_wen_comp),
      .out1_rsci_idat(nl_stage_run_out1_rsci_inst_out1_rsci_idat[79:0])
    );
  stage_run_mode1_triosy_obj stage_run_mode1_triosy_obj_inst (
      .mode1_triosy_lz(mode1_triosy_lz),
      .run_wten(run_wten),
      .mode1_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_in_f_d_triosy_obj stage_run_in_f_d_triosy_obj_inst (
      .in_f_d_triosy_lz(in_f_d_triosy_lz),
      .run_wten(run_wten),
      .in_f_d_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_in_u_triosy_obj stage_run_in_u_triosy_obj_inst (
      .in_u_triosy_lz(in_u_triosy_lz),
      .run_wten(run_wten),
      .in_u_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_out_f_d_triosy_obj stage_run_out_f_d_triosy_obj_inst (
      .out_f_d_triosy_lz(out_f_d_triosy_lz),
      .run_wten(run_wten),
      .out_f_d_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_out_u_triosy_obj stage_run_out_u_triosy_obj_inst (
      .out_u_triosy_lz(out_u_triosy_lz),
      .run_wten(run_wten),
      .out_u_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_staller stage_run_staller_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .ap_start_rsci_wen_comp(ap_start_rsci_wen_comp),
      .ap_done_rsci_wen_comp(ap_done_rsci_wen_comp),
      .out1_rsci_wen_comp(out1_rsci_wen_comp)
    );
  stage_run_run_fsm stage_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .for_C_0_tr0(nl_stage_run_run_fsm_inst_for_C_0_tr0),
      .BUTTERFLY_C_15_tr0(nl_stage_run_run_fsm_inst_BUTTERFLY_C_15_tr0),
      .BUTTERFLY_C_15_tr1(and_dcpl_42),
      .BUTTERFLY_1_C_15_tr0(nl_stage_run_run_fsm_inst_BUTTERFLY_1_C_15_tr0),
      .BUTTERFLY_1_C_15_tr1(and_dcpl_44),
      .for_1_C_2_tr0(nl_stage_run_run_fsm_inst_for_1_C_2_tr0)
    );
  assign for_1_if_and_ssc = run_wen & (or_tmp_26 | out1_rsci_idat_63_0_mx0c1 | out1_rsci_idat_63_0_mx0c2);
  assign or_670_rmff = (stage_PE_1_and_cse & or_dcpl_87) | (~(mode_lpi_1_dfm | (~(or_dcpl_89
      | (fsm_output[6]) | or_dcpl_88)))) | (operator_16_false_operator_16_false_nor_cse_sva
      & or_dcpl_92) | (and_dcpl_35 & (fsm_output[26]));
  assign or_671_rmff = (mode_lpi_1_dfm & ((fsm_output[4]) | (fsm_output[30]) | (fsm_output[31])
      | (fsm_output[6]) | or_dcpl_88 | (fsm_output[8]))) | (stage_PE_1_and_1_tmp
      & (or_dcpl_99 | or_dcpl_98)) | (or_dcpl_101 & or_dcpl_92) | (and_dcpl_1 & (or_dcpl_102
      | (fsm_output[34])));
  assign or_672_rmff = (and_dcpl_35 & (or_dcpl_104 | (fsm_output[15]))) | and_421_cse
      | (stage_PE_1_and_cse & (or_dcpl_107 | or_dcpl_106)) | (~(mode_lpi_1_dfm |
      (~(or_dcpl_109 | (fsm_output[21]))))) | (and_dcpl_91 & (fsm_output[37]));
  assign or_673_rmff = (mode_lpi_1_dfm & ((fsm_output[20]) | (fsm_output[24]) | or_dcpl_87
      | or_dcpl_111 | (fsm_output[15]))) | (stage_PE_1_and_1_tmp & ((fsm_output[11])
      | (fsm_output[13]) | or_dcpl_106)) | and_421_cse | (and_dcpl_1 & ((fsm_output[18:16]!=3'b000)));
  assign BUTTERFLY_i_or_3_cse = (fsm_output[18]) | ((~ (fsm_output[2])) & or_tmp_46);
  assign BUTTERFLY_i_or_4_ssc = (or_tmp_180 & (~ or_tmp_46)) | (or_tmp_180 & or_tmp_46);
  assign BUTTERFLY_i_or_5_ssc = (or_tmp_181 & (~ or_tmp_46)) | (or_tmp_181 & or_tmp_46);
  assign BUTTERFLY_i_div_cmp_b = {reg_BUTTERFLY_i_div_cmp_b_ftd , reg_BUTTERFLY_i_div_cmp_b_1_ftd
      , reg_BUTTERFLY_i_div_cmp_b_1_ftd_4 , reg_BUTTERFLY_i_div_cmp_b_1_ftd_3 , reg_BUTTERFLY_i_div_cmp_b_1_ftd_1
      , reg_BUTTERFLY_i_div_cmp_b_ftd_2 , reg_BUTTERFLY_i_div_cmp_b_ftd_3 , reg_BUTTERFLY_i_div_cmp_b_ftd_4
      , reg_BUTTERFLY_i_div_cmp_b_ftd_5 , reg_BUTTERFLY_i_div_cmp_b_ftd_6_5 , reg_BUTTERFLY_i_div_cmp_b_ftd_6_4
      , reg_BUTTERFLY_i_div_cmp_b_ftd_6_3 , reg_BUTTERFLY_i_div_cmp_b_ftd_6_2 , reg_BUTTERFLY_i_div_cmp_b_ftd_6_1
      , reg_BUTTERFLY_i_div_cmp_b_ftd_6_0 , reg_BUTTERFLY_i_div_cmp_b_ftd_7};
  assign nor_155_cse = ~((fsm_output[34]) | (fsm_output[18]));
  assign BUTTERFLY_i_div_cmp_a = {7'b0, reg_BUTTERFLY_i_div_cmp_a_reg};
  assign BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr = reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_addr_cse;
  assign nl_BUTTERFLY_1_else_1_if_acc_1_sdt = (z_out_61[15:0]) + conv_u2s_14_16(signext_14_13({(z_out_61[17])
      , 11'b00000000000 , (z_out_61[17])}));
  assign BUTTERFLY_1_else_1_if_acc_1_sdt = nl_BUTTERFLY_1_else_1_if_acc_1_sdt[15:0];
  assign or_683_ssc = (fsm_output[22]) | (fsm_output[5]) | and_450_cse;
  assign or_685_ssc = (fsm_output[25]) | (fsm_output[35]) | and_448_cse;
  assign BUTTERFLY_if_1_or_1_cse = (fsm_output[26]) | (fsm_output[31]);
  assign BUTTERFLY_if_1_or_3_cse = (fsm_output[32:31]!=2'b00);
  assign or_709_ssc = or_dcpl_111 | (fsm_output[9]);
  assign or_710_ssc = (fsm_output[36]) | (fsm_output[12]) | (fsm_output[35]) | (fsm_output[15]);
  assign operator_16_false_and_cse = run_wen & (~(and_dcpl_110 & (~ (fsm_output[1]))));
  assign t_in_mux_4_nl = MUX_s_1_2_2(and_dcpl_42, and_dcpl_44, fsm_output[34]);
  assign t_in_and_cse = run_wen & ((~(t_in_mux_4_nl | and_dcpl_147)) | (fsm_output[1]));
  assign mode_or_cse = (fsm_output[18]) | (fsm_output[34]);
  assign mode_and_cse = run_wen & (~(and_dcpl_150 & and_dcpl_149));
  assign stage_PE_1_and_2_cse = run_wen & (~(and_dcpl_170 & (fsm_output[38:37]==2'b00)
      & and_dcpl_149));
  assign stage_PE_qif_qelse_mux_15_itm = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_5, t_in_10_0_lpi_1_dfm_1_4,
      mode_lpi_1_dfm);
  assign nor_90_cse = ~((fsm_output[17]) | (fsm_output[4]));
  assign operator_11_true_return_26_sva_2 = (in_f_d_rsci_q_d[62:52]==11'b11111111111);
  assign nl_operator_6_false_49_acc_sdt = conv_u2s_11_12({drf_qr_lval_10_smx_lpi_3_dfm_mx2_10
      , drf_qr_lval_10_smx_lpi_3_dfm_mx2_9_6 , drf_qr_lval_10_smx_lpi_3_dfm_mx2_5_0})
      + conv_s2s_7_12({1'b1 , (~ leading_sign_57_0_1_0_21_out_3)}) + 12'b000000000001;
  assign operator_6_false_49_acc_sdt = nl_operator_6_false_49_acc_sdt[11:0];
  assign nor_88_cse = ~((fsm_output[9:8]!=2'b00));
  assign nor_87_cse = ~((fsm_output[15:14]!=2'b00));
  assign nor_145_cse = ~((fsm_output[19]) | (fsm_output[6]));
  assign BUTTERFLY_1_i_and_ssc = run_wen & ((inverse_lpi_1_dfm_1 & (~(return_add_generic_AC_RND_CONV_false_15_res_mant_or_1_cse
      | or_dcpl_320 | or_dcpl_305 | (fsm_output[25]) | (fsm_output[6]) | or_dcpl_316
      | or_dcpl_82 | or_dcpl_300))) | or_dcpl_83 | BUTTERFLY_1_i_9_0_sva_mx0c3);
  assign return_add_generic_AC_RND_CONV_false_10_op1_mu_mux1h_3_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1,
      (stage_PE_1_x_im_d_sva[52]), and_dcpl_196);
  assign and_255_tmp = (~((~(return_add_generic_AC_RND_CONV_false_25_else_4_return_add_generic_AC_RND_CONV_false_25_else_4_nand_tmp
      & (~ (operator_33_true_50_acc_tmp[11])))) & return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11))
      & (~(return_add_generic_AC_RND_CONV_false_25_if_5_return_add_generic_AC_RND_CONV_false_25_if_5_and_tmp
      & (return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp[53]))) & and_dcpl_197
      & (~ leading_sign_57_0_1_0_25_out_2);
  assign return_add_generic_AC_RND_CONV_false_14_op1_mu_and_1_cse = (~ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp)
      & (fsm_output[25]);
  assign return_add_generic_AC_RND_CONV_false_14_op1_mu_and_2_cse = return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp
      & (fsm_output[25]);
  assign return_add_generic_AC_RND_CONV_false_14_op1_mu_and_cse = run_wen & (~ or_dcpl_338);
  assign return_add_generic_AC_RND_CONV_false_14_op1_mu_and_5_cse = (~ return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp)
      & (fsm_output[9]);
  assign return_add_generic_AC_RND_CONV_false_14_op1_mu_and_6_cse = return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp
      & (fsm_output[9]);
  assign return_add_generic_AC_RND_CONV_false_14_op1_mu_and_8_cse = return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_tmp
      & (fsm_output[10]);
  assign return_add_generic_AC_RND_CONV_false_14_op1_mu_and_7_cse = (~ return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_tmp)
      & (fsm_output[10]);
  assign return_add_generic_AC_RND_CONV_false_14_op1_mu_and_12_cse = return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp
      & (fsm_output[26]);
  assign return_add_generic_AC_RND_CONV_false_14_op1_mu_and_11_cse = (~ return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp)
      & (fsm_output[26]);
  assign and_258_tmp = or_dcpl_356 & inverse_lpi_1_dfm_1;
  assign and_261_tmp = or_dcpl_359 & inverse_lpi_1_dfm_1;
  assign and_264_tmp = or_dcpl_360 & inverse_lpi_1_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_10_and_3_m1c = and_258_tmp & (fsm_output[6]);
  assign return_add_generic_AC_RND_CONV_false_10_and_5_m1c = or_dcpl_357 & (fsm_output[13]);
  assign return_add_generic_AC_RND_CONV_false_10_and_7_m1c = or_dcpl_358 & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_10_and_9_m1c = and_261_tmp & (fsm_output[22]);
  assign return_add_generic_AC_RND_CONV_false_10_and_11_m1c = and_264_tmp & (fsm_output[24]);
  assign return_add_generic_AC_RND_CONV_false_10_and_13_m1c = or_dcpl_361 & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_10_and_4_cse = (~ or_dcpl_357) & (fsm_output[13]);
  assign return_add_generic_AC_RND_CONV_false_10_and_6_cse = (~ or_dcpl_358) & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_10_and_12_cse = (~ or_dcpl_361) & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_10_and_16_cse = (~ return_add_generic_AC_RND_CONV_false_11_op1_smaller_return_add_generic_AC_RND_CONV_false_11_op1_smaller_or_cse)
      & return_add_generic_AC_RND_CONV_false_10_and_5_m1c;
  assign return_add_generic_AC_RND_CONV_false_10_and_17_cse = return_add_generic_AC_RND_CONV_false_11_op1_smaller_return_add_generic_AC_RND_CONV_false_11_op1_smaller_or_cse
      & return_add_generic_AC_RND_CONV_false_10_and_5_m1c;
  assign return_add_generic_AC_RND_CONV_false_10_and_18_cse = (~ return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse)
      & return_add_generic_AC_RND_CONV_false_10_and_7_m1c;
  assign return_add_generic_AC_RND_CONV_false_10_and_19_cse = return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse
      & return_add_generic_AC_RND_CONV_false_10_and_7_m1c;
  assign return_add_generic_AC_RND_CONV_false_10_and_24_cse = (~ return_add_generic_AC_RND_CONV_false_24_op1_smaller_return_add_generic_AC_RND_CONV_false_24_op1_smaller_or_cse)
      & return_add_generic_AC_RND_CONV_false_10_and_13_m1c;
  assign return_add_generic_AC_RND_CONV_false_10_and_25_cse = return_add_generic_AC_RND_CONV_false_24_op1_smaller_return_add_generic_AC_RND_CONV_false_24_op1_smaller_or_cse
      & return_add_generic_AC_RND_CONV_false_10_and_13_m1c;
  assign BUTTERFLY_and_ssc = run_wen & (fsm_output[9:7]==3'b000);
  assign return_add_generic_AC_RND_CONV_false_17_and_3_cse = return_add_generic_AC_RND_CONV_false_12_do_sub_sva
      & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_17_and_7_cse = (~ return_add_generic_AC_RND_CONV_false_4_do_sub_sva_1)
      & (fsm_output[22]);
  assign return_add_generic_AC_RND_CONV_false_17_and_8_cse = return_add_generic_AC_RND_CONV_false_4_do_sub_sva_1
      & (fsm_output[22]);
  assign return_add_generic_AC_RND_CONV_false_17_and_9_cse = (~ return_add_generic_AC_RND_CONV_false_12_do_sub_sva)
      & (fsm_output[29]);
  assign nl_BUTTERFLY_1_else_3_else_acc_4_sdt = (stage_u_add_9_acc_psp_sva_1[15:0])
      + conv_u2u_14_16(signext_14_13({(stage_u_add_9_acc_psp_sva_1[17]) , 11'b00000000000
      , (stage_u_add_9_acc_psp_sva_1[17])}));
  assign BUTTERFLY_1_else_3_else_acc_4_sdt = nl_BUTTERFLY_1_else_3_else_acc_4_sdt[15:0];
  assign BUTTERFLY_1_else_1_if_nor_cse = ~((fsm_output[11]) | (fsm_output[10]) |
      (fsm_output[8]));
  assign BUTTERFLY_1_else_1_if_and_ssc = run_wen & ((mode_lpi_1_dfm & BUTTERFLY_1_else_1_if_nor_cse)
      | BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c0 | BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c4
      | (fsm_output[22]) | (fsm_output[24]) | BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c7
      | (fsm_output[28]));
  assign BUTTERFLY_else_1_if_or_3_cse = (fsm_output[12]) | (fsm_output[28]);
  assign BUTTERFLY_else_1_if_and_cse = inverse_lpi_1_dfm_1 & (fsm_output[9]) & BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c7;
  assign BUTTERFLY_else_1_if_and_1_cse = (~ inverse_lpi_1_dfm_1) & BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c7;
  assign and_2638_cse = mode_lpi_1_dfm & (fsm_output[9]);
  assign nl_operator_33_true_37_acc_nl = (operator_6_false_40_acc_psp_1_sva_1[10:1])
      + 10'b0000000001;
  assign operator_33_true_37_acc_nl = nl_operator_33_true_37_acc_nl[9:0];
  assign and_1161_nl = (return_add_generic_AC_RND_CONV_false_18_res_rounded_acc_tmp[53])
      & (fsm_output[23]) & (~ or_1477_tmp);
  assign and_1163_nl = (~ (return_add_generic_AC_RND_CONV_false_18_res_rounded_acc_tmp[53]))
      & (fsm_output[23]) & (~ or_1477_tmp);
  assign and_1169_nl = (return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp[53])
      & (fsm_output[30]);
  assign and_1171_nl = (~ (return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp[53]))
      & (fsm_output[30]) & (~ or_1477_tmp);
  assign mux1h_3_nl = MUX1HOT_v_10_10_2((r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[61:52]),
      (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[61:52]), return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1,
      (stage_PE_1_x_re_d_sva[62:53]), operator_33_true_37_acc_nl, (operator_33_true_36_acc_psp_1_sva_1[10:1]),
      return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_mx1w0, (stage_PE_1_x_im_d_sva[62:53]),
      (return_add_generic_AC_RND_CONV_false_25_exp_plus_1_12_1_lpi_3_dfm_1[9:0]),
      (operator_33_true_50_acc_tmp[10:1]), {or_tmp_388 , or_tmp_389 , and_1132_ssc
      , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse , and_1161_nl
      , and_1163_nl , and_1813_cse , and_1808_cse , and_1169_nl , and_1171_nl});
  assign not_734_nl = ~ or_1477_tmp;
  assign and_2143_itm = MUX_v_10_2_2(10'b0000000000, mux1h_3_nl, not_734_nl);
  assign or_965_itm = (fsm_output[13]) | (fsm_output[23]) | (fsm_output[14]) | BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c4;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse = (fsm_output[6])
      | (fsm_output[22]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_cse = run_wen & (~(or_dcpl_437
      | or_dcpl_436));
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_4_cse = (~ and_dcpl_225)
      & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_5_cse = and_dcpl_225
      & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse = (~ and_dcpl_226)
      & (fsm_output[13]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse = and_dcpl_228
      & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse = (~ and_dcpl_227)
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse = (~ and_dcpl_228)
      & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_11_cse = and_dcpl_227
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse = and_dcpl_226
      & (fsm_output[13]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse = (~ return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp)
      & (fsm_output[24]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_13_cse = return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp
      & (fsm_output[24]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_cse = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_11_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_1_cse = run_wen &
      (~ (fsm_output[15]));
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_18_cse = (~ return_extract_12_return_extract_12_or_1_tmp)
      & (fsm_output[9]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_5_cse = (return_extract_12_return_extract_12_or_1_tmp
      & (fsm_output[9])) | (return_extract_44_return_extract_44_or_1_tmp & (fsm_output[25]));
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_24_cse = (~ return_extract_44_return_extract_44_or_1_tmp)
      & (fsm_output[25]);
  assign return_extract_41_and_cse = run_wen & (~((fsm_output[26]) | (fsm_output[24])
      | or_dcpl_443 | or_dcpl_442));
  assign return_extract_41_and_1_cse = return_extract_41_and_cse & mode_lpi_1_dfm;
  assign return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_2_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_226);
  assign return_add_generic_AC_RND_CONV_false_14_op1_mu_mux_1_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm, and_dcpl_227);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_cse = (~ return_add_generic_AC_RND_CONV_false_5_do_sub_sva_1)
      & (fsm_output[22]);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse = return_add_generic_AC_RND_CONV_false_5_do_sub_sva_1
      & (fsm_output[22]);
  assign return_add_generic_AC_RND_CONV_false_4_op_bigger_mux_3_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_4_op1_mu_52_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_4_op2_mu_52_lpi_3_dfm_mx0, and_dcpl_225);
  assign return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_cse = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[50]),
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0, and_dcpl_226);
  assign return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_cse = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0[50]),
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50, and_dcpl_227);
  assign nl_return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_acc_1_nl = ({1'b1
      , (stage_PE_1_x_im_d_sva[51:0])}) + conv_u2u_52_53({(~ return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm_mx2)
      , (~ return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_mx0w6)}) +
      53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_acc_1_nl = nl_return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_acc_1_nl[52:0];
  assign return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_and_cse
      = (readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_acc_1_nl))
      & return_add_generic_AC_RND_CONV_false_23_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_25_op1_smaller_return_add_generic_AC_RND_CONV_false_25_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_23_e_dif1_acc_1_tmp[11]);
  assign return_add_generic_AC_RND_CONV_false_11_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_11_op1_smaller_oelse_and_cse
      = z_out_2_52 & return_add_generic_AC_RND_CONV_false_9_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_11_op1_smaller_return_add_generic_AC_RND_CONV_false_11_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_11_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_11_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_9_e_dif1_acc_1_tmp[11]);
  assign return_add_generic_AC_RND_CONV_false_11_and_26_m1c = or_dcpl_356 & (fsm_output[6]);
  assign return_add_generic_AC_RND_CONV_false_11_and_28_m1c = or_dcpl_488 & (fsm_output[8]);
  assign return_add_generic_AC_RND_CONV_false_11_and_32_m1c = or_dcpl_359 & (fsm_output[22]);
  assign return_add_generic_AC_RND_CONV_false_11_and_34_m1c = or_dcpl_480 & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_11_and_27_cse = (~ or_dcpl_488) & (fsm_output[8]);
  assign return_add_generic_AC_RND_CONV_false_11_and_37_cse = (~ or_446_cse) & return_add_generic_AC_RND_CONV_false_11_and_28_m1c;
  assign return_add_generic_AC_RND_CONV_false_11_and_38_cse = or_446_cse & return_add_generic_AC_RND_CONV_false_11_and_28_m1c;
  assign return_add_generic_AC_RND_CONV_false_24_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_24_op1_smaller_oelse_and_cse
      = z_out_2_52 & return_add_generic_AC_RND_CONV_false_22_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_24_op1_smaller_return_add_generic_AC_RND_CONV_false_24_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_24_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_24_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_22_e_dif1_acc_1_tmp[11]);
  assign nl_return_add_generic_AC_RND_CONV_false_10_ma1_lt_ma2_acc_1_nl = ({1'b1
      , (stage_PE_1_x_im_d_sva[51:0])}) + conv_u2u_52_53({(~ return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm)
      , (~ return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0)}) + 53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_10_ma1_lt_ma2_acc_1_nl = nl_return_add_generic_AC_RND_CONV_false_10_ma1_lt_ma2_acc_1_nl[52:0];
  assign return_add_generic_AC_RND_CONV_false_10_ma1_lt_ma2_acc_1_itm_52 = readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_10_ma1_lt_ma2_acc_1_nl);
  assign return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_and_cse
      = return_add_generic_AC_RND_CONV_false_10_ma1_lt_ma2_acc_1_itm_52 & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva;
  assign return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_10_e_dif1_acc_1_tmp[11]);
  assign return_add_generic_AC_RND_CONV_false_12_and_6_m1c = or_dcpl_360 & (fsm_output[24]);
  assign return_extract_15_m_zero_mux1h_3_cse = ~((in_f_d_rsci_q_d[51:0]!=52'b0000000000000000000000000000000000000000000000000000));
  assign return_add_generic_AC_RND_CONV_false_11_mux_19_cse = MUX_s_1_2_2((stage_PE_1_tmp_im_d_1_sva_1_63_51[12]),
      return_add_generic_AC_RND_CONV_false_11_mux_itm, inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_5_e_dif_sat_or_2_nl = (return_add_generic_AC_RND_CONV_false_4_e_dif_qif_acc_pmx_lpi_3_dfm_mx0_9_0[9:6]!=4'b0000)
      | ((return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt[10]) & (return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp[10]));
  assign return_add_generic_AC_RND_CONV_false_4_e_dif_sat_or_cse = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_4_e_dif_qif_acc_pmx_lpi_3_dfm_mx0_9_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_5_e_dif_sat_or_2_nl);
  assign return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_3_itm = MUX_v_6_2_2((drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_0[5:0]),
      leading_sign_57_0_1_0_6_out_3, return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_10_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_5_itm = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_10_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_9_itm = MUX_v_6_2_2((drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_0[5:0]),
      leading_sign_57_0_1_0_19_out_3, return_add_generic_AC_RND_CONV_false_19_acc_2_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_14_and_cse = run_wen & (~(or_dcpl_320
      | (fsm_output[11]) | or_dcpl_511));
  assign return_add_generic_AC_RND_CONV_false_14_or_cse = (fsm_output[7]) | (fsm_output[23]);
  assign return_add_generic_AC_RND_CONV_false_3_op_bigger_mux_1_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_1_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_3_op_bigger_mux_2_cse = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0,
      return_add_generic_AC_RND_CONV_false_1_op2_mu_51_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_1_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_op_bigger_mux_1_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm, or_446_cse);
  assign return_add_generic_AC_RND_CONV_false_op_bigger_mux_2_cse = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_1_op2_mu_51_1_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0, or_446_cse);
  assign return_add_generic_AC_RND_CONV_false_16_op_bigger_mux_1_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm_1, or_452_cse);
  assign return_add_generic_AC_RND_CONV_false_16_op_bigger_mux_2_cse = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0,
      return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm_mx1, or_452_cse);
  assign return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_1_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm, or_445_cse);
  assign return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_cse = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm_mx1,
      return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0, or_445_cse);
  assign return_add_generic_AC_RND_CONV_false_15_res_mant_or_1_cse = (fsm_output[26])
      | (fsm_output[28]);
  assign return_add_generic_AC_RND_CONV_false_15_res_mant_or_cse = (fsm_output[6])
      | (fsm_output[8]) | (fsm_output[22]) | (fsm_output[24]);
  assign or_1143_itm = or_dcpl_338 | (fsm_output[9]);
  assign stage_PE_1_tmp_im_d_and_ssc = run_wen & (~((fsm_output[24]) | (fsm_output[8])));
  assign and_1132_ssc = return_add_generic_AC_RND_CONV_false_11_op1_smaller_return_add_generic_AC_RND_CONV_false_11_op1_smaller_or_cse
      & (fsm_output[13]);
  assign and_1141_ssc = (return_add_generic_AC_RND_CONV_false_17_res_rounded_acc_tmp[53])
      & (fsm_output[23]);
  assign and_1143_ssc = (~ (return_add_generic_AC_RND_CONV_false_17_res_rounded_acc_tmp[53]))
      & (fsm_output[23]);
  assign and_1145_ssc = return_add_generic_AC_RND_CONV_false_24_op1_smaller_return_add_generic_AC_RND_CONV_false_24_op1_smaller_or_cse
      & (fsm_output[29]);
  assign and_1149_ssc = (~ (return_add_generic_AC_RND_CONV_false_24_res_rounded_acc_tmp[53]))
      & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_7_exp_and_ssc = run_wen & (~(or_dcpl_99
      | or_dcpl_523));
  assign and_2120_cse = return_add_generic_AC_RND_CONV_false_17_op1_smaller_lor_lpi_3_dfm_2
      & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  assign and_1134_cse = and_dcpl_241 & (fsm_output[29]);
  assign and_2123_cse = and_1134_cse | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse;
  assign and_2126_cse = and_1141_ssc & (~ or_dcpl_629);
  assign and_2127_cse = and_1143_ssc & (~ or_dcpl_629);
  assign and_2129_cse = (return_add_generic_AC_RND_CONV_false_24_res_rounded_acc_tmp[53])
      & (fsm_output[30]);
  assign and_2130_cse = and_1149_ssc & (~ or_dcpl_629);
  assign BUTTERFLY_else_2_and_ssc = run_wen & (~ or_dcpl_471);
  assign or_954_rgt = and_1014_cse | (and_dcpl_214 & (fsm_output[8]));
  assign or_955_rgt = (and_dcpl_215 & (fsm_output[22])) | (and_dcpl_216 & (fsm_output[6]));
  assign or_959_rgt = and_1029_cse | (or_451_cse & (fsm_output[12]));
  assign or_960_rgt = and_1032_cse | (and_dcpl_224 & (fsm_output[24]));
  assign BUTTERFLY_else_2_and_2_rgt = (~ mode_lpi_1_dfm) & (fsm_output[12]);
  assign nor_99_ssc = ~(inverse_lpi_1_dfm_1 | return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_18_and_4_cse = nor_99_ssc & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_18_and_8_cse = inverse_lpi_1_dfm_1
      & (fsm_output[29]);
  assign and_1813_cse = return_add_generic_AC_RND_CONV_false_25_op1_smaller_return_add_generic_AC_RND_CONV_false_25_op1_smaller_or_cse
      & (fsm_output[29]);
  assign and_1808_cse = and_dcpl_196 & (fsm_output[29]);
  assign and_1804_cse = return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse
      & (fsm_output[14]);
  assign nl_operator_32_false_acc_nl = (~ (z_out_25[3:0])) + ({(z_out_25[1:0]) ,
      2'b01});
  assign operator_32_false_acc_nl = nl_operator_32_false_acc_nl[3:0];
  assign nl_in_u_mux1h_1_itm = ({operator_32_false_acc_nl , 12'b000000000001}) +
      (~ (z_out_25[15:0]));
  assign in_u_mux1h_1_itm = nl_in_u_mux1h_1_itm[15:0];
  assign return_add_generic_AC_RND_CONV_false_14_op1_mu_and_13_cse = (~ and_dcpl_196)
      & (fsm_output[29]);
  assign BUTTERFLY_1_fiy_and_4_cse = return_add_generic_AC_RND_CONV_false_24_op1_smaller_return_add_generic_AC_RND_CONV_false_24_op1_smaller_or_cse
      & (~ inverse_lpi_1_dfm_1) & (fsm_output[29]);
  assign BUTTERFLY_1_fiy_and_5_cse = or_dcpl_441 & (~((return_add_generic_AC_RND_CONV_false_22_e_dif1_acc_1_tmp[11])
      | inverse_lpi_1_dfm_1)) & (fsm_output[29]);
  assign and_336_cse = and_dcpl_281 & and_dcpl_254 & (~ leading_sign_57_0_1_0_2_out_2);
  assign return_add_generic_AC_RND_CONV_false_9_exp_mux1h_2_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1,
      (stage_PE_1_x_re_d_sva[52]), and_dcpl_226);
  assign and_342_tmp = (~((~(return_add_generic_AC_RND_CONV_false_23_else_4_return_add_generic_AC_RND_CONV_false_23_else_4_nand_tmp
      & (~ (operator_33_true_46_acc_tmp[11])))) & return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1))
      & (~(return_add_generic_AC_RND_CONV_false_23_if_5_return_add_generic_AC_RND_CONV_false_23_if_5_and_tmp
      & (return_add_generic_AC_RND_CONV_false_23_res_rounded_acc_tmp[53]))) & and_dcpl_197
      & (~ leading_sign_57_0_1_0_15_out_2);
  assign stage_PE_1_tmp_im_d_and_6_cse = inverse_lpi_1_dfm_1 & (fsm_output[23]);
  assign return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse = (fsm_output[12])
      | (fsm_output[16]);
  assign or_1266_cse = (fsm_output[24]) | (fsm_output[22]);
  assign return_add_generic_AC_RND_CONV_false_20_ls_or_cse = (fsm_output[7]) | (fsm_output[14]);
  assign operator_6_false_18_or_cse = (fsm_output[12]) | (fsm_output[26]) | (fsm_output[28]);
  assign and_1585_rgt = inverse_lpi_1_dfm_1 & (fsm_output[7]);
  assign and_1587_rgt = (~ inverse_lpi_1_dfm_1) & return_add_generic_AC_RND_CONV_false_14_or_cse;
  assign stage_PE_tmp_im_d_mux1h_nl = MUX1HOT_v_10_6_2(stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1,
      (stage_PE_1_tmp_im_d_1_sva_1_63_51[11:2]), (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_1[10:1]),
      (z_out_24[10:1]), stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w4_10_1, (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_1[10:1]),
      {and_1585_rgt , and_1587_rgt , stage_PE_tmp_im_d_and_cse , stage_PE_tmp_im_d_or_cse
      , stage_PE_1_tmp_im_d_and_6_cse , stage_PE_tmp_im_d_and_2_cse});
  assign not_726_nl = ~ or_tmp_830;
  assign operator_6_false_18_mux1h_itm_10_1 = MUX_v_10_2_2(10'b0000000000, stage_PE_tmp_im_d_mux1h_nl,
      not_726_nl);
  assign or_1285_itm = or_dcpl_320 | or_dcpl_523 | or_dcpl_442;
  assign return_extract_15_and_3_cse = run_wen & (~ return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_2_cse);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_mux_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0, and_dcpl_226);
  assign return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_1_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm, and_dcpl_227);
  assign and_352_tmp = (~((~((~ (operator_33_true_48_acc_tmp[11])) & return_add_generic_AC_RND_CONV_false_24_else_4_return_add_generic_AC_RND_CONV_false_24_else_4_nand_tmp))
      & return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11)) & (~(return_add_generic_AC_RND_CONV_false_24_if_5_return_add_generic_AC_RND_CONV_false_24_if_5_and_tmp
      & (return_add_generic_AC_RND_CONV_false_24_res_rounded_acc_tmp[53]))) & and_dcpl_294
      & (~ leading_sign_57_0_1_0_24_out_2);
  assign return_add_generic_AC_RND_CONV_false_11_exp_and_1_cse = (~ return_add_generic_AC_RND_CONV_false_21_unequal_tmp)
      & (fsm_output[10]);
  assign return_add_generic_AC_RND_CONV_false_11_exp_and_2_cse = return_add_generic_AC_RND_CONV_false_21_unequal_tmp
      & (fsm_output[10]);
  assign return_add_generic_AC_RND_CONV_false_17_m_r_and_cse = run_wen & (~(or_dcpl_89
      | (fsm_output[9])));
  assign return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_2_cse = (fsm_output[9])
      | (fsm_output[25]);
  assign nl_stage_u_add_3_mux1h_2_itm = conv_u2s_16_17(z_out_64_31_16) + 17'b11100111111111111;
  assign stage_u_add_3_mux1h_2_itm = nl_stage_u_add_3_mux1h_2_itm[16:0];
  assign or_1367_cse = (fsm_output[22:21]!=2'b00);
  assign BUTTERFLY_1_if_mux_itm = MUX_v_14_2_2(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out,
      BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out, inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1 = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[49:0]),
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_226);
  assign return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0[49:0]),
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0, and_dcpl_227);
  assign nl_return_mult_generic_AC_RND_CONV_false_2_if_acc_1_nl =  -operator_6_false_16_acc_psp_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_2_if_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_2_if_acc_1_nl[12:0];
  assign return_mult_generic_AC_RND_CONV_false_2_if_acc_1_itm_12_1 = readslicef_13_1_12(return_mult_generic_AC_RND_CONV_false_2_if_acc_1_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_1_if_acc_1_nl =  -z_out_57;
  assign return_mult_generic_AC_RND_CONV_false_1_if_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_1_if_acc_1_nl[12:0];
  assign return_mult_generic_AC_RND_CONV_false_1_if_acc_1_itm_12_1 = readslicef_13_1_12(return_mult_generic_AC_RND_CONV_false_1_if_acc_1_nl);
  assign return_add_generic_AC_RND_CONV_false_1_if_5_or_2_nl = return_add_generic_AC_RND_CONV_false_2_acc_3_itm_11_1
      | (~((operator_33_true_4_acc_tmp!=13'b0000000000000)));
  assign return_add_generic_AC_RND_CONV_false_1_mux_29_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_2_acc_3_itm_11_1,
      return_add_generic_AC_RND_CONV_false_1_if_5_or_2_nl, return_add_generic_AC_RND_CONV_false_2_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0 = leading_sign_57_0_1_0_2_out_2
      | (~ return_add_generic_AC_RND_CONV_false_1_mux_29_nl);
  assign return_add_generic_AC_RND_CONV_false_2_else_4_return_add_generic_AC_RND_CONV_false_2_else_4_nand_tmp
      = ~((operator_33_true_4_acc_tmp[11:0]==12'b011111111111));
  assign return_add_generic_AC_RND_CONV_false_3_if_5_or_2_nl = return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1
      | (~((z_out_13!=13'b0000000000000)));
  assign return_add_generic_AC_RND_CONV_false_3_mux_23_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1,
      return_add_generic_AC_RND_CONV_false_3_if_5_or_2_nl, return_add_generic_AC_RND_CONV_false_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w0 = leading_sign_57_0_1_0_15_out_2
      | (~ return_add_generic_AC_RND_CONV_false_3_mux_23_nl);
  assign return_add_generic_AC_RND_CONV_false_15_else_4_return_add_generic_AC_RND_CONV_false_15_else_4_nand_tmp
      = ~((z_out_13[11:0]==12'b011111111111));
  assign return_add_generic_AC_RND_CONV_false_6_mux_32_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva,
      return_add_generic_AC_RND_CONV_false_6_if_5_or_3, return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1 = return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_6_mux_32_nl);
  assign return_add_generic_AC_RND_CONV_false_7_mux_17_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1,
      return_add_generic_AC_RND_CONV_false_7_if_5_or_3, return_add_generic_AC_RND_CONV_false_7_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs_mx0w0 = return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_7_mux_17_nl);
  assign return_add_generic_AC_RND_CONV_false_10_else_4_return_add_generic_AC_RND_CONV_false_10_else_4_nand_tmp
      = ~((stage_u_add_3_acc_itm_rsp_1[11:0]==12'b011111111111));
  assign return_add_generic_AC_RND_CONV_false_8_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1,
      return_add_generic_AC_RND_CONV_false_8_if_5_or_3, z_out_46[53]);
  assign return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs_mx0w0 = return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_8_mux_13_nl);
  assign return_add_generic_AC_RND_CONV_false_21_else_4_return_add_generic_AC_RND_CONV_false_21_else_4_nand_tmp
      = ~(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0 & (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0==9'b111111111)
      & reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1 & (~ (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_2_1[0])));
  assign nl_return_mult_generic_AC_RND_CONV_false_5_if_acc_1_nl =  -operator_6_false_45_acc_psp_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_5_if_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_5_if_acc_1_nl[12:0];
  assign return_mult_generic_AC_RND_CONV_false_5_if_acc_1_itm_12_1 = readslicef_13_1_12(return_mult_generic_AC_RND_CONV_false_5_if_acc_1_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_4_if_acc_1_nl =  -z_out_63;
  assign return_mult_generic_AC_RND_CONV_false_4_if_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_4_if_acc_1_nl[12:0];
  assign return_mult_generic_AC_RND_CONV_false_4_if_acc_1_itm_12_1 = readslicef_13_1_12(return_mult_generic_AC_RND_CONV_false_4_if_acc_1_nl);
  assign return_add_generic_AC_RND_CONV_false_20_mux_17_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1,
      return_add_generic_AC_RND_CONV_false_7_if_5_or_3, return_add_generic_AC_RND_CONV_false_20_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs_mx0w0 = return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_20_mux_17_nl);
  assign return_add_generic_AC_RND_CONV_false_21_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1,
      return_add_generic_AC_RND_CONV_false_8_if_5_or_3, return_add_generic_AC_RND_CONV_false_21_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs_mx0w0 = return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_21_mux_13_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl =  -operator_6_false_58_acc_psp_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl[11:0];
  assign return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1 = readslicef_12_1_11(return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl);
  assign return_add_generic_AC_RND_CONV_false_9_if_5_or_2_nl = return_add_generic_AC_RND_CONV_false_22_acc_3_itm_11_1
      | (~((operator_33_true_44_acc_tmp!=13'b0000000000000)));
  assign return_add_generic_AC_RND_CONV_false_9_mux_32_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_22_acc_3_itm_11_1,
      return_add_generic_AC_RND_CONV_false_9_if_5_or_2_nl, z_out_47[53]);
  assign return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs_mx0w0 = leading_sign_57_0_1_0_2_out_2
      | (~ return_add_generic_AC_RND_CONV_false_9_mux_32_nl);
  assign return_add_generic_AC_RND_CONV_false_10_mux_16_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1,
      return_add_generic_AC_RND_CONV_false_7_if_5_or_3, z_out_46[53]);
  assign return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs_mx0w0 = return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_10_mux_16_nl);
  assign return_add_generic_AC_RND_CONV_false_11_mux_9_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva,
      return_add_generic_AC_RND_CONV_false_6_if_5_or_3, z_out_46[53]);
  assign return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w0 = return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_11_mux_9_nl);
  assign return_add_generic_AC_RND_CONV_false_24_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11
      | (~((operator_33_true_48_acc_tmp!=13'b0000000000000)));
  assign return_add_generic_AC_RND_CONV_false_24_mux_9_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11,
      return_add_generic_AC_RND_CONV_false_24_if_5_or_1_nl, return_add_generic_AC_RND_CONV_false_24_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs_mx0w0 = leading_sign_57_0_1_0_24_out_2
      | (~ return_add_generic_AC_RND_CONV_false_24_mux_9_nl);
  assign return_add_generic_AC_RND_CONV_false_25_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11
      | (~((operator_33_true_50_acc_tmp!=13'b0000000000000)));
  assign return_add_generic_AC_RND_CONV_false_25_mux_9_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11,
      return_add_generic_AC_RND_CONV_false_25_if_5_or_1_nl, return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs_mx0w0 = leading_sign_57_0_1_0_25_out_2
      | (~ return_add_generic_AC_RND_CONV_false_25_mux_9_nl);
  assign return_add_generic_AC_RND_CONV_false_23_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1
      | (~((operator_33_true_46_acc_tmp!=13'b0000000000000)));
  assign return_add_generic_AC_RND_CONV_false_23_mux_16_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1,
      return_add_generic_AC_RND_CONV_false_23_if_5_or_1_nl, return_add_generic_AC_RND_CONV_false_23_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs_mx0w0 = leading_sign_57_0_1_0_15_out_2
      | (~ return_add_generic_AC_RND_CONV_false_23_mux_16_nl);
  assign return_add_generic_AC_RND_CONV_false_23_else_4_return_add_generic_AC_RND_CONV_false_23_else_4_nand_tmp
      = ~((operator_33_true_46_acc_tmp[11:0]==12'b011111111111));
  assign return_add_generic_AC_RND_CONV_false_24_else_4_return_add_generic_AC_RND_CONV_false_24_else_4_nand_tmp
      = ~((operator_33_true_48_acc_tmp[11:0]==12'b011111111111));
  assign return_add_generic_AC_RND_CONV_false_25_else_4_return_add_generic_AC_RND_CONV_false_25_else_4_nand_tmp
      = ~((operator_33_true_50_acc_tmp[11:0]==12'b011111111111));
  assign operator_16_false_1_operator_16_false_1_and_mdf_sva_1 = (mode1_rsci_idat==16'b0000000000000001);
  assign operator_16_false_operator_16_false_nor_tmp = ~((mode1_rsci_idat!=16'b0000000000000000));
  assign mode_lpi_1_dfm_mx0w0 = operator_16_false_1_operator_16_false_1_and_mdf_sva_1
      | operator_16_false_operator_16_false_nor_tmp;
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_8 = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_1,
      t_in_10_0_lpi_1_dfm_1_0, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_7 = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_2,
      t_in_10_0_lpi_1_dfm_1_1, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_6 = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_3,
      t_in_10_0_lpi_1_dfm_1_2, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_5 = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_4,
      t_in_10_0_lpi_1_dfm_1_3, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_2 = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_7,
      t_in_10_0_lpi_1_dfm_1_6, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_1 = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_8,
      t_in_10_0_lpi_1_dfm_1_7, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_0 = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_9,
      t_in_10_0_lpi_1_dfm_1_8, mode_lpi_1_dfm);
  assign stage_PE_1_and_1_tmp = mode_lpi_1_dfm & inverse_lpi_1_dfm_1;
  assign stage_PE_asn_13_mx0w0 = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_10, t_in_10_0_lpi_1_dfm_1_9,
      mode_lpi_1_dfm);
  assign stage_PE_index_const_15_lpi_2_dfm_mx0w0 = m_in_15_1_lpi_1_dfm_1_rsp_0_13
      & (~ mode_lpi_1_dfm) & inverse_lpi_1_dfm_1;
  assign stage_PE_qif_qelse_mux_11_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_0, m_in_15_1_lpi_1_dfm_1_rsp_0_9,
      mode_lpi_1_dfm);
  assign stage_PE_index_const_10_lpi_2_dfm_mx0w0 = stage_PE_qif_qelse_mux_11_nl &
      inverse_lpi_1_dfm_1;
  assign stage_PE_1_and_cse = (~ mode_lpi_1_dfm) & inverse_lpi_1_dfm_1;
  assign operator_11_true_return_3_sva_mx1w0 = (out_f_d_rsci_q_d[62:52]==11'b11111111111);
  assign nl_BUTTERFLY_i_9_0_sva_1 = conv_u2u_9_10(operator_6_false_49_acc_psp_sva_8_0)
      + (z_out_26[9:0]);
  assign BUTTERFLY_i_9_0_sva_1 = nl_BUTTERFLY_i_9_0_sva_1[9:0];
  assign return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp
      = (out_f_d_rsci_q_d[62:52]!=11'b00000000000);
  assign return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1 = (out_f_d_rsci_q_d[51])
      | return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1 = (stage_PE_1_x_im_d_sva[0])
      & return_add_generic_AC_RND_CONV_false_10_mux_7_itm;
  assign return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm_1 = (in_f_d_rsci_q_d[51])
      | return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_10_if_2_return_add_generic_AC_RND_CONV_false_10_if_2_and_1_mx3w0
      = operator_11_true_return_15_sva & (stage_PE_1_x_im_d_sva[63]);
  assign return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp
      = (in_f_d_rsci_q_d[62:52]!=11'b00000000000);
  assign return_extract_3_m_zero_sva_1 = ~((out_f_d_rsci_q_d[51:0]!=52'b0000000000000000000000000000000000000000000000000000));
  assign return_extract_17_m_zero_sva_mx0w3 = ~(BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx1
      | (return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_add_generic_AC_RND_CONV_false_18_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_18_acc_2_itm_10
      | (~((operator_33_true_36_acc_psp_1_sva_1!=12'b000000000000)));
  assign return_add_generic_AC_RND_CONV_false_18_mux_9_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_18_acc_2_itm_10,
      return_add_generic_AC_RND_CONV_false_18_if_5_or_1_nl, return_add_generic_AC_RND_CONV_false_18_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_svs_1 = leading_sign_57_0_1_0_18_out_2
      | (~ return_add_generic_AC_RND_CONV_false_18_mux_9_nl);
  assign return_add_generic_AC_RND_CONV_false_9_op1_inf_sva_1 = operator_11_true_return_24_sva
      & return_extract_1_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_1_else_2_else_else_mux_nl = MUX_v_11_2_2((return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_1[10:0]),
      (z_out_55[10:0]), return_mult_generic_AC_RND_CONV_false_1_e_incr_lpi_3_dfm_2);
  assign return_mult_generic_AC_RND_CONV_false_1_else_2_else_return_mult_generic_AC_RND_CONV_false_1_else_2_else_and_nl
      = MUX_v_11_2_2(11'b00000000000, return_mult_generic_AC_RND_CONV_false_1_else_2_else_else_mux_nl,
      return_mult_generic_AC_RND_CONV_false_1_zero_m_return_mult_generic_AC_RND_CONV_false_1_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_1_r_zero_return_mult_generic_AC_RND_CONV_false_1_r_zero_nor_mdf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w3
      = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_1_else_2_else_return_mult_generic_AC_RND_CONV_false_1_else_2_else_and_nl,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_1_lor_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_3_else_2_else_return_mult_generic_AC_RND_CONV_false_3_else_2_else_and_nl
      = MUX_v_11_2_2(11'b00000000000, return_mult_generic_AC_RND_CONV_false_else_2_else_else_mux_2,
      return_mult_generic_AC_RND_CONV_false_3_zero_m_return_mult_generic_AC_RND_CONV_false_3_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_3_r_zero_return_mult_generic_AC_RND_CONV_false_3_r_zero_nor_mdf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_3_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w7
      = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_3_else_2_else_return_mult_generic_AC_RND_CONV_false_3_else_2_else_and_nl,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_3_lor_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_3_do_sub_sva_1 = ~((stage_PE_1_x_im_d_sva[63])
      ^ (out_f_d_rsci_q_d[63]));
  assign return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1 = (stage_PE_1_x_im_d_sva[63])
      ^ (out_f_d_rsci_q_d[63]);
  assign return_extract_41_return_extract_41_or_1_cse_sva_1 = (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[61:52]!=10'b0000000000);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_18,
      z_out_17, z_out_18[11]);
  assign return_add_generic_AC_RND_CONV_false_1_op2_mu_51_1_lpi_3_dfm_mx0 = MUX_v_51_2_2((out_f_d_rsci_q_d[50:0]),
      (out_f_d_rsci_q_d[51:1]), return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp);
  assign return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1 = (out_f_d_rsci_q_d[0])
      & return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1,
      and_dcpl_216);
  assign return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0
      = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0, return_add_generic_AC_RND_CONV_false_1_op2_mu_51_1_lpi_3_dfm_mx0,
      and_dcpl_216);
  assign return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_0_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1, and_dcpl_216);
  assign return_add_generic_AC_RND_CONV_false_1_e1_eq_e2_equal_tmp = (stage_PE_1_x_im_d_sva[62:52])
      == (out_f_d_rsci_q_d[62:52]);
  assign return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_and_1_cse
      = z_out_3_52 & return_add_generic_AC_RND_CONV_false_1_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_1_op1_smaller_lor_lpi_3_dfm_2 = return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_and_1_cse
      | (z_out_18[11]);
  assign return_add_generic_AC_RND_CONV_false_1_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_40[54]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_40[53]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_40[52]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_40[51]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_40[50]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_40[49]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_40[48]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_40[47]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_40[46]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_40[45]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_40[44]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_40[43]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_40[42]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_40[41]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_40[40]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_40[39]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_40[38]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_40[37]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_40[36]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_40[35]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_40[34]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_40[33]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_40[32]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_40[31]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_40[30]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_40[29]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_40[28]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_40[27]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_40[26]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_40[25]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_40[24]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_40[23]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_40[22]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_40[21]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_40[20]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_40[19]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_40[18]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_40[17]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_40[16]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_40[15]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_40[14]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_40[13]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_40[12]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_40[11]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_40[10]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_40[9]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_40[8]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_40[7]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_40[6]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_40[5]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_40[4]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_40[3]))) | (return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_40[2])));
  assign return_add_generic_AC_RND_CONV_false_3_e_dif_qr_lpi_3_dfm_mx0_10_0 = MUX_v_11_2_2((z_out_18[10:0]),
      (z_out_17[10:0]), z_out_18[11]);
  assign return_add_generic_AC_RND_CONV_false_3_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_38[54]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_38[53]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_38[52]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_38[51]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_38[50]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_38[49]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_38[48]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_38[47]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_38[46]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_38[45]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_38[44]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_38[43]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_38[42]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_38[41]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_38[40]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_38[39]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_38[38]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_38[37]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_38[36]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_38[35]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_38[34]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_38[33]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_38[32]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_38[31]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_38[30]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_38[29]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_38[28]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_38[27]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_38[26]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_38[25]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_38[24]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_38[23]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_38[22]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_38[21]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_38[20]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_38[19]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_38[18]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_38[17]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_38[16]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_38[15]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_38[14]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_38[13]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_38[12]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_38[11]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_38[10]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_38[9]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_38[8]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_38[7]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_38[6]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_38[5]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_38[4]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_38[3]))) | (return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_38[2])));
  assign return_add_generic_AC_RND_CONV_false_1_e_dif_qelse_return_add_generic_AC_RND_CONV_false_1_e_dif_qelse_and_cse
      = (z_out_17[11]) & (z_out_18[11]);
  assign return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_3_e_dif_qr_lpi_3_dfm_mx0_10_0[10:6]!=5'b00000)
      | return_add_generic_AC_RND_CONV_false_1_e_dif_qelse_return_add_generic_AC_RND_CONV_false_1_e_dif_qelse_and_cse;
  assign return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_3_e_dif_qr_lpi_3_dfm_mx0_10_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_1_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif_sat_or_cse = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_1_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_1_e_dif_sat_or_1_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt = ({1'b1 ,
      (~ (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[61:52]))}) + conv_u2s_10_11(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[61:52])
      + 11'b00000000001;
  assign return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt = nl_return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt[10:0];
  assign return_add_generic_AC_RND_CONV_false_4_e_dif_qif_acc_pmx_lpi_3_dfm_mx0_9_0
      = MUX_v_10_2_2((return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp[9:0]),
      (return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt[9:0]), return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp[10]);
  assign nl_return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp = ({1'b1 , (~ (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[61:52]))})
      + conv_u2s_10_11(BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[61:52])
      + 11'b00000000001;
  assign return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp = nl_return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp[10:0];
  assign return_add_generic_AC_RND_CONV_false_4_op1_mu_52_lpi_3_dfm_1 = (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[51])
      | return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_or_tmp;
  assign return_add_generic_AC_RND_CONV_false_4_op1_mu_51_1_lpi_3_dfm_mx0 = MUX_v_51_2_2((BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[50:0]),
      (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[51:1]), return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_or_tmp);
  assign return_add_generic_AC_RND_CONV_false_4_op1_mu_0_lpi_3_dfm_1 = (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[0])
      & return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_or_tmp;
  assign return_add_generic_AC_RND_CONV_false_4_op2_mu_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_extract_41_return_extract_41_or_1_cse_sva_1,
      (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[51]), return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_if_1_return_add_generic_AC_RND_CONV_false_17_op2_normal_return_extract_41_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_4_op2_mu_51_1_lpi_3_dfm_mx0 = MUX_v_51_2_2((r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[51:1]),
      (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[50:0]), return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_if_1_return_add_generic_AC_RND_CONV_false_17_op2_normal_return_extract_41_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_4_op2_mu_0_lpi_3_dfm_1 = (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[0])
      & (~ return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_if_1_return_add_generic_AC_RND_CONV_false_17_op2_normal_return_extract_41_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_17_e1_eq_e2_equal_tmp = (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[61:52])
      == (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[61:52]);
  assign nl_return_add_generic_AC_RND_CONV_false_18_ma1_lt_ma2_acc_2_nl = ({1'b1
      , (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[51:0])}) + conv_u2u_52_53(~
      (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[51:0])) +
      53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_18_ma1_lt_ma2_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_18_ma1_lt_ma2_acc_2_nl[52:0];
  assign return_add_generic_AC_RND_CONV_false_4_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_4_op1_smaller_oelse_and_1_cse
      = (readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_18_ma1_lt_ma2_acc_2_nl))
      & return_add_generic_AC_RND_CONV_false_17_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_17_op1_smaller_lor_lpi_3_dfm_2 = return_add_generic_AC_RND_CONV_false_4_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_4_op1_smaller_oelse_and_1_cse
      | (return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp[10]);
  assign return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_if_1_return_add_generic_AC_RND_CONV_false_17_op2_normal_return_extract_41_nor_tmp
      = ~((r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[61:52]!=10'b0000000000));
  assign return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_or_tmp
      = (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[61:52]!=10'b0000000000);
  assign return_add_generic_AC_RND_CONV_false_7_op_bigger_mux_6_itm = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1,
      BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0, and_dcpl_220);
  assign or_1477_tmp = ((~ return_add_generic_AC_RND_CONV_false_18_acc_2_itm_10)
      & (fsm_output[23])) | ((~(return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11
      | (return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp[53]))) & (fsm_output[30]));
  assign return_mult_generic_AC_RND_CONV_false_1_if_nor_ovfl_sva_1 = ~((return_mult_generic_AC_RND_CONV_false_1_exp_acc_tmp[9:6]==4'b1111));
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_4_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_4_op2_mu_0_lpi_3_dfm_1,
      and_dcpl_225);
  assign and_287_nl = and_dcpl_231 & (~(return_extract_12_m_zero_sva & operator_11_true_return_13_sva))
      & and_dcpl_229 & (~(return_extract_15_return_extract_15_nor_cse_sva & return_extract_15_m_zero_sva));
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2 =
      MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_r_nan_sva_1, (z_out[51]),
      and_287_nl);
  assign and_292_nl = or_dcpl_450 & (~(operator_11_true_return_1_sva | operator_11_true_49_operator_11_true_49_and_tmp))
      & (~((z_out_55[11]) | return_mult_generic_AC_RND_CONV_false_4_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_4_exp_ovf_oif_aelse_and_tmp))
      & (~(return_extract_49_m_zero_return_extract_49_m_zero_nor_tmp & return_extract_49_return_extract_49_nor_tmp));
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx6 =
      MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_4_r_nan_sva_1, (r_rnd_dummy_4_51_0_sva_1[51]),
      and_292_nl);
  assign return_add_generic_AC_RND_CONV_false_4_do_sub_sva_1 = ~((BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[63])
      ^ inverse_lpi_1_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_1_r_nan_sva_1 = return_add_generic_AC_RND_CONV_false_14_op2_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_8_op1_nan_sva_1 | (return_mult_generic_AC_RND_CONV_false_op1_zero_sva_1
      & return_extract_17_and_tmp) | (return_extract_16_and_tmp & return_extract_22_and_1_tmp);
  assign return_mult_generic_AC_RND_CONV_false_2_r_nan_sva_1 = (operator_11_true_19_operator_11_true_19_and_tmp
      & (~ return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp)) | (return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1
      & return_mult_generic_AC_RND_CONV_false_2_op2_inf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_5_r_nan_sva_1 = (operator_11_true_51_operator_11_true_51_and_tmp
      & (~ return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp)) | (return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1
      & return_mult_generic_AC_RND_CONV_false_5_op2_inf_sva_1);
  assign return_add_generic_AC_RND_CONV_false_12_if_2_return_add_generic_AC_RND_CONV_false_12_if_2_nor_mx3w0
      = ~(operator_11_true_return_15_sva | (~ (stage_PE_1_x_im_d_sva[63])));
  assign return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_tmp
      = (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1!=11'b00000000000);
  assign return_add_generic_AC_RND_CONV_false_11_if_2_return_add_generic_AC_RND_CONV_false_11_if_2_nor_mx3w0
      = ~(return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 | (~ (stage_PE_1_x_re_d_sva[63])));
  assign return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp
      = (return_mult_generic_AC_RND_CONV_false_3_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w7!=11'b00000000000);
  assign return_add_generic_AC_RND_CONV_false_5_do_sub_sva_1 = (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[63])
      ^ inverse_lpi_1_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_7_if_2_return_add_generic_AC_RND_CONV_false_7_if_2_and_1_mx1w0
      = stage_PE_1_tmp_im_d_1_lpi_3_dfm_63 & stage_PE_1_tmp_re_d_1_lpi_3_dfm_63;
  assign return_add_generic_AC_RND_CONV_false_7_r_sign_mux_1_nl = MUX_s_1_2_2(stage_PE_1_tmp_re_d_1_lpi_3_dfm_63,
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_63, return_add_generic_AC_RND_CONV_false_7_op1_smaller_lor_lpi_3_dfm_2);
  assign nand_84_nl = ~(return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm , return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm
      , reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1
      , return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1
      , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1})));
  assign return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_if_2_return_add_generic_AC_RND_CONV_false_7_if_2_and_1_mx1w0,
      return_add_generic_AC_RND_CONV_false_7_r_sign_mux_1_nl, nand_84_nl);
  assign return_add_generic_AC_RND_CONV_false_8_if_2_return_add_generic_AC_RND_CONV_false_8_if_2_and_1_mx2w0
      = stage_PE_1_tmp_im_d_1_lpi_3_dfm_63 & stage_PE_1_tmp_im_d_1_lpi_3_dfm_51;
  assign return_add_generic_AC_RND_CONV_false_20_r_sign_mux_1_nl = MUX_s_1_2_2(stage_PE_1_tmp_im_d_1_lpi_3_dfm_51,
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_63, or_450_cse);
  assign nand_85_nl = ~(return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm
      , reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1
      , return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1
      , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1})));
  assign return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_if_2_return_add_generic_AC_RND_CONV_false_8_if_2_and_1_mx2w0,
      return_add_generic_AC_RND_CONV_false_20_r_sign_mux_1_nl, nand_85_nl);
  assign return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp
      = ~((stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_1!=10'b0000000000) | stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0);
  assign return_add_generic_AC_RND_CONV_false_7_op1_inf_sva_1 = operator_11_true_return_1_sva
      & return_extract_12_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_2_lor_lpi_3_dfm_1 = return_mult_generic_AC_RND_CONV_false_2_op2_inf_sva_1
      | ((return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_1==12'b011111111110)
      & return_mult_generic_AC_RND_CONV_false_2_e_incr_lpi_3_dfm_2) | (z_out_24[11])
      | return_mult_generic_AC_RND_CONV_false_2_r_nan_sva_1;
  assign return_add_generic_AC_RND_CONV_false_10_op1_inf_sva_1 = operator_11_true_return_26_sva
      & return_extract_44_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_5_lor_lpi_3_dfm_1 = return_mult_generic_AC_RND_CONV_false_5_op2_inf_sva_1
      | ((return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_1==12'b011111111110)
      & return_mult_generic_AC_RND_CONV_false_5_e_incr_lpi_3_dfm_2) | (z_out_24[11])
      | return_mult_generic_AC_RND_CONV_false_5_r_nan_sva_1;
  assign return_add_generic_AC_RND_CONV_false_2_do_sub_sva_1 = ~((out_f_d_rsci_q_d[63])
      ^ (stage_PE_1_tmp_im_d_1_sva_1_63_51[12]));
  assign return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1 = (stage_PE_1_x_im_d_sva[63])
      ^ (in_f_d_rsci_q_d[63]);
  assign return_add_generic_AC_RND_CONV_false_13_do_sub_sva_1 = (in_f_d_rsci_q_d[63])
      ^ (stage_PE_1_tmp_im_d_1_sva_1_63_51[12]);
  assign return_add_generic_AC_RND_CONV_false_do_sub_sva_1 = (out_f_d_rsci_q_d[63])
      ^ (stage_PE_1_tmp_im_d_1_sva_1_63_51[12]);
  assign return_add_generic_AC_RND_CONV_false_16_do_sub_sva_1 = ~((stage_PE_1_x_im_d_sva[63])
      ^ (in_f_d_rsci_q_d[63]));
  assign return_add_generic_AC_RND_CONV_false_15_do_sub_sva_1 = ~((in_f_d_rsci_q_d[63])
      ^ (stage_PE_1_tmp_im_d_1_sva_1_63_51[12]));
  assign return_add_generic_AC_RND_CONV_false_5_if_7_not_7_nl = ~ return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (r_rnd_dummy_1_51_0_sva_1[50:0]), return_add_generic_AC_RND_CONV_false_5_if_7_not_7_nl);
  assign return_mult_generic_AC_RND_CONV_false_3_oelse_3_return_mult_generic_AC_RND_CONV_false_3_if_3_nor_nl
      = ~((~ return_mult_generic_AC_RND_CONV_false_3_zero_m_return_mult_generic_AC_RND_CONV_false_3_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_3_r_zero_return_mult_generic_AC_RND_CONV_false_3_r_zero_nor_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_3_lor_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (z_out[50:0]), return_mult_generic_AC_RND_CONV_false_3_oelse_3_return_mult_generic_AC_RND_CONV_false_3_if_3_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_4_if_7_not_6_nl = ~ return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_mx0w2 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_4_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_4_if_7_not_6_nl);
  assign return_add_generic_AC_RND_CONV_false_8_if_7_return_add_generic_AC_RND_CONV_false_8_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_8_exception_sva_1 | return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_mx0w4 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_5_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_8_if_7_return_add_generic_AC_RND_CONV_false_8_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_5_if_7_not_5_nl = ~ return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_mx0w5 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_2, return_add_generic_AC_RND_CONV_false_5_if_7_not_5_nl);
  assign return_add_generic_AC_RND_CONV_false_21_if_7_return_add_generic_AC_RND_CONV_false_21_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_21_exception_sva_1 | return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_mx0w6 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_21_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_21_if_7_return_add_generic_AC_RND_CONV_false_21_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_5_mux_20_nl = MUX_v_56_2_2((z_out_31[56:1]),
      (~ (z_out_31[56:1])), return_add_generic_AC_RND_CONV_false_12_mux_itm);
  assign return_add_generic_AC_RND_CONV_false_5_mux_19_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_5_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_5_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_12_mux_itm);
  assign nl_return_add_generic_AC_RND_CONV_false_5_res_mant_4_sva_1 = ({return_add_generic_AC_RND_CONV_false_5_mux_20_nl
      , return_add_generic_AC_RND_CONV_false_5_mux_19_nl}) + conv_u2u_56_57({return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm
      , return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm
      , return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm , 3'b000}) +
      conv_u2u_1_57(return_add_generic_AC_RND_CONV_false_12_mux_itm);
  assign return_add_generic_AC_RND_CONV_false_5_res_mant_4_sva_1 = nl_return_add_generic_AC_RND_CONV_false_5_res_mant_4_sva_1[56:0];
  assign return_add_generic_AC_RND_CONV_false_6_mux_31_nl = MUX_v_56_2_2((z_out_32[56:1]),
      (~ (z_out_32[56:1])), return_add_generic_AC_RND_CONV_false_13_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_6_mux_30_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_6_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_13_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_6_op_bigger_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm,
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50, return_add_generic_AC_RND_CONV_false_19_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_6_op_bigger_mux_2_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_19_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_6_op_bigger_mux_9_nl = MUX_v_50_2_2(reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1,
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0, return_add_generic_AC_RND_CONV_false_19_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_6_op_bigger_mux_3_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_19_op1_smaller_lor_lpi_3_dfm_2);
  assign nl_return_add_generic_AC_RND_CONV_false_6_res_mant_4_sva_1 = ({return_add_generic_AC_RND_CONV_false_6_mux_31_nl
      , return_add_generic_AC_RND_CONV_false_6_mux_30_nl}) + conv_u2u_56_57({return_add_generic_AC_RND_CONV_false_6_op_bigger_mux_1_nl
      , return_add_generic_AC_RND_CONV_false_6_op_bigger_mux_2_nl , return_add_generic_AC_RND_CONV_false_6_op_bigger_mux_9_nl
      , return_add_generic_AC_RND_CONV_false_6_op_bigger_mux_3_nl , 3'b000}) + conv_u2u_1_57(return_add_generic_AC_RND_CONV_false_13_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_6_res_mant_4_sva_1 = nl_return_add_generic_AC_RND_CONV_false_6_res_mant_4_sva_1[56:0];
  assign return_add_generic_AC_RND_CONV_false_8_mux_25_nl = MUX_v_56_2_2((z_out_33[56:1]),
      (~ (z_out_33[56:1])), return_add_generic_AC_RND_CONV_false_15_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_8_mux_24_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_8_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_15_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_8_op_bigger_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1, or_451_cse);
  assign return_add_generic_AC_RND_CONV_false_8_op_bigger_mux_2_nl = MUX_s_1_2_2(drf_qr_lval_14_smx_0_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0, or_451_cse);
  assign return_add_generic_AC_RND_CONV_false_8_op_bigger_mux_4_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1, or_451_cse);
  assign nl_return_add_generic_AC_RND_CONV_false_8_res_mant_4_sva_1 = ({return_add_generic_AC_RND_CONV_false_8_mux_25_nl
      , return_add_generic_AC_RND_CONV_false_8_mux_24_nl}) + conv_u2u_56_57({return_add_generic_AC_RND_CONV_false_8_op_bigger_mux_1_nl
      , return_add_generic_AC_RND_CONV_false_8_op_bigger_mux_2_nl , z_out_10 , return_add_generic_AC_RND_CONV_false_8_op_bigger_mux_4_nl
      , 3'b000}) + conv_u2u_1_57(return_add_generic_AC_RND_CONV_false_15_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_8_res_mant_4_sva_1 = nl_return_add_generic_AC_RND_CONV_false_8_res_mant_4_sva_1[56:0];
  assign return_add_generic_AC_RND_CONV_false_5_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_5_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_5_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign nl_return_add_generic_AC_RND_CONV_false_4_res_mant_4_sva_1 = ({return_add_generic_AC_RND_CONV_false_4_res_mant_conc_2_itm_56_1
      , return_add_generic_AC_RND_CONV_false_5_mux_nl}) + conv_u2u_56_57({return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm
      , return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm
      , return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm , 3'b000}) +
      conv_u2u_1_57(return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_4_res_mant_4_sva_1 = nl_return_add_generic_AC_RND_CONV_false_4_res_mant_4_sva_1[56:0];
  assign return_add_generic_AC_RND_CONV_false_10_mux_26_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_10_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_10_op_bigger_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse);
  assign return_add_generic_AC_RND_CONV_false_10_op_bigger_mux_1_nl = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0[50]),
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50, return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse);
  assign return_add_generic_AC_RND_CONV_false_10_op_bigger_mux_2_nl = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0[49:0]),
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0, return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse);
  assign return_add_generic_AC_RND_CONV_false_10_op_bigger_mux_3_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse);
  assign nl_return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_2 = ({return_add_generic_AC_RND_CONV_false_4_res_mant_conc_2_itm_56_1
      , return_add_generic_AC_RND_CONV_false_10_mux_26_nl}) + conv_u2u_56_57({return_add_generic_AC_RND_CONV_false_10_op_bigger_mux_nl
      , return_add_generic_AC_RND_CONV_false_10_op_bigger_mux_1_nl , return_add_generic_AC_RND_CONV_false_10_op_bigger_mux_2_nl
      , return_add_generic_AC_RND_CONV_false_10_op_bigger_mux_3_nl , 3'b000}) + conv_u2u_1_57(return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_2 = nl_return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_2[56:0];
  assign return_add_generic_AC_RND_CONV_false_21_mux_23_nl = MUX_v_56_2_2((z_out_33[56:1]),
      (~ (z_out_33[56:1])), return_add_generic_AC_RND_CONV_false_13_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_21_mux_22_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_21_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_13_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_21_op_bigger_mux_1_nl = MUX_s_1_2_2(drf_qr_lval_14_smx_0_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_21_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_21_op_bigger_mux_2_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_21_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_21_op_bigger_mux_4_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_21_op1_smaller_lor_lpi_3_dfm_2);
  assign nl_return_add_generic_AC_RND_CONV_false_21_res_mant_4_sva_1 = ({return_add_generic_AC_RND_CONV_false_21_mux_23_nl
      , return_add_generic_AC_RND_CONV_false_21_mux_22_nl}) + conv_u2u_56_57({return_add_generic_AC_RND_CONV_false_21_op_bigger_mux_1_nl
      , return_add_generic_AC_RND_CONV_false_21_op_bigger_mux_2_nl , z_out_10 , return_add_generic_AC_RND_CONV_false_21_op_bigger_mux_4_nl
      , 3'b000}) + conv_u2u_1_57(return_add_generic_AC_RND_CONV_false_13_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_21_res_mant_4_sva_1 = nl_return_add_generic_AC_RND_CONV_false_21_res_mant_4_sva_1[56:0];
  assign return_mult_generic_AC_RND_CONV_false_else_2_else_return_mult_generic_AC_RND_CONV_false_else_2_else_and_nl
      = MUX_v_11_2_2(11'b00000000000, return_mult_generic_AC_RND_CONV_false_else_2_else_else_mux_2,
      return_mult_generic_AC_RND_CONV_false_zero_m_return_mult_generic_AC_RND_CONV_false_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_r_zero_return_mult_generic_AC_RND_CONV_false_r_zero_nor_mdf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1 = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_else_2_else_return_mult_generic_AC_RND_CONV_false_else_2_else_and_nl,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_lor_lpi_3_dfm_1);
  assign drf_qr_lval_10_smx_lpi_3_dfm_mx1_10 = MUX_s_1_2_2((return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd, and_dcpl_248);
  assign drf_qr_lval_10_smx_lpi_3_dfm_mx1_9_6 = MUX_v_4_2_2((return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[9:6]),
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1, and_dcpl_248);
  assign drf_qr_lval_10_smx_lpi_3_dfm_mx1_5_0 = MUX_v_6_2_2((return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[5:0]),
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2, and_dcpl_248);
  assign return_mult_generic_AC_RND_CONV_false_4_else_2_else_else_mux_nl = MUX_v_11_2_2((return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_1_cse[10:0]),
      (z_out_55[10:0]), return_mult_generic_AC_RND_CONV_false_4_e_incr_lpi_3_dfm_2);
  assign return_mult_generic_AC_RND_CONV_false_4_else_2_else_return_mult_generic_AC_RND_CONV_false_4_else_2_else_and_nl
      = MUX_v_11_2_2(11'b00000000000, return_mult_generic_AC_RND_CONV_false_4_else_2_else_else_mux_nl,
      return_mult_generic_AC_RND_CONV_false_4_zero_m_return_mult_generic_AC_RND_CONV_false_4_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_4_r_zero_return_mult_generic_AC_RND_CONV_false_4_r_zero_nor_mdf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_4_exp_1_11_0_lpi_3_dfm_3_10_0_1 =
      MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_4_else_2_else_return_mult_generic_AC_RND_CONV_false_4_else_2_else_and_nl,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_4_lor_lpi_3_dfm_1);
  assign drf_qr_lval_10_smx_lpi_3_dfm_mx2_10 = MUX_s_1_2_2((return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd, and_dcpl_249);
  assign drf_qr_lval_10_smx_lpi_3_dfm_mx2_9_6 = MUX_v_4_2_2((return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[9:6]),
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1, and_dcpl_249);
  assign drf_qr_lval_10_smx_lpi_3_dfm_mx2_5_0 = MUX_v_6_2_2((return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[5:0]),
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2, and_dcpl_249);
  assign nl_return_add_generic_AC_RND_CONV_false_8_ma1_lt_ma2_acc_1_nl = ({1'b1 ,
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm , return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm})
      + conv_u2u_52_53({(~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx1)
      , (~ return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1)}) + 53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_8_ma1_lt_ma2_acc_1_nl = nl_return_add_generic_AC_RND_CONV_false_8_ma1_lt_ma2_acc_1_nl[52:0];
  assign and_276_cse = return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp
      & (readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_8_ma1_lt_ma2_acc_1_nl));
  assign or_451_cse = and_276_cse | (return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp[11]);
  assign nl_return_add_generic_AC_RND_CONV_false_20_ma1_lt_ma2_acc_1_nl = ({1'b1
      , BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm , return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm})
      + conv_u2u_52_53({(~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx1)
      , (~ return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1)}) + 53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_20_ma1_lt_ma2_acc_1_nl = nl_return_add_generic_AC_RND_CONV_false_20_ma1_lt_ma2_acc_1_nl[52:0];
  assign and_275_cse = return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp
      & (readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_20_ma1_lt_ma2_acc_1_nl));
  assign or_450_cse = and_275_cse | (return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp[11]);
  assign nl_return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl = ({1'b1 ,
      (out_f_d_rsci_q_d[51:0])}) + conv_u2u_52_53({(~ (stage_PE_1_tmp_im_d_1_sva_1_63_51[0]))
      , (~ stage_PE_1_tmp_im_d_1_sva_1_50_0)}) + 53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl[52:0];
  assign and_272_cse = (readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl))
      & return_add_generic_AC_RND_CONV_false_e1_eq_e2_equal_tmp;
  assign and_277_cse = return_add_generic_AC_RND_CONV_false_14_e1_eq_e2_equal_tmp
      & z_out_3_52;
  assign nl_return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl = ({1'b1
      , (in_f_d_rsci_q_d[51:0])}) + conv_u2u_52_53({(~ (stage_PE_1_tmp_im_d_1_sva_1_63_51[0]))
      , (~ stage_PE_1_tmp_im_d_1_sva_1_50_0)}) + 53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl[52:0];
  assign and_271_cse = return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp
      & (readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl));
  assign or_446_cse = and_272_cse | (z_out_17[11]);
  assign or_452_cse = and_277_cse | (z_out_18[11]);
  assign or_445_cse = and_271_cse | (z_out_17[11]);
  assign and_1029_cse = or_450_cse & (fsm_output[28]);
  assign and_1014_cse = return_add_generic_AC_RND_CONV_false_1_op1_smaller_lor_lpi_3_dfm_2
      & (fsm_output[6]);
  assign and_1032_cse = or_452_cse & (fsm_output[22]);
  assign or_956_cse = (or_445_cse & (fsm_output[24])) | (or_446_cse & (fsm_output[8]));
  assign return_add_generic_AC_RND_CONV_false_3_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_14_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_14_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_15_do_sub_sva);
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_51_mx0 = MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_3_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_3_res_rounded_lpi_3_dfm_51_0_1[51]),
      (stage_PE_1_tmp_im_d_1_sva_1_63_51[0]), {and_344_cse , and_347_cse , (~ inverse_lpi_1_dfm_1)});
  assign return_add_generic_AC_RND_CONV_false_3_if_7_return_add_generic_AC_RND_CONV_false_3_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_3_exception_sva_1 | leading_sign_57_0_1_0_15_out_2);
  assign return_add_generic_AC_RND_CONV_false_3_return_add_generic_AC_RND_CONV_false_3_and_4_nl
      = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000, (return_add_generic_AC_RND_CONV_false_3_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_3_if_7_return_add_generic_AC_RND_CONV_false_3_if_7_nor_nl);
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0 = MUX_v_51_2_2(stage_PE_1_tmp_im_d_1_sva_1_50_0,
      return_add_generic_AC_RND_CONV_false_3_return_add_generic_AC_RND_CONV_false_3_and_4_nl,
      inverse_lpi_1_dfm_1);
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_3_exception_sva_1);
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs, or_dcpl_168);
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_0 = (return_add_generic_AC_RND_CONV_false_3_mux_26
      & (~ return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_1_nl)) | return_add_generic_AC_RND_CONV_false_3_exception_sva_1;
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_1 = MUX_v_10_2_2((stage_PE_1_tmp_im_d_1_sva_1_63_51[11:2]),
      stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1, inverse_lpi_1_dfm_1);
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0 = MUX_s_1_2_2((stage_PE_1_tmp_im_d_1_sva_1_63_51[1]),
      stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_0, inverse_lpi_1_dfm_1);
  assign return_extract_13_return_extract_13_or_1_cse_sva_1 = (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_1!=10'b0000000000)
      | stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0;
  assign and_2152_nl = (return_add_generic_AC_RND_CONV_false_2_res_rounded_acc_tmp[53])
      & (~ return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0);
  assign mux_16_nl = MUX_v_10_2_2((operator_33_true_4_acc_tmp[10:1]), (return_add_generic_AC_RND_CONV_false_1_exp_plus_1_12_1_lpi_3_dfm_1[9:0]),
      and_2152_nl);
  assign not_736_nl = ~ return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0;
  assign return_add_generic_AC_RND_CONV_false_1_e_r_qelse_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(10'b0000000000,
      mux_16_nl, not_736_nl);
  assign nl_operator_33_true_4_acc_tmp = conv_s2s_7_13({operator_6_false_2_operator_6_false_2_conc_2_6_1
      , (~ (leading_sign_57_0_1_0_2_out_3[0]))}) + conv_u2s_11_13(BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0);
  assign operator_33_true_4_acc_tmp = nl_operator_33_true_4_acc_tmp[12:0];
  assign return_add_generic_AC_RND_CONV_false_1_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      z_out_21, return_add_generic_AC_RND_CONV_false_2_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_1_res_rounded_and_1_cse = (z_out_36[3])
      & ((z_out_36[0]) | (z_out_36[1]) | (z_out_36[2]) | (z_out_36[4]));
  assign nl_return_add_generic_AC_RND_CONV_false_2_res_rounded_acc_tmp = conv_u2u_53_54(z_out_36[56:4])
      + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_1_res_rounded_and_1_cse);
  assign return_add_generic_AC_RND_CONV_false_2_res_rounded_acc_tmp = nl_return_add_generic_AC_RND_CONV_false_2_res_rounded_acc_tmp[53:0];
  assign return_add_generic_AC_RND_CONV_false_14_op1_nan_sva_1 = operator_11_true_return_1_sva
      & (~ return_extract_17_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 = operator_11_true_return_13_sva
      & (~ return_extract_15_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_14_op1_inf_sva_1 = operator_11_true_return_1_sva
      & return_extract_17_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 = operator_11_true_return_13_sva
      & return_extract_15_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_1_not_6_nl = ~ (return_add_generic_AC_RND_CONV_false_2_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_1_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_2_res_rounded_acc_tmp[51:0]), return_add_generic_AC_RND_CONV_false_1_not_6_nl);
  assign and_2154_nl = (return_add_generic_AC_RND_CONV_false_res_rounded_acc_tmp[53])
      & (~ return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w0);
  assign mux_17_nl = MUX_v_10_2_2((z_out_13[10:1]), (return_add_generic_AC_RND_CONV_false_3_exp_plus_1_12_1_lpi_3_dfm_1[9:0]),
      and_2154_nl);
  assign not_738_nl = ~ return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w0;
  assign return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(10'b0000000000,
      mux_17_nl, not_738_nl);
  assign nl_operator_33_true_7_acc_1_nl = conv_s2s_11_12(z_out_52[11:1]) + 12'b000000000001;
  assign operator_33_true_7_acc_1_nl = nl_operator_33_true_7_acc_1_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_3_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      operator_33_true_7_acc_1_nl, return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_3_res_rounded_and_1_nl = (return_add_generic_AC_RND_CONV_false_3_res_rounded_asn_rndc_sva_1[3])
      & ((return_add_generic_AC_RND_CONV_false_3_res_rounded_asn_rndc_sva_1[0]) |
      (return_add_generic_AC_RND_CONV_false_3_res_rounded_asn_rndc_sva_1[1]) | (return_add_generic_AC_RND_CONV_false_3_res_rounded_asn_rndc_sva_1[2])
      | (return_add_generic_AC_RND_CONV_false_3_res_rounded_asn_rndc_sva_1[4]));
  assign nl_return_add_generic_AC_RND_CONV_false_res_rounded_acc_tmp = conv_u2u_53_54(return_add_generic_AC_RND_CONV_false_3_res_rounded_asn_rndc_sva_1[56:4])
      + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_3_res_rounded_and_1_nl);
  assign return_add_generic_AC_RND_CONV_false_res_rounded_acc_tmp = nl_return_add_generic_AC_RND_CONV_false_res_rounded_acc_tmp[53:0];
  assign return_add_generic_AC_RND_CONV_false_3_not_6_nl = ~ (return_add_generic_AC_RND_CONV_false_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_3_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_res_rounded_acc_tmp[51:0]), return_add_generic_AC_RND_CONV_false_3_not_6_nl);
  assign return_add_generic_AC_RND_CONV_false_3_if_5_or_nl = return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_15_if_5_return_add_generic_AC_RND_CONV_false_15_if_5_and_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_3_mux_10_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_3_if_5_or_nl, return_add_generic_AC_RND_CONV_false_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_3_exception_sva_1 = return_add_generic_AC_RND_CONV_false_14_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_3_mux_10_cse;
  assign return_add_generic_AC_RND_CONV_false_3_exp_plus_1_0_lpi_3_dfm_1 = (z_out_52[0])
      | (~ return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2 = ((z_out_13[11])
      | (~ return_add_generic_AC_RND_CONV_false_15_else_4_return_add_generic_AC_RND_CONV_false_15_else_4_nand_tmp))
      & return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_1_exp_plus_1_0_lpi_3_dfm_1 = (z_out_51[0])
      | (~ return_add_generic_AC_RND_CONV_false_2_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_1_if_5_or_nl = return_add_generic_AC_RND_CONV_false_1_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_2_if_5_return_add_generic_AC_RND_CONV_false_2_if_5_and_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_1_mux_16_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_1_if_5_or_nl, return_add_generic_AC_RND_CONV_false_2_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_1_exception_sva_1 = return_add_generic_AC_RND_CONV_false_14_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_1_mux_16_cse;
  assign return_add_generic_AC_RND_CONV_false_1_r_inf_lpi_3_dfm_2 = ((operator_33_true_4_acc_tmp[11])
      | (~ return_add_generic_AC_RND_CONV_false_2_else_4_return_add_generic_AC_RND_CONV_false_2_else_4_nand_tmp))
      & return_add_generic_AC_RND_CONV_false_2_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_5_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm
      & (~ (z_out_39[54]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[50])
      & (~ (z_out_39[53]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[49])
      & (~ (z_out_39[52]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[48])
      & (~ (z_out_39[51]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[47])
      & (~ (z_out_39[50]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[46])
      & (~ (z_out_39[49]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[45])
      & (~ (z_out_39[48]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[44])
      & (~ (z_out_39[47]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[43])
      & (~ (z_out_39[46]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[42])
      & (~ (z_out_39[45]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[41])
      & (~ (z_out_39[44]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[40])
      & (~ (z_out_39[43]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[39])
      & (~ (z_out_39[42]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[38])
      & (~ (z_out_39[41]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[37])
      & (~ (z_out_39[40]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[36])
      & (~ (z_out_39[39]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[35])
      & (~ (z_out_39[38]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[34])
      & (~ (z_out_39[37]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[33])
      & (~ (z_out_39[36]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[32])
      & (~ (z_out_39[35]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[31])
      & (~ (z_out_39[34]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[30])
      & (~ (z_out_39[33]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[29])
      & (~ (z_out_39[32]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[28])
      & (~ (z_out_39[31]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[27])
      & (~ (z_out_39[30]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[26])
      & (~ (z_out_39[29]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[25])
      & (~ (z_out_39[28]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[24])
      & (~ (z_out_39[27]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[23])
      & (~ (z_out_39[26]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[22])
      & (~ (z_out_39[25]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[21])
      & (~ (z_out_39[24]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[20])
      & (~ (z_out_39[23]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[19])
      & (~ (z_out_39[22]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[18])
      & (~ (z_out_39[21]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[17])
      & (~ (z_out_39[20]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[16])
      & (~ (z_out_39[19]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[15])
      & (~ (z_out_39[18]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[14])
      & (~ (z_out_39[17]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[13])
      & (~ (z_out_39[16]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[12])
      & (~ (z_out_39[15]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[11])
      & (~ (z_out_39[14]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[10])
      & (~ (z_out_39[13]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[9])
      & (~ (z_out_39[12]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[8])
      & (~ (z_out_39[11]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[7])
      & (~ (z_out_39[10]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[6])
      & (~ (z_out_39[9]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[5])
      & (~ (z_out_39[8]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[4])
      & (~ (z_out_39[7]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[3])
      & (~ (z_out_39[6]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[2])
      & (~ (z_out_39[5]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[1])
      & (~ (z_out_39[4]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[0])
      & (~ (z_out_39[3]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm
      & (~ (z_out_39[2])));
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_mx0w1 = MUX_s_1_2_2(stage_PE_1_tmp_im_d_1_lpi_3_dfm_51,
      (stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0[50]), return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_cse_sva);
  assign return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_mx0w4[0])
      & (~ return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1 = (stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0[0])
      & (~ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_cse_sva);
  assign return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50_mx2 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm_mx1,
      (return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_mx0w4[50]), return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp);
  assign return_extract_12_return_extract_12_or_1_tmp = (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_1!=10'b0000000000)
      | stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0;
  assign BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx1 = MUX_s_1_2_2((r_rnd_dummy_1_51_0_sva_1[51]),
      return_add_generic_AC_RND_CONV_false_10_do_sub_sva, return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_extract_45_return_extract_45_or_1_cse_sva_1 = (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_1!=10'b0000000000)
      | stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0;
  assign return_extract_44_return_extract_44_or_1_tmp = (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx1_10_1!=10'b0000000000)
      | stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx1_0;
  assign and_328_nl = and_dcpl_231 & or_dcpl_450 & and_dcpl_229 & (~(return_extract_17_m_zero_sva
      & return_extract_15_return_extract_15_nor_cse_sva));
  assign BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx3 = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_3_r_nan_sva_1,
      (z_out[51]), and_328_nl);
  assign return_add_generic_AC_RND_CONV_false_7_e_r_qelse_not_2_nl = ~ return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs_mx0w0;
  assign return_add_generic_AC_RND_CONV_false_7_e_r_qelse_return_add_generic_AC_RND_CONV_false_7_e_r_qelse_and_nl
      = MUX_v_10_2_2(10'b0000000000, z_out_44, return_add_generic_AC_RND_CONV_false_7_e_r_qelse_not_2_nl);
  assign return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_7_e_r_qelse_return_add_generic_AC_RND_CONV_false_7_e_r_qelse_and_nl,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_7_exception_sva_1);
  assign return_add_generic_AC_RND_CONV_false_21_mux_16_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_and_10_9,
      (return_add_generic_AC_RND_CONV_false_21_exp_plus_1_12_1_lpi_3_dfm_1[9]), return_add_generic_AC_RND_CONV_false_21_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_21_e_r_qelse_return_add_generic_AC_RND_CONV_false_21_e_r_qelse_and_nl
      = return_add_generic_AC_RND_CONV_false_21_mux_16_nl & (~ return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs_mx0w0);
  assign return_add_generic_AC_RND_CONV_false_21_mux_24_nl = MUX_v_9_2_2(return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_and_10_8_0,
      (return_add_generic_AC_RND_CONV_false_21_exp_plus_1_12_1_lpi_3_dfm_1[8:0]),
      return_add_generic_AC_RND_CONV_false_21_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_21_e_r_qelse_not_3_nl = ~ return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs_mx0w0;
  assign return_add_generic_AC_RND_CONV_false_21_e_r_qelse_return_add_generic_AC_RND_CONV_false_21_e_r_qelse_and_2_nl
      = MUX_v_9_2_2(9'b000000000, return_add_generic_AC_RND_CONV_false_21_mux_24_nl,
      return_add_generic_AC_RND_CONV_false_21_e_r_qelse_not_3_nl);
  assign return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_mx1w0 = MUX_v_10_2_2(({return_add_generic_AC_RND_CONV_false_21_e_r_qelse_return_add_generic_AC_RND_CONV_false_21_e_r_qelse_and_nl
      , return_add_generic_AC_RND_CONV_false_21_e_r_qelse_return_add_generic_AC_RND_CONV_false_21_e_r_qelse_and_2_nl}),
      10'b1111111111, return_add_generic_AC_RND_CONV_false_21_exception_sva_1);
  assign return_add_generic_AC_RND_CONV_false_6_exp_plus_1_0_lpi_3_dfm_1 = (operator_6_false_13_acc_psp_sva_1[0])
      | (~ return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_8_mux_17_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_and_8,
      return_add_generic_AC_RND_CONV_false_8_exp_plus_1_0_lpi_3_dfm_1, z_out_46[53]);
  assign or_230_nl = or_dcpl_201 | and_dcpl_127 | operator_11_true_return_17_sva;
  assign return_add_generic_AC_RND_CONV_false_8_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs, or_230_nl);
  assign return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_8_mux_17_nl
      & (~ return_add_generic_AC_RND_CONV_false_8_e_r_qelse_mux_1_nl)) | return_add_generic_AC_RND_CONV_false_8_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm_mx1
      = MUX_s_1_2_2((stage_PE_1_x_im_d_sva[52]), return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm,
      return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse);
  assign return_add_generic_AC_RND_CONV_false_21_mux_17_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_and_8,
      return_add_generic_AC_RND_CONV_false_21_exp_plus_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_21_res_rounded_acc_tmp[53]);
  assign or_249_nl = or_dcpl_201 | and_dcpl_132 | operator_11_true_return_17_sva;
  assign return_add_generic_AC_RND_CONV_false_21_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs, or_249_nl);
  assign return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_21_mux_17_nl
      & (~ return_add_generic_AC_RND_CONV_false_21_e_r_qelse_mux_1_nl)) | return_add_generic_AC_RND_CONV_false_21_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_and_nl
      = (({return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm , return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm
      , reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1
      , return_add_generic_AC_RND_CONV_false_6_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50
      , return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0
      , return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1})) & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva;
  assign return_add_generic_AC_RND_CONV_false_6_mux_6_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_r_sign_mux_2,
      return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_nor_2,
      return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_and_nl);
  assign stage_d_mul_return_d_2_63_sva_1 = inverse_lpi_1_dfm_1 ^ return_add_generic_AC_RND_CONV_false_6_mux_6_nl;
  assign return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_and_nl
      = (({return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm
      , reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1
      , return_add_generic_AC_RND_CONV_false_19_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50 , return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0
      , return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm})) & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva;
  assign return_add_generic_AC_RND_CONV_false_19_mux_6_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_r_sign_mux_2,
      return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_nor_2,
      return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_and_nl);
  assign stage_d_mul_return_d_5_63_sva_1 = inverse_lpi_1_dfm_1 ^ return_add_generic_AC_RND_CONV_false_19_mux_6_nl;
  assign stage_d_mul_return_d_1_63_sva_1 = stage_PE_1_tmp_im_d_1_lpi_3_dfm_63 ^ return_add_generic_AC_RND_CONV_false_18_mux_itm;
  assign and_344_cse = (or_dcpl_167 | and_dcpl_114 | operator_11_true_return_13_sva
      | leading_sign_57_0_1_0_15_out_2) & inverse_lpi_1_dfm_1;
  assign and_347_cse = (~((~((~ (z_out_13[11])) & return_add_generic_AC_RND_CONV_false_15_else_4_return_add_generic_AC_RND_CONV_false_15_else_4_nand_tmp))
      & return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1)) & (~(return_add_generic_AC_RND_CONV_false_15_if_5_return_add_generic_AC_RND_CONV_false_15_if_5_and_1_tmp
      & (return_add_generic_AC_RND_CONV_false_res_rounded_acc_tmp[53]))) & and_dcpl_254
      & (~ leading_sign_57_0_1_0_15_out_2) & inverse_lpi_1_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_16_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_14_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_14_op1_inf_sva_1
      & return_mult_generic_AC_RND_CONV_false_op1_zero_sva_1 & return_add_generic_AC_RND_CONV_false_15_do_sub_sva);
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_51_mx1 = MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_16_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_3_res_rounded_lpi_3_dfm_51_0_1[51]),
      (stage_PE_1_tmp_im_d_1_sva_1_63_51[0]), {and_344_cse , and_347_cse , (~ inverse_lpi_1_dfm_1)});
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w4_10_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_16_exception_sva_1);
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_5_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs, or_dcpl_168);
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w4_0 = (return_add_generic_AC_RND_CONV_false_3_mux_26
      & (~ return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_5_nl)) | return_add_generic_AC_RND_CONV_false_16_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_1_return_add_generic_AC_RND_CONV_false_6_op2_normal_return_extract_13_nor_tmp
      = ~((stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_1!=10'b0000000000) | stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0);
  assign return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_tmp
      = ~((stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_1!=10'b0000000000) | stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0);
  assign return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp
      = ~((stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx1_10_1!=10'b0000000000) | stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx1_0);
  assign return_add_generic_AC_RND_CONV_false_25_if_5_return_add_generic_AC_RND_CONV_false_25_if_5_and_tmp
      = (return_add_generic_AC_RND_CONV_false_25_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_25_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_25_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_25_if_5_or_nl = return_add_generic_AC_RND_CONV_false_25_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_25_if_5_return_add_generic_AC_RND_CONV_false_25_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_25_mux_10_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_25_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_25_if_5_or_nl, return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_25_exception_sva_1 = return_add_generic_AC_RND_CONV_false_23_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_23_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_25_mux_10_nl;
  assign return_add_generic_AC_RND_CONV_false_17_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10
      | (~((operator_33_true_34_acc_psp_1_sva_1!=12'b000000000000)));
  assign return_add_generic_AC_RND_CONV_false_17_mux_15_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10,
      return_add_generic_AC_RND_CONV_false_17_if_5_or_1_nl, return_add_generic_AC_RND_CONV_false_17_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qelse_or_svs_1 = leading_sign_57_0_1_0_17_out_2
      | (~ return_add_generic_AC_RND_CONV_false_17_mux_15_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_6_acc_2_nl =  -(operator_33_true_12_acc_tmp[11:0]);
  assign return_add_generic_AC_RND_CONV_false_6_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_6_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_6_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_11_acc_2_nl =  -(z_out_48[11:0]);
  assign return_add_generic_AC_RND_CONV_false_11_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_11_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_11_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_19_acc_2_nl =  -(z_out_16[11:0]);
  assign return_add_generic_AC_RND_CONV_false_19_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_19_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_19_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_19_acc_2_nl);
  assign return_add_generic_AC_RND_CONV_false_16_if_7_return_add_generic_AC_RND_CONV_false_16_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_16_exception_sva_1 | leading_sign_57_0_1_0_15_out_2);
  assign return_add_generic_AC_RND_CONV_false_16_return_add_generic_AC_RND_CONV_false_16_and_4_nl
      = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000, (return_add_generic_AC_RND_CONV_false_3_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_16_if_7_return_add_generic_AC_RND_CONV_false_16_if_7_nor_nl);
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx1 = MUX_v_51_2_2(stage_PE_1_tmp_im_d_1_sva_1_50_0,
      return_add_generic_AC_RND_CONV_false_16_return_add_generic_AC_RND_CONV_false_16_and_4_nl,
      inverse_lpi_1_dfm_1);
  assign nl_operator_33_true_13_acc_nl = conv_s2s_11_12(operator_6_false_13_acc_psp_sva_1[11:1])
      + 12'b000000000001;
  assign operator_33_true_13_acc_nl = nl_operator_33_true_13_acc_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_6_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      operator_33_true_13_acc_nl, return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1);
  assign nl_return_add_generic_AC_RND_CONV_false_9_e_dif1_acc_1_tmp = ({1'b1 , (stage_PE_1_x_re_d_sva[62:52])})
      + conv_u2s_11_12({(~ return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1)
      , (~ return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1)}) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_9_e_dif1_acc_1_tmp = nl_return_add_generic_AC_RND_CONV_false_9_e_dif1_acc_1_tmp[11:0];
  assign nl_return_add_generic_AC_RND_CONV_false_10_e_dif1_acc_1_tmp = ({1'b1 , (stage_PE_1_x_im_d_sva[62:52])})
      + conv_u2s_11_12({(~ in_u_rsc_merge_sva_rsp_1_rsp_0) , (~ in_u_rsc_merge_sva_rsp_1_rsp_1)
      , (~ return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm)})
      + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_10_e_dif1_acc_1_tmp = nl_return_add_generic_AC_RND_CONV_false_10_e_dif1_acc_1_tmp[11:0];
  assign nl_return_mult_generic_AC_RND_CONV_false_1_exp_acc_1_nl = conv_u2s_11_12({return_add_generic_AC_RND_CONV_false_5_e_r_qelse_qr_10_1_lpi_3_dfm_1
      , return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1}) + conv_s2s_11_12({10'b1000000000
      , (~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm)}) + 12'b000000000001;
  assign return_mult_generic_AC_RND_CONV_false_1_exp_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_1_exp_acc_1_nl[11:0];
  assign nl_return_mult_generic_AC_RND_CONV_false_1_exp_acc_tmp = conv_s2s_12_13(return_mult_generic_AC_RND_CONV_false_1_exp_acc_1_nl)
      + conv_u2s_11_13({operator_6_false_18_acc_psp_sva_10_0_rsp_0 , operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0
      , operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1}) + conv_u2s_1_13(return_extract_17_return_extract_17_nor_tmp);
  assign return_mult_generic_AC_RND_CONV_false_1_exp_acc_tmp = nl_return_mult_generic_AC_RND_CONV_false_1_exp_acc_tmp[12:0];
  assign return_extract_17_return_extract_17_or_sva_1 = (return_add_generic_AC_RND_CONV_false_5_e_r_qelse_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_5_res_rounded_lpi_3_dfm_51_0_1[51])
      & (~ return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_5_if_7_not_6_nl = ~ return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_5_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_5_if_7_not_6_nl);
  assign return_extract_17_return_extract_17_nor_tmp = ~((return_add_generic_AC_RND_CONV_false_5_e_r_qelse_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_9_op1_nan_sva_1 = operator_11_true_return_24_sva
      & (~ return_extract_1_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (z_out_49[10:1]), return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1));
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_1_nl = ~(MUX_v_10_2_2(10'b0000000000,
      z_out_12, return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1));
  assign return_add_generic_AC_RND_CONV_false_4_mux_18_nl = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_nl,
      return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_1_nl, z_out_47[53]);
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_qr_10_1_lpi_3_dfm_1 = ~(MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_4_mux_18_nl,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_4_e_r_qelse_or_svs_1));
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_2_nl = ~((z_out_49[0])
      & return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1);
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nor_nl = ~((z_out_14[0])
      | (~ return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1));
  assign return_add_generic_AC_RND_CONV_false_4_mux_19_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_2_nl,
      return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nor_nl, z_out_47[53]);
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1 = ~(return_add_generic_AC_RND_CONV_false_4_mux_19_nl
      | return_add_generic_AC_RND_CONV_false_4_e_r_qelse_or_svs_1);
  assign return_add_generic_AC_RND_CONV_false_4_m_r_51_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_4_res_rounded_lpi_3_dfm_51_0_1[51])
      & (~ return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_7_op1_nan_sva_1 = operator_11_true_return_1_sva
      & (~ return_extract_12_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_8_r_sign_mux_1_nl = MUX_s_1_2_2(stage_PE_1_tmp_im_d_1_lpi_3_dfm_51,
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_63, or_451_cse);
  assign nand_87_nl = ~(return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm , drf_qr_lval_14_smx_0_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1})));
  assign operator_11_true_return_15_sva_mx1 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_if_2_return_add_generic_AC_RND_CONV_false_8_if_2_and_1_mx2w0,
      return_add_generic_AC_RND_CONV_false_8_r_sign_mux_1_nl, nand_87_nl);
  assign return_add_generic_AC_RND_CONV_false_10_op1_nan_sva_1 = operator_11_true_return_26_sva
      & (~ return_extract_44_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1 = operator_11_true_return_1_sva
      & (~ return_extract_44_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_21_r_sign_mux_1_nl = MUX_s_1_2_2(stage_PE_1_tmp_re_d_1_lpi_3_dfm_63,
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_63, return_add_generic_AC_RND_CONV_false_21_op1_smaller_lor_lpi_3_dfm_2);
  assign nand_88_nl = ~(return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp
      & (({drf_qr_lval_14_smx_0_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm
      , return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1})));
  assign operator_11_true_return_15_sva_mx2 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_if_2_return_add_generic_AC_RND_CONV_false_7_if_2_and_1_mx1w0,
      return_add_generic_AC_RND_CONV_false_21_r_sign_mux_1_nl, nand_88_nl);
  assign return_add_generic_AC_RND_CONV_false_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_17,
      z_out_18, z_out_17[11]);
  assign return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1 = (stage_PE_1_tmp_im_d_1_sva_1_50_0[0])
      & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva;
  assign return_add_generic_AC_RND_CONV_false_op_smaller_qr_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm, and_dcpl_214);
  assign return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0 =
      MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_1_op2_mu_51_1_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0, and_dcpl_214);
  assign return_add_generic_AC_RND_CONV_false_op_smaller_qr_0_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1, and_dcpl_214);
  assign return_add_generic_AC_RND_CONV_false_e1_eq_e2_equal_tmp = (out_f_d_rsci_q_d[62:52])
      == (stage_PE_1_tmp_im_d_1_sva_1_63_51[11:1]);
  assign return_add_generic_AC_RND_CONV_false_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_40[54]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_40[53]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_40[52]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_40[51]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_40[50]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_40[49]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_40[48]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_40[47]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_40[46]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_40[45]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_40[44]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_40[43]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_40[42]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_40[41]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_40[40]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_40[39]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_40[38]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_40[37]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_40[36]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_40[35]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_40[34]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_40[33]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_40[32]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_40[31]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_40[30]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_40[29]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_40[28]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_40[27]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_40[26]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_40[25]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_40[24]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_40[23]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_40[22]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_40[21]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_40[20]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_40[19]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_40[18]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_40[17]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_40[16]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_40[15]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_40[14]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_40[13]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_40[12]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_40[11]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_40[10]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_40[9]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_40[8]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_40[7]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_40[6]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_40[5]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_40[4]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_40[3]))) | (return_add_generic_AC_RND_CONV_false_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_40[2])));
  assign return_add_generic_AC_RND_CONV_false_2_e_dif_qr_lpi_3_dfm_mx0_10_0 = MUX_v_11_2_2((z_out_17[10:0]),
      (z_out_18[10:0]), z_out_17[11]);
  assign return_add_generic_AC_RND_CONV_false_2_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_38[54]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_38[53]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_38[52]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_38[51]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_38[50]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_38[49]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_38[48]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_38[47]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_38[46]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_38[45]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_38[44]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_38[43]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_38[42]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_38[41]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_38[40]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_38[39]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_38[38]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_38[37]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_38[36]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_38[35]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_38[34]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_38[33]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_38[32]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_38[31]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_38[30]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_38[29]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_38[28]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_38[27]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_38[26]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_38[25]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_38[24]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_38[23]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_38[22]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_38[21]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_38[20]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_38[19]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_38[18]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_38[17]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_38[16]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_38[15]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_38[14]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_38[13]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_38[12]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_38[11]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_38[10]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_38[9]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_38[8]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_38[7]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_38[6]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_38[5]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_38[4]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_38[3]))) | (return_add_generic_AC_RND_CONV_false_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_38[2])));
  assign return_add_generic_AC_RND_CONV_false_2_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_2_e_dif_qr_lpi_3_dfm_mx0_10_0[10:6]!=5'b00000)
      | return_add_generic_AC_RND_CONV_false_1_e_dif_qelse_return_add_generic_AC_RND_CONV_false_1_e_dif_qelse_and_cse;
  assign return_add_generic_AC_RND_CONV_false_2_e_dif_sat_or_cse = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_2_e_dif_qr_lpi_3_dfm_mx0_10_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_2_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_e_dif_sat_or_cse = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (operator_33_true_10_acc_psp_1_sva_1[10:1]), return_add_generic_AC_RND_CONV_false_5_acc_2_itm_10_1));
  assign nl_operator_33_true_11_acc_nl = (z_out_13[10:1]) + 10'b0000000001;
  assign operator_33_true_11_acc_nl = nl_operator_33_true_11_acc_nl[9:0];
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_1_nl = ~(MUX_v_10_2_2(10'b0000000000,
      operator_33_true_11_acc_nl, return_add_generic_AC_RND_CONV_false_5_acc_2_itm_10_1));
  assign return_add_generic_AC_RND_CONV_false_5_mux_12_nl = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_nl,
      return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_1_nl, z_out_46[53]);
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qelse_qr_10_1_lpi_3_dfm_1 = ~(MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_5_mux_12_nl,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_5_e_r_qelse_or_svs_1));
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_2_nl = ~((operator_33_true_10_acc_psp_1_sva_1[0])
      & return_add_generic_AC_RND_CONV_false_5_acc_2_itm_10_1);
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nor_nl = ~((z_out_13[0])
      | (~ return_add_generic_AC_RND_CONV_false_5_acc_2_itm_10_1));
  assign return_add_generic_AC_RND_CONV_false_5_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_2_nl,
      return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nor_nl, z_out_46[53]);
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1 = ~(return_add_generic_AC_RND_CONV_false_5_mux_13_nl
      | return_add_generic_AC_RND_CONV_false_5_e_r_qelse_or_svs_1);
  assign return_add_generic_AC_RND_CONV_false_5_not_3_nl = ~ (z_out_46[53]);
  assign return_add_generic_AC_RND_CONV_false_5_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (z_out_46[51:0]), return_add_generic_AC_RND_CONV_false_5_not_3_nl);
  assign nl_operator_33_true_10_acc_psp_1_sva_1 = conv_s2s_7_12({operator_6_false_10_operator_6_false_10_conc_2_6_1
      , (~ (return_add_generic_AC_RND_CONV_false_20_ls_sva[0]))}) + conv_u2s_10_12({reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0
      , reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1});
  assign operator_33_true_10_acc_psp_1_sva_1 = nl_operator_33_true_10_acc_psp_1_sva_1[11:0];
  assign nl_return_add_generic_AC_RND_CONV_false_5_acc_2_nl =  -(operator_33_true_10_acc_psp_1_sva_1[10:0]);
  assign return_add_generic_AC_RND_CONV_false_5_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_5_acc_2_nl[10:0];
  assign return_add_generic_AC_RND_CONV_false_5_acc_2_itm_10_1 = readslicef_11_1_10(return_add_generic_AC_RND_CONV_false_5_acc_2_nl);
  assign return_add_generic_AC_RND_CONV_false_5_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_5_acc_2_itm_10_1
      | (~((operator_33_true_10_acc_psp_1_sva_1!=12'b000000000000)));
  assign return_add_generic_AC_RND_CONV_false_5_mux_9_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_5_acc_2_itm_10_1,
      return_add_generic_AC_RND_CONV_false_5_if_5_or_1_nl, z_out_46[53]);
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qelse_or_svs_1 = return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_5_mux_9_nl);
  assign return_add_generic_AC_RND_CONV_false_4_not_3_nl = ~ (z_out_47[53]);
  assign return_add_generic_AC_RND_CONV_false_4_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (z_out_47[51:0]), return_add_generic_AC_RND_CONV_false_4_not_3_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_4_acc_2_nl =  -(z_out_49[10:0]);
  assign return_add_generic_AC_RND_CONV_false_4_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_4_acc_2_nl[10:0];
  assign return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1 = readslicef_11_1_10(return_add_generic_AC_RND_CONV_false_4_acc_2_nl);
  assign return_add_generic_AC_RND_CONV_false_4_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1
      | (~((z_out_49!=12'b000000000000)));
  assign return_add_generic_AC_RND_CONV_false_4_mux_15_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1,
      return_add_generic_AC_RND_CONV_false_4_if_5_or_1_nl, z_out_47[53]);
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_or_svs_1 = return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_4_mux_15_nl);
  assign return_extract_27_return_extract_27_or_2_nl = (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_mx0w2!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx1 = MUX_s_1_2_2(return_extract_27_return_extract_27_or_2_nl,
      return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm_mx1, return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_8_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_8_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 | (return_extract_22_and_1_tmp
      & return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_15_do_sub_sva);
  assign and_357_nl = or_dcpl_597 & (~((z_out_46[53]) & return_add_generic_AC_RND_CONV_false_8_if_5_return_add_generic_AC_RND_CONV_false_8_if_5_and_tmp))
      & and_dcpl_300;
  assign return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm_mx1 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_5_res_rounded_lpi_3_dfm_51_0_1[51]),
      and_357_nl);
  assign return_add_generic_AC_RND_CONV_false_21_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_21_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_21_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_13_do_sub_sva);
  assign and_359_nl = or_dcpl_597 & (~(return_add_generic_AC_RND_CONV_false_21_if_5_return_add_generic_AC_RND_CONV_false_21_if_5_and_tmp
      & (return_add_generic_AC_RND_CONV_false_21_res_rounded_acc_tmp[53]))) & and_dcpl_300;
  assign return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm_mx2 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_21_res_rounded_lpi_3_dfm_51_0_1[51]),
      and_359_nl);
  assign return_add_generic_AC_RND_CONV_false_8_mux_16_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_and_10_9,
      (return_add_generic_AC_RND_CONV_false_8_exp_plus_1_12_1_lpi_3_dfm_1[9]), z_out_46[53]);
  assign return_add_generic_AC_RND_CONV_false_8_e_r_qelse_return_add_generic_AC_RND_CONV_false_8_e_r_qelse_and_nl
      = return_add_generic_AC_RND_CONV_false_8_mux_16_nl & (~ return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs_mx0w0);
  assign return_add_generic_AC_RND_CONV_false_8_mux_28_nl = MUX_v_9_2_2(return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_and_10_8_0,
      (return_add_generic_AC_RND_CONV_false_8_exp_plus_1_12_1_lpi_3_dfm_1[8:0]),
      z_out_46[53]);
  assign return_add_generic_AC_RND_CONV_false_8_e_r_qelse_not_3_nl = ~ return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs_mx0w0;
  assign return_add_generic_AC_RND_CONV_false_8_e_r_qelse_return_add_generic_AC_RND_CONV_false_8_e_r_qelse_and_2_nl
      = MUX_v_9_2_2(9'b000000000, return_add_generic_AC_RND_CONV_false_8_mux_28_nl,
      return_add_generic_AC_RND_CONV_false_8_e_r_qelse_not_3_nl);
  assign return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_mx0w2 = MUX_v_10_2_2(({return_add_generic_AC_RND_CONV_false_8_e_r_qelse_return_add_generic_AC_RND_CONV_false_8_e_r_qelse_and_nl
      , return_add_generic_AC_RND_CONV_false_8_e_r_qelse_return_add_generic_AC_RND_CONV_false_8_e_r_qelse_and_2_nl}),
      10'b1111111111, return_add_generic_AC_RND_CONV_false_8_exception_sva_1);
  assign return_extract_13_return_extract_13_return_extract_13_m_zero_not_6_nl =
      ~ return_extract_12_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_mx0w4_9_6
      = MUX_v_4_2_2(4'b0000, reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1, return_extract_13_return_extract_13_return_extract_13_m_zero_not_6_nl);
  assign return_extract_13_return_extract_13_return_extract_13_m_zero_not_5_nl =
      ~ return_extract_12_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_mx0w4_5_0
      = MUX_v_6_2_2(6'b000000, reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2, return_extract_13_return_extract_13_return_extract_13_m_zero_not_5_nl);
  assign return_add_generic_AC_RND_CONV_false_7_mux_21_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_and_11,
      return_add_generic_AC_RND_CONV_false_7_exp_plus_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_7_res_rounded_acc_tmp[53]);
  assign or_222_nl = or_dcpl_193 | and_dcpl_125 | operator_11_true_return_13_sva;
  assign return_add_generic_AC_RND_CONV_false_7_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs, or_222_nl);
  assign return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_7_mux_21_nl
      & (~ return_add_generic_AC_RND_CONV_false_7_e_r_qelse_mux_1_nl)) | return_add_generic_AC_RND_CONV_false_7_exception_sva_1;
  assign nl_operator_6_false_12_acc_nl = ({1'b1 , (~ (leading_sign_57_0_1_0_6_out_3[5:1]))})
      + 6'b000001;
  assign operator_6_false_12_acc_nl = nl_operator_6_false_12_acc_nl[5:0];
  assign nl_operator_33_true_12_acc_tmp = conv_s2s_7_13({operator_6_false_12_acc_nl
      , (~ (leading_sign_57_0_1_0_6_out_3[0]))}) + conv_u2s_11_13({drf_qr_lval_6_smx_lpi_3_dfm_mx0_10
      , drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_0});
  assign operator_33_true_12_acc_tmp = nl_operator_33_true_12_acc_tmp[12:0];
  assign return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm_mx1 = MUX_v_51_2_2((in_f_d_rsci_q_d[50:0]),
      (in_f_d_rsci_q_d[51:1]), return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp);
  assign return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0_mx2 =
      MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_mx0w4[50:1]),
      (return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_mx0w4[49:0]), return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_2_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_13_do_sub_sva);
  assign and_362_nl = (or_dcpl_158 | and_dcpl_112 | operator_11_true_return_24_sva
      | leading_sign_57_0_1_0_2_out_2) & inverse_lpi_1_dfm_1;
  assign and_365_nl = and_dcpl_281 & and_dcpl_294 & (~ leading_sign_57_0_1_0_2_out_2)
      & inverse_lpi_1_dfm_1;
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_51_mx0 = MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_2_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_1_res_rounded_lpi_3_dfm_51_0_1[51]),
      (stage_PE_1_tmp_im_d_1_sva_1_63_51[0]), {and_362_nl , and_365_nl , (~ inverse_lpi_1_dfm_1)});
  assign return_add_generic_AC_RND_CONV_false_2_if_7_return_add_generic_AC_RND_CONV_false_2_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_2_exception_sva_1 | leading_sign_57_0_1_0_2_out_2);
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0w0 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_1_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_2_if_7_return_add_generic_AC_RND_CONV_false_2_if_7_nor_nl);
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0 = MUX_v_51_2_2(stage_PE_1_tmp_im_d_1_sva_1_50_0,
      stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0w0, inverse_lpi_1_dfm_1);
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx1_50 = MUX_s_1_2_2((stage_PE_1_tmp_im_d_1_sva_1_50_0[50]),
      (stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0w0[50]), inverse_lpi_1_dfm_1);
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w0_10_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_1_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_2_exception_sva_1);
  assign or_206_nl = or_dcpl_158 | and_dcpl_112 | operator_11_true_return_24_sva;
  assign return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_3_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs, or_206_nl);
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w0_0 = (return_add_generic_AC_RND_CONV_false_1_mux_32
      & (~ return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_3_nl)) | return_add_generic_AC_RND_CONV_false_2_exception_sva_1;
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_1 = MUX_v_10_2_2((stage_PE_1_tmp_im_d_1_sva_1_63_51[11:2]),
      stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w0_10_1, inverse_lpi_1_dfm_1);
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0 = MUX_s_1_2_2((stage_PE_1_tmp_im_d_1_sva_1_63_51[1]),
      stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w0_0, inverse_lpi_1_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_op1_zero_sva_1 = operator_11_true_return_13_sva
      & return_extract_12_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_14_op2_nan_sva_1 = operator_11_true_return_13_sva
      & (~ return_extract_12_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_op1_nan_sva_1 = operator_11_true_return_24_sva
      & (~ return_extract_44_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_op2_nan_sva_1 = operator_11_true_return_1_sva
      & (~ return_extract_1_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_op1_inf_sva_1 = operator_11_true_return_24_sva
      & return_extract_44_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_op2_inf_sva_1 = operator_11_true_return_1_sva
      & return_extract_1_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_2_exception_sva_1 = return_add_generic_AC_RND_CONV_false_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_1_mux_16_cse;
  assign return_add_generic_AC_RND_CONV_false_exception_sva_1 = return_add_generic_AC_RND_CONV_false_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_3_mux_10_cse;
  assign return_add_generic_AC_RND_CONV_false_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_exception_sva_1
      | leading_sign_57_0_1_0_15_out_2;
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_1_if_acc_1_itm_12_1) | (z_out_54[105]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_if_not_nl = ~ (z_out_57[12]);
  assign return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      (z_out_57[11:0]), return_mult_generic_AC_RND_CONV_false_1_if_if_not_nl);
  assign return_mult_generic_AC_RND_CONV_false_1_e_incr_lpi_3_dfm_2 = ~((~(((z_out_54[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((z_out_54[51]) | return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_or_2))
      | (z_out_54[105]))) | (stage_u_add_3_acc_itm_rsp_1[12]));
  assign return_mult_generic_AC_RND_CONV_false_1_zero_m_return_mult_generic_AC_RND_CONV_false_1_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_1_r_zero_return_mult_generic_AC_RND_CONV_false_1_r_zero_nor_mdf_sva_1
      = ~(return_extract_16_and_tmp | return_extract_17_and_tmp);
  assign return_mult_generic_AC_RND_CONV_false_1_lor_lpi_3_dfm_1 = return_mult_generic_AC_RND_CONV_false_op1_zero_sva_1
      | return_extract_22_and_1_tmp | ((return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_1==12'b011111111110)
      & return_mult_generic_AC_RND_CONV_false_1_e_incr_lpi_3_dfm_2) | (z_out_55[11])
      | return_mult_generic_AC_RND_CONV_false_1_r_nan_sva_1;
  assign return_extract_22_and_1_tmp = operator_11_true_return_17_sva & return_extract_17_m_zero_sva;
  assign return_extract_16_and_tmp = return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_cse_sva
      & return_extract_12_m_zero_sva;
  assign return_extract_17_and_tmp = return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm
      & return_extract_17_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_mux_1_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_1_if_acc_1_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva, stage_u_add_3_acc_itm_rsp_1[12]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_mux_1_nl
      & (~ (z_out_54[105]));
  assign return_mult_generic_AC_RND_CONV_false_1_shift_right_conc_3_5 = (~ (stage_u_add_3_acc_itm_rsp_1[5]))
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm;
  assign return_mult_generic_AC_RND_CONV_false_1_shift_right_conc_3_0 = (~ (stage_u_add_3_acc_itm_rsp_1[0]))
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm;
  assign stage_d_mul_return_d_63_sva_1 = stage_PE_1_tmp_re_d_1_lpi_3_dfm_63 ^ return_add_generic_AC_RND_CONV_false_17_mux_6_itm;
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_63_mx1 = MUX_s_1_2_2((stage_PE_1_tmp_im_d_1_sva_1_63_51[12]),
      return_add_generic_AC_RND_CONV_false_12_mux_itm, inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_15_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_7_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_7_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_15_do_sub_sva);
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_51_mx1 = MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_15_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_3_res_rounded_lpi_3_dfm_51_0_1[51]),
      (stage_PE_1_tmp_im_d_1_sva_1_63_51[0]), {and_344_cse , and_347_cse , (~ inverse_lpi_1_dfm_1)});
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w2_10_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_15_exception_sva_1);
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_7_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs, or_dcpl_168);
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w2_0 = (return_add_generic_AC_RND_CONV_false_3_mux_26
      & (~ return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_7_nl)) | return_add_generic_AC_RND_CONV_false_15_exception_sva_1;
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx1_10_1 = MUX_v_10_2_2((stage_PE_1_tmp_im_d_1_sva_1_63_51[11:2]),
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w2_10_1, inverse_lpi_1_dfm_1);
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx1_0 = MUX_s_1_2_2((stage_PE_1_tmp_im_d_1_sva_1_63_51[1]),
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w2_0, inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp
      = (return_mult_generic_AC_RND_CONV_false_4_exp_1_11_0_lpi_3_dfm_3_10_0_1!=11'b00000000000);
  assign return_add_generic_AC_RND_CONV_false_24_if_5_return_add_generic_AC_RND_CONV_false_24_if_5_and_tmp
      = (return_add_generic_AC_RND_CONV_false_24_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_24_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_24_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_24_if_5_or_nl = return_add_generic_AC_RND_CONV_false_24_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_24_if_5_return_add_generic_AC_RND_CONV_false_24_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_24_mux_14_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_24_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_24_if_5_or_nl, return_add_generic_AC_RND_CONV_false_24_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_24_exception_sva_1 = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1 | return_add_generic_AC_RND_CONV_false_22_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_24_mux_14_nl;
  assign return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1 = operator_11_true_return_1_sva
      & return_extract_44_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_15_if_7_return_add_generic_AC_RND_CONV_false_15_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_15_exception_sva_1 | leading_sign_57_0_1_0_15_out_2);
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx0w2 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_3_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_15_if_7_return_add_generic_AC_RND_CONV_false_15_if_7_nor_nl);
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1 = MUX_v_51_2_2(stage_PE_1_tmp_im_d_1_sva_1_50_0,
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx0w2, inverse_lpi_1_dfm_1);
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx2_50 = MUX_s_1_2_2((stage_PE_1_tmp_im_d_1_sva_1_50_0[50]),
      (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx0w2[50]), inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_18_not_3_nl = ~ (return_add_generic_AC_RND_CONV_false_18_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_18_res_rounded_acc_tmp[51:0]), return_add_generic_AC_RND_CONV_false_18_not_3_nl);
  assign return_mult_generic_AC_RND_CONV_false_oelse_3_return_mult_generic_AC_RND_CONV_false_if_3_nor_nl
      = ~((~ return_mult_generic_AC_RND_CONV_false_zero_m_return_mult_generic_AC_RND_CONV_false_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_r_zero_return_mult_generic_AC_RND_CONV_false_r_zero_nor_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_lor_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (z_out[50:0]), return_mult_generic_AC_RND_CONV_false_oelse_3_return_mult_generic_AC_RND_CONV_false_if_3_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_6_op1_mu_0_lpi_3_dfm_1 = (stage_PE_1_tmp_im_d_1_sva_1_50_0[0])
      & (~ operator_11_true_return_13_sva);
  assign drf_qr_lval_6_smx_lpi_3_dfm_mx0_10 = MUX_s_1_2_2(operator_6_false_18_acc_psp_sva_10_0_rsp_0,
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0, and_dcpl_312);
  assign return_mult_generic_AC_RND_CONV_false_2_exp_mux_1_nl = MUX_v_9_2_2(operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0,
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0, and_dcpl_312);
  assign return_mult_generic_AC_RND_CONV_false_2_exp_mux_2_nl = MUX_s_1_2_2(operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1,
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1, and_dcpl_312);
  assign drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_0 = {return_mult_generic_AC_RND_CONV_false_2_exp_mux_1_nl
      , return_mult_generic_AC_RND_CONV_false_2_exp_mux_2_nl};
  assign return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm, return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50,
      and_dcpl_312);
  assign return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_50_mx0
      = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm, and_dcpl_312);
  assign return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0
      = MUX_v_50_2_2(reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1,
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0, and_dcpl_312);
  assign return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_0_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1, and_dcpl_312);
  assign nl_return_add_generic_AC_RND_CONV_false_19_ma1_lt_ma2_acc_2_nl = ({1'b1
      , stage_PE_1_tmp_re_d_1_lpi_3_dfm_51 , stage_PE_1_tmp_im_d_1_sva_1_50_0}) +
      conv_u2u_52_53({(~ stage_PE_1_tmp_im_d_1_lpi_3_dfm_51) , (~ stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0)})
      + 53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_19_ma1_lt_ma2_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_19_ma1_lt_ma2_acc_2_nl[52:0];
  assign return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_and_1_cse
      = (readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_19_ma1_lt_ma2_acc_2_nl))
      & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva;
  assign return_add_generic_AC_RND_CONV_false_19_op1_smaller_lor_lpi_3_dfm_2 = return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_and_1_cse
      | return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm;
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_2_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[49])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[52]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_3_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[48])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[51]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_4_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[47])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[50]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_5_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[46])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[49]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_6_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[45])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[48]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_7_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[44])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[47]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_8_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[43])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[46]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_9_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[42])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[45]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_10_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[41])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[44]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_11_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[40])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[43]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_12_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[39])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[42]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_13_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[38])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[41]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_14_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[37])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[40]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_15_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[36])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[39]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_16_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[35])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[38]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_17_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[34])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[37]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_18_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[33])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[36]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_19_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[32])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[35]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_20_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[31])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[34]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_21_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[30])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[33]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_22_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[29])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[32]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_23_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[28])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[31]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_24_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[27])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[30]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_25_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[26])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[29]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_26_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[25])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[28]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_27_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[24])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[27]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_28_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[23])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[26]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_29_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[22])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[25]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_30_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[21])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[24]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_31_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[20])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[23]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_32_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[19])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[22]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_33_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[18])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[21]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_34_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[17])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[20]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_35_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[16])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[19]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_36_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[15])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[18]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_37_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[14])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[17]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_38_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[13])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[16]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_39_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[12])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[15]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_40_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[11])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[14]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_41_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[10])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[13]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_42_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[9])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[12]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_43_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[8])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[11]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_44_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[7])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[10]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_45_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[6])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[9]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_46_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[5])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[8]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_47_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[4])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[7]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_48_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[3])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[6]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_49_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[2])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[5]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_50_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[1])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[4]));
  assign return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_51_cse = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[0])
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[3]));
  assign return_add_generic_AC_RND_CONV_false_6_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[54]))) | (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_50_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[53]))) | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_2_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_3_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_4_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_5_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_6_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_7_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_8_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_9_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_10_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_11_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_12_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_13_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_14_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_15_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_16_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_17_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_18_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_19_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_20_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_21_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_22_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_23_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_24_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_25_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_26_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_27_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_28_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_29_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_30_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_31_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_32_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_33_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_34_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_35_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_36_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_37_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_38_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_39_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_40_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_41_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_42_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_43_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_44_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_45_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_46_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_47_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_48_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_49_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_50_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_51_cse | (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[2])));
  assign return_mult_generic_AC_RND_CONV_false_if_1_aelse_return_mult_generic_AC_RND_CONV_false_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_3_if_acc_2_itm_12_1) | (return_mult_generic_AC_RND_CONV_false_3_p_sva_1[105]);
  assign return_mult_generic_AC_RND_CONV_false_if_if_not_1_nl = ~ (z_out_63[12]);
  assign return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_1_cse
      = MUX_v_12_2_2(12'b000000000000, (z_out_63[11:0]), return_mult_generic_AC_RND_CONV_false_if_if_not_1_nl);
  assign return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1 = ~((z_out_45[9:6]==4'b1111));
  assign return_mult_generic_AC_RND_CONV_false_3_e_incr_lpi_3_dfm_2 = ~((~(((return_mult_generic_AC_RND_CONV_false_3_p_sva_1[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((return_mult_generic_AC_RND_CONV_false_3_p_sva_1[51]) | return_mult_generic_AC_RND_CONV_false_if_1_aelse_return_mult_generic_AC_RND_CONV_false_if_1_aelse_or_2))
      | (return_mult_generic_AC_RND_CONV_false_3_p_sva_1[105]))) | (z_out_45[12]));
  assign return_mult_generic_AC_RND_CONV_false_zero_m_return_mult_generic_AC_RND_CONV_false_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_r_zero_return_mult_generic_AC_RND_CONV_false_r_zero_nor_mdf_sva_1
      = ~(return_mult_generic_AC_RND_CONV_false_op1_zero_sva_1 | return_mult_generic_AC_RND_CONV_false_op2_zero_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_1_and_3_nl = (return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_2[0])
      & return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm;
  assign nl_r_rnd_dummy_1_51_0_sva_1 = ({return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_1
      , (return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_2[50:1])}) +
      conv_u2u_1_52(return_mult_generic_AC_RND_CONV_false_1_and_3_nl);
  assign r_rnd_dummy_1_51_0_sva_1 = nl_r_rnd_dummy_1_51_0_sva_1[51:0];
  assign return_mult_generic_AC_RND_CONV_false_r_nan_sva_1 = return_add_generic_AC_RND_CONV_false_7_op1_nan_sva_1
      | (operator_11_true_return_15_sva & (~ return_extract_15_m_zero_sva)) | (return_add_generic_AC_RND_CONV_false_7_op1_inf_sva_1
      & return_mult_generic_AC_RND_CONV_false_op2_zero_sva_1) | (return_mult_generic_AC_RND_CONV_false_op1_zero_sva_1
      & return_mult_generic_AC_RND_CONV_false_op2_inf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_3_exp_ovf_lor_lpi_3_dfm_2 = return_mult_generic_AC_RND_CONV_false_3_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_3_exp_ovf_oif_aelse_and_1_tmp
      | (z_out_55[11]);
  assign return_mult_generic_AC_RND_CONV_false_lor_lpi_3_dfm_1 = return_add_generic_AC_RND_CONV_false_7_op1_inf_sva_1
      | return_mult_generic_AC_RND_CONV_false_op2_inf_sva_1 | return_mult_generic_AC_RND_CONV_false_3_exp_ovf_lor_lpi_3_dfm_2
      | return_mult_generic_AC_RND_CONV_false_r_nan_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_return_mult_generic_AC_RND_CONV_false_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_if_1_and_1_tmp_1 | (z_out_45[12]));
  assign return_mult_generic_AC_RND_CONV_false_and_2_nl = return_mult_generic_AC_RND_CONV_false_if_1_and_1_tmp_1
      & (~ (z_out_45[12]));
  assign return_mult_generic_AC_RND_CONV_false_res_bef_rnd_3_53_1_lpi_3_dfm_1 = MUX1HOT_v_53_3_2((return_mult_generic_AC_RND_CONV_false_3_p_sva_1[104:52]),
      (return_mult_generic_AC_RND_CONV_false_3_p_sva_1[103:51]), (z_out_35[53:1]),
      {return_mult_generic_AC_RND_CONV_false_return_mult_generic_AC_RND_CONV_false_nor_nl
      , return_mult_generic_AC_RND_CONV_false_and_2_nl , (z_out_45[12])});
  assign return_mult_generic_AC_RND_CONV_false_op2_inf_sva_1 = operator_11_true_return_15_sva
      & return_extract_15_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_op2_zero_sva_1 = return_extract_15_return_extract_15_nor_cse_sva
      & return_extract_15_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_1_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_3_if_acc_2_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva, z_out_45[12]);
  assign return_mult_generic_AC_RND_CONV_false_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_1_nl
      & (~ (return_mult_generic_AC_RND_CONV_false_3_p_sva_1[105]));
  assign nl_operator_6_false_13_acc_psp_sva_1 = conv_u2s_11_12({drf_qr_lval_6_smx_lpi_3_dfm_mx0_10
      , drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_0}) + conv_s2s_7_12({1'b1 , (~ leading_sign_57_0_1_0_6_out_3)})
      + 12'b000000000001;
  assign operator_6_false_13_acc_psp_sva_1 = nl_operator_6_false_13_acc_psp_sva_1[11:0];
  assign return_add_generic_AC_RND_CONV_false_6_e_dif_sat_or_2_nl = (z_out_19[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_19_e_dif_sat_sva_1 = MUX_v_6_2_2((z_out_19[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_6_e_dif_sat_or_2_nl);
  assign return_mult_generic_AC_RND_CONV_false_if_or_3_cse = (~ (z_out_45[5])) |
      return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_3_if_not_1_nl = ~ return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_if_nand_1_cse = ~(MUX_v_4_2_2(4'b0000,
      (z_out_45[4:1]), return_mult_generic_AC_RND_CONV_false_3_if_not_1_nl));
  assign return_mult_generic_AC_RND_CONV_false_if_or_cse = (~ (z_out_45[0])) | return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_4_oelse_3_return_mult_generic_AC_RND_CONV_false_4_if_3_nor_nl
      = ~((~ return_mult_generic_AC_RND_CONV_false_4_zero_m_return_mult_generic_AC_RND_CONV_false_4_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_4_r_zero_return_mult_generic_AC_RND_CONV_false_4_r_zero_nor_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_4_lor_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (r_rnd_dummy_4_51_0_sva_1[50:0]), return_mult_generic_AC_RND_CONV_false_4_oelse_3_return_mult_generic_AC_RND_CONV_false_4_if_3_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_6_res_rounded_and_1_nl = (return_add_generic_AC_RND_CONV_false_6_res_rounded_asn_rndc_sva_1[3])
      & ((return_add_generic_AC_RND_CONV_false_6_res_rounded_asn_rndc_sva_1[0]) |
      (return_add_generic_AC_RND_CONV_false_6_res_rounded_asn_rndc_sva_1[1]) | (return_add_generic_AC_RND_CONV_false_6_res_rounded_asn_rndc_sva_1[2])
      | (return_add_generic_AC_RND_CONV_false_6_res_rounded_asn_rndc_sva_1[4]));
  assign nl_return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp = conv_u2u_53_54(return_add_generic_AC_RND_CONV_false_6_res_rounded_asn_rndc_sva_1[56:4])
      + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_6_res_rounded_and_1_nl);
  assign return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp = nl_return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[53:0];
  assign return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_2_if_acc_1_itm_12_1) | (return_mult_generic_AC_RND_CONV_false_2_p_sva_1[105]);
  assign return_mult_generic_AC_RND_CONV_false_2_if_if_not_nl = ~ (operator_6_false_16_acc_psp_sva_1[12]);
  assign return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      (operator_6_false_16_acc_psp_sva_1[11:0]), return_mult_generic_AC_RND_CONV_false_2_if_if_not_nl);
  assign return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1 = ({return_extract_41_return_extract_41_or_1_cse_sva
      , (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[51:0])}) * ({return_extract_19_return_extract_19_or_sva_1
      , return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1});
  assign nl_return_mult_generic_AC_RND_CONV_false_2_exp_acc_1_nl = conv_u2u_11_12({return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1_9_1
      , return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1_0 , return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1})
      + conv_u2u_1_12(~ return_extract_41_return_extract_41_or_1_cse_sva) + 12'b000000000001;
  assign return_mult_generic_AC_RND_CONV_false_2_exp_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_2_exp_acc_1_nl[11:0];
  assign nl_return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp = conv_u2s_12_13(return_mult_generic_AC_RND_CONV_false_2_exp_acc_1_nl)
      + conv_s2s_11_13({1'b1 , (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[61:52])}) + conv_u2s_1_13(return_extract_19_return_extract_19_nor_tmp);
  assign return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp = nl_return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp[12:0];
  assign nl_operator_6_false_16_acc_psp_sva_1 = return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp
      + conv_s2s_7_13({1'b1 , (~ leading_sign_53_0_2_out_1)}) + 13'b0000000000001;
  assign operator_6_false_16_acc_psp_sva_1 = nl_operator_6_false_16_acc_psp_sva_1[12:0];
  assign return_mult_generic_AC_RND_CONV_false_2_if_nor_ovfl_sva_1 = ~((return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp[9:6]==4'b1111));
  assign return_mult_generic_AC_RND_CONV_false_2_e_incr_lpi_3_dfm_2 = ~((~(((return_mult_generic_AC_RND_CONV_false_2_p_sva_1[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((return_mult_generic_AC_RND_CONV_false_2_p_sva_1[51]) | return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_or_2))
      | (return_mult_generic_AC_RND_CONV_false_2_p_sva_1[105]))) | (return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp[12]));
  assign return_mult_generic_AC_RND_CONV_false_2_zero_m_return_mult_generic_AC_RND_CONV_false_2_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_2_r_zero_return_mult_generic_AC_RND_CONV_false_2_r_zero_nor_mdf_sva_1
      = ~(return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 | (return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp
      & return_extract_19_return_extract_19_nor_tmp));
  assign return_mult_generic_AC_RND_CONV_false_2_op2_inf_sva_1 = operator_11_true_19_operator_11_true_19_and_tmp
      & return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp;
  assign return_extract_19_return_extract_19_nor_tmp = ~((return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1_9_1!=9'b000000000)
      | return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1_0 | return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1);
  assign return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp = ~(return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_mux_1_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_2_if_acc_1_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva, return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp[12]);
  assign return_mult_generic_AC_RND_CONV_false_2_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_mux_1_nl
      & (~ (return_mult_generic_AC_RND_CONV_false_2_p_sva_1[105]));
  assign return_extract_19_return_extract_19_or_sva_1 = (return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1_9_1!=9'b000000000)
      | return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1_0 | return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_6_r_nan_or_1_nl = operator_11_true_return_15_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | (operator_11_true_return_13_sva
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva & return_add_generic_AC_RND_CONV_false_13_do_sub_sva);
  assign and_369_nl = and_dcpl_121 & and_dcpl_314;
  assign return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_6_res_rounded_lpi_3_dfm_51_0_1[51]),
      and_369_nl);
  assign return_add_generic_AC_RND_CONV_false_6_if_7_return_add_generic_AC_RND_CONV_false_6_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_6_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_6_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_6_if_7_return_add_generic_AC_RND_CONV_false_6_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_6_mux_18_nl = MUX_v_9_2_2((return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_and_9[9:1]),
      operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0, return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_not_6_nl = ~ return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1;
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_return_add_generic_AC_RND_CONV_false_6_e_r_qelse_and_nl
      = MUX_v_9_2_2(9'b000000000, return_add_generic_AC_RND_CONV_false_6_mux_18_nl,
      return_add_generic_AC_RND_CONV_false_6_e_r_qelse_not_6_nl);
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1_9_1 = MUX_v_9_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_return_add_generic_AC_RND_CONV_false_6_e_r_qelse_and_nl,
      9'b111111111, return_add_generic_AC_RND_CONV_false_6_exception_sva_1);
  assign return_add_generic_AC_RND_CONV_false_6_mux_35_nl = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_and_9[0]),
      operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1, return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1_0 = (return_add_generic_AC_RND_CONV_false_6_mux_35_nl
      & (~ return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1)) | return_add_generic_AC_RND_CONV_false_6_exception_sva_1;
  assign and_178_cse = ((stage_u_add_3_acc_itm_rsp_1[11]) | (~ return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva;
  assign return_add_generic_AC_RND_CONV_false_6_mux_19_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_and_11,
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm,
      return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[53]);
  assign or_214_nl = and_178_cse | or_dcpl_25 | or_dcpl_183 | (return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm
      & (return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[53]));
  assign return_add_generic_AC_RND_CONV_false_19_e_r_qelse_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs, or_214_nl);
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_6_mux_19_nl
      & (~ return_add_generic_AC_RND_CONV_false_19_e_r_qelse_mux_nl)) | return_add_generic_AC_RND_CONV_false_6_exception_sva_1;
  assign operator_11_true_19_operator_11_true_19_and_tmp = (return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1_9_1==9'b111111111)
      & return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1_0 & return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_6_not_4_nl = ~ (return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_6_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[51:0]), return_add_generic_AC_RND_CONV_false_6_not_4_nl);
  assign return_add_generic_AC_RND_CONV_false_6_if_5_or_nl = and_178_cse | return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm;
  assign return_add_generic_AC_RND_CONV_false_6_mux_16_nl = MUX_s_1_2_2(and_178_cse,
      return_add_generic_AC_RND_CONV_false_6_if_5_or_nl, return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_6_exception_sva_1 = operator_11_true_return_13_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | operator_11_true_return_15_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_6_mux_16_nl;
  assign return_mult_generic_AC_RND_CONV_false_2_shift_right_conc_3_5 = (~ (return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp[5]))
      | return_mult_generic_AC_RND_CONV_false_2_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_2_if_not_nl = ~ return_mult_generic_AC_RND_CONV_false_2_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_2_shift_right_conc_3_4_1 = ~(MUX_v_4_2_2(4'b0000,
      (return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp[4:1]), return_mult_generic_AC_RND_CONV_false_2_if_not_nl));
  assign return_mult_generic_AC_RND_CONV_false_2_shift_right_conc_3_0 = (~ (return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp[0]))
      | return_mult_generic_AC_RND_CONV_false_2_if_nor_ovfl_sva_1;
  assign nl_return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp = ({1'b1 , reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd
      , reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1 , reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2})
      + conv_u2s_11_12(~ return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1)
      + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp = nl_return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp[11:0];
  assign nl_return_add_generic_AC_RND_CONV_false_7_e_dif_qif_acc_1_nl = ({1'b1 ,
      return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1}) + conv_u2s_11_12({(~
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd) , (~ reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1)
      , (~ reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2)}) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_7_e_dif_qif_acc_1_nl = nl_return_add_generic_AC_RND_CONV_false_7_e_dif_qif_acc_1_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_7_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp,
      return_add_generic_AC_RND_CONV_false_7_e_dif_qif_acc_1_nl, return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp[11]);
  assign return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1 =
      MUX_v_11_2_2(({operator_6_false_18_acc_psp_sva_10_0_rsp_0 , operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0
      , operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1}), 11'b11111111111, operator_11_true_return_13_sva);
  assign return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1 = (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm[0])
      & return_add_generic_AC_RND_CONV_false_11_mux_itm;
  assign return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1 = BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx1
      | return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0 = MUX_s_1_2_2((return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1[50]),
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx1, return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp);
  assign return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0 = MUX_v_50_2_2((return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1[49:0]),
      (return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1[50:1]), return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp);
  assign return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1 = (return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1[0])
      & return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1,
      and_dcpl_248);
  assign return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_51_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0,
      and_dcpl_248);
  assign return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2(reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_248);
  assign return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_0_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_248);
  assign return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp = ({reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd
      , reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1 , reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2})
      == (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1);
  assign nl_return_add_generic_AC_RND_CONV_false_7_ma1_lt_ma2_acc_1_nl = ({1'b1 ,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm , return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm})
      + conv_u2u_52_53({(~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx1)
      , (~ return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1)}) + 53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_7_ma1_lt_ma2_acc_1_nl = nl_return_add_generic_AC_RND_CONV_false_7_ma1_lt_ma2_acc_1_nl[52:0];
  assign return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_and_cse
      = (readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_7_ma1_lt_ma2_acc_1_nl))
      & return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_7_op1_smaller_lor_lpi_3_dfm_2 = return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp[11]);
  assign return_add_generic_AC_RND_CONV_false_7_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[54]))) | (return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[53]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[52]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[51]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[50]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[49]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[48]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[47]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[46]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[45]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[44]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[43]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[42]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[41]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[40]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[39]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[38]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[37]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[36]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[35]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[34]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[33]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[32]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[31]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[30]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[29]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[28]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[27]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[26]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[25]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[24]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[23]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[22]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[21]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[20]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[19]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[18]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[17]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[16]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[15]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[14]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[13]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[12]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[11]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[10]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[9]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[8]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[7]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[6]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[5]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[4]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[3]))) | (return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_7_lshift_itm[2])));
  assign nl_return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp = ({1'b1 , BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0})
      + conv_u2s_11_12(~ return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1)
      + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp = nl_return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp[11:0];
  assign nl_return_add_generic_AC_RND_CONV_false_8_e_dif_qif_acc_1_nl = ({1'b1 ,
      return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1}) + conv_u2s_11_12(~
      BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_8_e_dif_qif_acc_1_nl = nl_return_add_generic_AC_RND_CONV_false_8_e_dif_qif_acc_1_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_8_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp,
      return_add_generic_AC_RND_CONV_false_8_e_dif_qif_acc_1_nl, return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp[11]);
  assign return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[0])
      & return_add_generic_AC_RND_CONV_false_21_unequal_tmp;
  assign return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1,
      and_dcpl_220);
  assign return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_51_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(drf_qr_lval_14_smx_0_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0,
      and_dcpl_220);
  assign return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_220);
  assign return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_0_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_220);
  assign return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp = (BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0)
      == (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1);
  assign return_add_generic_AC_RND_CONV_false_8_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_37[54]))) | (return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (z_out_37[53]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_37[52]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_37[51]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_37[50]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_37[49]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_37[48]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_37[47]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_37[46]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_37[45]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_37[44]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_37[43]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_37[42]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_37[41]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_37[40]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_37[39]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_37[38]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_37[37]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_37[36]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_37[35]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_37[34]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_37[33]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_37[32]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_37[31]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_37[30]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_37[29]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_37[28]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_37[27]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_37[26]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_37[25]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_37[24]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_37[23]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_37[22]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_37[21]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_37[20]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_37[19]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_37[18]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_37[17]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_37[16]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_37[15]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_37[14]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_37[13]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_37[12]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_37[11]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_37[10]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_37[9]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_37[8]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_37[7]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_37[6]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_37[5]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_37[4]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_37[3]))) | (return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_37[2])));
  assign return_add_generic_AC_RND_CONV_false_8_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_8_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_8_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_8_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_7_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_7_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_7_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_7_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp
      = (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1!=11'b00000000000);
  assign return_add_generic_AC_RND_CONV_false_7_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      operator_33_true_15_acc_2, return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_7_res_rounded_and_nl = (return_add_generic_AC_RND_CONV_false_7_res_rounded_asn_rndc_sva_1[3])
      & ((return_add_generic_AC_RND_CONV_false_7_res_rounded_asn_rndc_sva_1[0]) |
      (return_add_generic_AC_RND_CONV_false_7_res_rounded_asn_rndc_sva_1[1]) | (return_add_generic_AC_RND_CONV_false_7_res_rounded_asn_rndc_sva_1[2])
      | (return_add_generic_AC_RND_CONV_false_7_res_rounded_asn_rndc_sva_1[4]));
  assign nl_return_add_generic_AC_RND_CONV_false_7_res_rounded_acc_tmp = conv_u2u_53_54(return_add_generic_AC_RND_CONV_false_7_res_rounded_asn_rndc_sva_1[56:4])
      + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_7_res_rounded_and_nl);
  assign return_add_generic_AC_RND_CONV_false_7_res_rounded_acc_tmp = nl_return_add_generic_AC_RND_CONV_false_7_res_rounded_acc_tmp[53:0];
  assign return_add_generic_AC_RND_CONV_false_7_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_7_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_7_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_12_mux_itm);
  assign and_373_nl = or_dcpl_625 & (~(return_add_generic_AC_RND_CONV_false_20_if_5_return_add_generic_AC_RND_CONV_false_20_if_5_and_1_tmp
      & (return_add_generic_AC_RND_CONV_false_7_res_rounded_acc_tmp[53]))) & and_dcpl_316;
  assign return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_7_res_rounded_lpi_3_dfm_51_0_1[51]),
      and_373_nl);
  assign return_add_generic_AC_RND_CONV_false_7_not_3_nl = ~ (return_add_generic_AC_RND_CONV_false_7_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_7_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_7_res_rounded_acc_tmp[51:0]), return_add_generic_AC_RND_CONV_false_7_not_3_nl);
  assign nl_operator_33_true_17_acc_nl = conv_s2s_11_12(z_out_49[11:1]) + 12'b000000000001;
  assign operator_33_true_17_acc_nl = nl_operator_33_true_17_acc_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_8_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      operator_33_true_17_acc_nl, return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_8_op1_nan_sva_1 = operator_11_true_return_17_sva
      & (~ return_extract_17_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_7_if_7_return_add_generic_AC_RND_CONV_false_7_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_7_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_7_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_7_if_7_return_add_generic_AC_RND_CONV_false_7_if_7_nor_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_9_e_dif_qif_acc_1_nl = ({1'b1 ,
      return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1})
      + conv_u2s_11_12(~ (stage_PE_1_x_re_d_sva[62:52])) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_9_e_dif_qif_acc_1_nl = nl_return_add_generic_AC_RND_CONV_false_9_e_dif_qif_acc_1_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_9_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(return_add_generic_AC_RND_CONV_false_9_e_dif1_acc_1_tmp,
      return_add_generic_AC_RND_CONV_false_9_e_dif_qif_acc_1_nl, return_add_generic_AC_RND_CONV_false_9_e_dif1_acc_1_tmp[11]);
  assign return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1 = (stage_PE_1_x_re_d_sva[0])
      & return_add_generic_AC_RND_CONV_false_22_unequal_tmp;
  assign return_extract_25_return_extract_25_or_2_nl = (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_extract_25_return_extract_25_or_2_nl,
      return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1[50]), return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0 = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1[50:1]),
      (return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1[49:0]), return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1[0])
      & (~ return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_9_e1_eq_e2_equal_tmp = (stage_PE_1_x_re_d_sva[62:52])
      == ({return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1});
  assign return_add_generic_AC_RND_CONV_false_9_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_mux_cse
      & (~ (z_out_40[54]))) | (return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_cse
      & (~ (z_out_40[53]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[49])
      & (~ (z_out_40[52]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[48])
      & (~ (z_out_40[51]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[47])
      & (~ (z_out_40[50]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[46])
      & (~ (z_out_40[49]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[45])
      & (~ (z_out_40[48]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[44])
      & (~ (z_out_40[47]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[43])
      & (~ (z_out_40[46]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[42])
      & (~ (z_out_40[45]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[41])
      & (~ (z_out_40[44]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[40])
      & (~ (z_out_40[43]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[39])
      & (~ (z_out_40[42]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[38])
      & (~ (z_out_40[41]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[37])
      & (~ (z_out_40[40]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[36])
      & (~ (z_out_40[39]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[35])
      & (~ (z_out_40[38]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[34])
      & (~ (z_out_40[37]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[33])
      & (~ (z_out_40[36]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[32])
      & (~ (z_out_40[35]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[31])
      & (~ (z_out_40[34]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[30])
      & (~ (z_out_40[33]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[29])
      & (~ (z_out_40[32]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[28])
      & (~ (z_out_40[31]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[27])
      & (~ (z_out_40[30]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[26])
      & (~ (z_out_40[29]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[25])
      & (~ (z_out_40[28]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[24])
      & (~ (z_out_40[27]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[23])
      & (~ (z_out_40[26]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[22])
      & (~ (z_out_40[25]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[21])
      & (~ (z_out_40[24]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[20])
      & (~ (z_out_40[23]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[19])
      & (~ (z_out_40[22]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[18])
      & (~ (z_out_40[21]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[17])
      & (~ (z_out_40[20]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[16])
      & (~ (z_out_40[19]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[15])
      & (~ (z_out_40[18]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[14])
      & (~ (z_out_40[17]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[13])
      & (~ (z_out_40[16]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[12])
      & (~ (z_out_40[15]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[11])
      & (~ (z_out_40[14]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[10])
      & (~ (z_out_40[13]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[9])
      & (~ (z_out_40[12]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[8])
      & (~ (z_out_40[11]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[7])
      & (~ (z_out_40[10]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[6])
      & (~ (z_out_40[9]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[5])
      & (~ (z_out_40[8]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[4])
      & (~ (z_out_40[7]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[3])
      & (~ (z_out_40[6]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[2])
      & (~ (z_out_40[5]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[1])
      & (~ (z_out_40[4]))) | ((return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1[0])
      & (~ (z_out_40[3]))) | (return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_2_cse
      & (~ (z_out_40[2])));
  assign nl_return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0w1 = ({1'b1
      , (stage_PE_1_x_im_d_sva[62:52])}) + conv_u2s_11_12({(~ return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_mx0w2)
      , (~ return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1)}) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0w1 = nl_return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0w1[11:0];
  assign nl_return_add_generic_AC_RND_CONV_false_10_e_dif_qif_acc_1_nl = ({1'b1 ,
      return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_mx0w2 , return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1})
      + conv_u2s_11_12(~ (stage_PE_1_x_im_d_sva[62:52])) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_10_e_dif_qif_acc_1_nl = nl_return_add_generic_AC_RND_CONV_false_10_e_dif_qif_acc_1_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0w1,
      return_add_generic_AC_RND_CONV_false_10_e_dif_qif_acc_1_nl, return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0w1[11]);
  assign return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp
      = ~((return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_mx0w2!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_9_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_9_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_9_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp
      = ~((return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_8_if_5_return_add_generic_AC_RND_CONV_false_8_if_5_and_tmp
      = (return_add_generic_AC_RND_CONV_false_8_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_8_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_8_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_8_if_5_or_nl = return_add_generic_AC_RND_CONV_false_8_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_8_if_5_return_add_generic_AC_RND_CONV_false_8_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_8_mux_14_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_8_if_5_or_nl, z_out_46[53]);
  assign return_add_generic_AC_RND_CONV_false_8_exception_sva_1 = return_extract_22_and_1_tmp
      | return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_8_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_8_mux_14_nl;
  assign return_add_generic_AC_RND_CONV_false_8_exp_plus_1_0_lpi_3_dfm_1 = (z_out_49[0])
      | (~ return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_8_r_inf_lpi_3_dfm_2 = ((reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_2_1[0])
      | (~ return_add_generic_AC_RND_CONV_false_21_else_4_return_add_generic_AC_RND_CONV_false_21_else_4_nand_tmp))
      & return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_8_mux_8_itm = MUX_v_6_2_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[5:0]),
      return_add_generic_AC_RND_CONV_false_20_ls_sva, return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_7_if_5_or_cse = return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_20_if_5_return_add_generic_AC_RND_CONV_false_20_if_5_and_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_7_mux_18_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_7_if_5_or_cse, return_add_generic_AC_RND_CONV_false_7_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_7_exception_sva_1 = return_add_generic_AC_RND_CONV_false_7_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_7_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_7_mux_18_nl;
  assign return_add_generic_AC_RND_CONV_false_7_exp_plus_1_0_lpi_3_dfm_1 = operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1
      | (~ return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2 = ((stage_u_add_3_acc_itm_rsp_1[11])
      | (~ return_add_generic_AC_RND_CONV_false_10_else_4_return_add_generic_AC_RND_CONV_false_10_else_4_nand_tmp))
      & return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1;
  assign nl_operator_33_true_44_acc_tmp = conv_s2s_7_13({operator_6_false_2_operator_6_false_2_conc_2_6_1
      , (~ (leading_sign_57_0_1_0_2_out_3[0]))}) + conv_u2s_11_13({reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1
      , reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2 , drf_qr_lval_12_smx_0_lpi_3_dfm});
  assign operator_33_true_44_acc_tmp = nl_operator_33_true_44_acc_tmp[12:0];
  assign return_add_generic_AC_RND_CONV_false_9_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      z_out_21, return_add_generic_AC_RND_CONV_false_22_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_10_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_1_cse
      & (~ (z_out_39[54]))) | (return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_cse
      & (~ (z_out_39[53]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[49])
      & (~ (z_out_39[52]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[48])
      & (~ (z_out_39[51]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[47])
      & (~ (z_out_39[50]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[46])
      & (~ (z_out_39[49]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[45])
      & (~ (z_out_39[48]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[44])
      & (~ (z_out_39[47]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[43])
      & (~ (z_out_39[46]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[42])
      & (~ (z_out_39[45]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[41])
      & (~ (z_out_39[44]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[40])
      & (~ (z_out_39[43]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[39])
      & (~ (z_out_39[42]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[38])
      & (~ (z_out_39[41]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[37])
      & (~ (z_out_39[40]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[36])
      & (~ (z_out_39[39]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[35])
      & (~ (z_out_39[38]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[34])
      & (~ (z_out_39[37]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[33])
      & (~ (z_out_39[36]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[32])
      & (~ (z_out_39[35]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[31])
      & (~ (z_out_39[34]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[30])
      & (~ (z_out_39[33]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[29])
      & (~ (z_out_39[32]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[28])
      & (~ (z_out_39[31]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[27])
      & (~ (z_out_39[30]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[26])
      & (~ (z_out_39[29]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[25])
      & (~ (z_out_39[28]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[24])
      & (~ (z_out_39[27]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[23])
      & (~ (z_out_39[26]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[22])
      & (~ (z_out_39[25]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[21])
      & (~ (z_out_39[24]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[20])
      & (~ (z_out_39[23]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[19])
      & (~ (z_out_39[22]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[18])
      & (~ (z_out_39[21]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[17])
      & (~ (z_out_39[20]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[16])
      & (~ (z_out_39[19]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[15])
      & (~ (z_out_39[18]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[14])
      & (~ (z_out_39[17]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[13])
      & (~ (z_out_39[16]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[12])
      & (~ (z_out_39[15]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[11])
      & (~ (z_out_39[14]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[10])
      & (~ (z_out_39[13]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[9])
      & (~ (z_out_39[12]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[8])
      & (~ (z_out_39[11]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[7])
      & (~ (z_out_39[10]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[6])
      & (~ (z_out_39[9]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[5])
      & (~ (z_out_39[8]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[4])
      & (~ (z_out_39[7]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[3])
      & (~ (z_out_39[6]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[2])
      & (~ (z_out_39[5]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[1])
      & (~ (z_out_39[4]))) | ((return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse[0])
      & (~ (z_out_39[3]))) | (return_add_generic_AC_RND_CONV_false_14_op1_mu_mux_1_cse
      & (~ (z_out_39[2])));
  assign nl_return_add_generic_AC_RND_CONV_false_11_e_dif_qif_acc_1_sdt = ({1'b1
      , return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_itm
      , return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm})
      + conv_u2s_11_12(~ (stage_PE_1_x_re_d_sva[62:52])) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_11_e_dif_qif_acc_1_sdt = nl_return_add_generic_AC_RND_CONV_false_11_e_dif_qif_acc_1_sdt[11:0];
  assign return_add_generic_AC_RND_CONV_false_11_e_dif_qr_lpi_3_dfm_mx0_9_1 = MUX_v_9_2_2(operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0,
      (return_add_generic_AC_RND_CONV_false_11_e_dif_qif_acc_1_sdt[9:1]), operator_6_false_18_acc_psp_sva_11);
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_return_add_generic_AC_RND_CONV_false_11_sticky_bit_return_add_generic_AC_RND_CONV_false_11_sticky_bit_or_cse
      = (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm & (~
      (z_out_43[54]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm
      & (~ (z_out_43[53]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[49])
      & (~ (z_out_43[52]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[48])
      & (~ (z_out_43[51]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[47])
      & (~ (z_out_43[50]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[46])
      & (~ (z_out_43[49]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[45])
      & (~ (z_out_43[48]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[44])
      & (~ (z_out_43[47]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[43])
      & (~ (z_out_43[46]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[42])
      & (~ (z_out_43[45]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[41])
      & (~ (z_out_43[44]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[40])
      & (~ (z_out_43[43]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[39])
      & (~ (z_out_43[42]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[38])
      & (~ (z_out_43[41]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[37])
      & (~ (z_out_43[40]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[36])
      & (~ (z_out_43[39]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[35])
      & (~ (z_out_43[38]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[34])
      & (~ (z_out_43[37]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[33])
      & (~ (z_out_43[36]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[32])
      & (~ (z_out_43[35]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[31])
      & (~ (z_out_43[34]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[30])
      & (~ (z_out_43[33]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[29])
      & (~ (z_out_43[32]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[28])
      & (~ (z_out_43[31]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[27])
      & (~ (z_out_43[30]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[26])
      & (~ (z_out_43[29]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[25])
      & (~ (z_out_43[28]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[24])
      & (~ (z_out_43[27]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[23])
      & (~ (z_out_43[26]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[22])
      & (~ (z_out_43[25]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[21])
      & (~ (z_out_43[24]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[20])
      & (~ (z_out_43[23]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[19])
      & (~ (z_out_43[22]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[18])
      & (~ (z_out_43[21]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[17])
      & (~ (z_out_43[20]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[16])
      & (~ (z_out_43[19]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[15])
      & (~ (z_out_43[18]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[14])
      & (~ (z_out_43[17]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[13])
      & (~ (z_out_43[16]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[12])
      & (~ (z_out_43[15]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[11])
      & (~ (z_out_43[14]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[10])
      & (~ (z_out_43[13]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[9])
      & (~ (z_out_43[12]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[8])
      & (~ (z_out_43[11]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[7])
      & (~ (z_out_43[10]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[6])
      & (~ (z_out_43[9]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[5])
      & (~ (z_out_43[8]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[4])
      & (~ (z_out_43[7]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[3])
      & (~ (z_out_43[6]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[2])
      & (~ (z_out_43[5]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[1])
      & (~ (z_out_43[4]))) | ((return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm[0])
      & (~ (z_out_43[3]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm
      & (~ (z_out_43[2])));
  assign return_add_generic_AC_RND_CONV_false_11_e_dif_qelse_mux_nl = MUX_s_1_2_2(operator_6_false_18_acc_psp_sva_10_0_rsp_0,
      (return_add_generic_AC_RND_CONV_false_11_e_dif_qif_acc_1_sdt[10]), operator_6_false_18_acc_psp_sva_11);
  assign return_add_generic_AC_RND_CONV_false_11_e_dif_sat_or_1_seb = (return_add_generic_AC_RND_CONV_false_11_e_dif_qr_lpi_3_dfm_mx0_9_1[8:5]!=4'b0000)
      | return_add_generic_AC_RND_CONV_false_11_e_dif_qelse_mux_nl | ((return_add_generic_AC_RND_CONV_false_11_e_dif_qif_acc_1_sdt[11])
      & operator_6_false_18_acc_psp_sva_11);
  assign return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1_5_1 = MUX_v_5_2_2((return_add_generic_AC_RND_CONV_false_11_e_dif_qr_lpi_3_dfm_mx0_9_1[4:0]),
      5'b11111, return_add_generic_AC_RND_CONV_false_11_e_dif_sat_or_1_seb);
  assign return_add_generic_AC_RND_CONV_false_11_e_dif_qelse_mux_2_nl = MUX_s_1_2_2(operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1,
      (return_add_generic_AC_RND_CONV_false_11_e_dif_qif_acc_1_sdt[0]), operator_6_false_18_acc_psp_sva_11);
  assign return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1_0 = return_add_generic_AC_RND_CONV_false_11_e_dif_qelse_mux_2_nl
      | return_add_generic_AC_RND_CONV_false_11_e_dif_sat_or_1_seb;
  assign return_add_generic_AC_RND_CONV_false_9_if_5_or_nl = return_add_generic_AC_RND_CONV_false_9_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_22_if_5_return_add_generic_AC_RND_CONV_false_22_if_5_and_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_9_mux_17_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_9_if_5_or_nl, z_out_47[53]);
  assign return_add_generic_AC_RND_CONV_false_9_exception_sva_1 = return_add_generic_AC_RND_CONV_false_9_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op1_inf_sva_1 | return_add_generic_AC_RND_CONV_false_9_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op1_nan_sva_1 | return_add_generic_AC_RND_CONV_false_9_mux_17_cse;
  assign return_add_generic_AC_RND_CONV_false_9_exp_plus_1_0_lpi_3_dfm_1 = (z_out_51[0])
      | (~ return_add_generic_AC_RND_CONV_false_22_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_9_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_9_exception_sva_1
      | leading_sign_57_0_1_0_2_out_2;
  assign return_add_generic_AC_RND_CONV_false_9_r_inf_lpi_3_dfm_2 = ((operator_33_true_44_acc_tmp[11])
      | ((operator_33_true_44_acc_tmp[10:0]==11'b11111111111))) & return_add_generic_AC_RND_CONV_false_22_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_10_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      z_out_56, return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_10_if_5_return_add_generic_AC_RND_CONV_false_10_if_5_and_tmp
      = (return_add_generic_AC_RND_CONV_false_10_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_10_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_10_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_10_if_5_or_nl = return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_10_if_5_return_add_generic_AC_RND_CONV_false_10_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_10_mux_17_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_10_if_5_or_nl, z_out_46[53]);
  assign return_add_generic_AC_RND_CONV_false_10_exception_sva_1 = return_add_generic_AC_RND_CONV_false_10_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_10_mux_17_cse;
  assign return_add_generic_AC_RND_CONV_false_10_exp_plus_1_0_lpi_3_dfm_1 = (z_out_13[0])
      | (~ return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_10_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_10_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_11_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      z_out_56, return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva);
  assign nl_return_add_generic_AC_RND_CONV_false_12_e_dif_qif_acc_1_sdt = ({1'b1
      , in_u_rsc_merge_sva_rsp_1_rsp_0 , in_u_rsc_merge_sva_rsp_1_rsp_1 , return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm})
      + conv_u2s_11_12(~ (stage_PE_1_x_im_d_sva[62:52])) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_12_e_dif_qif_acc_1_sdt = nl_return_add_generic_AC_RND_CONV_false_12_e_dif_qif_acc_1_sdt[11:0];
  assign return_add_generic_AC_RND_CONV_false_12_e_dif_qr_lpi_3_dfm_mx0_9_1 = MUX_v_9_2_2(operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0,
      (return_add_generic_AC_RND_CONV_false_12_e_dif_qif_acc_1_sdt[9:1]), operator_6_false_18_acc_psp_sva_11);
  assign return_add_generic_AC_RND_CONV_false_12_e_dif_qelse_mux_nl = MUX_s_1_2_2(operator_6_false_18_acc_psp_sva_10_0_rsp_0,
      (return_add_generic_AC_RND_CONV_false_12_e_dif_qif_acc_1_sdt[10]), operator_6_false_18_acc_psp_sva_11);
  assign return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_1_seb = (return_add_generic_AC_RND_CONV_false_12_e_dif_qr_lpi_3_dfm_mx0_9_1[8:5]!=4'b0000)
      | return_add_generic_AC_RND_CONV_false_12_e_dif_qelse_mux_nl | ((return_add_generic_AC_RND_CONV_false_12_e_dif_qif_acc_1_sdt[11])
      & operator_6_false_18_acc_psp_sva_11);
  assign return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1_5_1 = MUX_v_5_2_2((return_add_generic_AC_RND_CONV_false_12_e_dif_qr_lpi_3_dfm_mx0_9_1[4:0]),
      5'b11111, return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_1_seb);
  assign return_add_generic_AC_RND_CONV_false_12_e_dif_qelse_mux_2_nl = MUX_s_1_2_2(operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1,
      (return_add_generic_AC_RND_CONV_false_12_e_dif_qif_acc_1_sdt[0]), operator_6_false_18_acc_psp_sva_11);
  assign return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1_0 = return_add_generic_AC_RND_CONV_false_12_e_dif_qelse_mux_2_nl
      | return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_1_seb;
  assign return_add_generic_AC_RND_CONV_false_11_if_5_return_add_generic_AC_RND_CONV_false_11_if_5_and_tmp
      = (return_add_generic_AC_RND_CONV_false_11_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_11_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_11_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_11_if_5_or_nl = return_add_generic_AC_RND_CONV_false_11_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_11_if_5_return_add_generic_AC_RND_CONV_false_11_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_11_mux_10_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_11_if_5_or_nl, z_out_46[53]);
  assign return_add_generic_AC_RND_CONV_false_11_exception_sva_1 = operator_11_true_return_1_sva
      | operator_11_true_return_24_sva | operator_11_true_return_17_sva | return_add_generic_AC_RND_CONV_false_15_do_sub_sva
      | return_add_generic_AC_RND_CONV_false_11_mux_10_nl;
  assign return_add_generic_AC_RND_CONV_false_11_exp_plus_1_0_lpi_3_dfm_1 = (z_out_13[0])
      | (~ return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva);
  assign return_add_generic_AC_RND_CONV_false_11_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_11_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_11_r_inf_lpi_3_dfm_2 = ((stage_u_add_3_acc_itm_rsp_1[11])
      | (~ return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva;
  assign return_add_generic_AC_RND_CONV_false_12_exception_sva_1 = operator_11_true_return_13_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | operator_11_true_return_15_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_10_mux_17_cse;
  assign return_add_generic_AC_RND_CONV_false_12_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_12_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1 = (in_f_d_rsci_q_d[0])
      & return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm_1,
      and_dcpl_215);
  assign return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0
      = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0, return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm_mx1,
      and_dcpl_215);
  assign return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1,
      and_dcpl_215);
  assign return_add_generic_AC_RND_CONV_false_14_e1_eq_e2_equal_tmp = (stage_PE_1_x_im_d_sva[62:52])
      == (in_f_d_rsci_q_d[62:52]);
  assign return_add_generic_AC_RND_CONV_false_14_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_40[54]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_40[53]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_40[52]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_40[51]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_40[50]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_40[49]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_40[48]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_40[47]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_40[46]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_40[45]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_40[44]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_40[43]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_40[42]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_40[41]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_40[40]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_40[39]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_40[38]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_40[37]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_40[36]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_40[35]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_40[34]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_40[33]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_40[32]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_40[31]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_40[30]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_40[29]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_40[28]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_40[27]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_40[26]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_40[25]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_40[24]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_40[23]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_40[22]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_40[21]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_40[20]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_40[19]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_40[18]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_40[17]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_40[16]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_40[15]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_40[14]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_40[13]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_40[12]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_40[11]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_40[10]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_40[9]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_40[8]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_40[7]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_40[6]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_40[5]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_40[4]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_40[3]))) | (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_40[2])));
  assign return_add_generic_AC_RND_CONV_false_16_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_38[54]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_38[53]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_38[52]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_38[51]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_38[50]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_38[49]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_38[48]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_38[47]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_38[46]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_38[45]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_38[44]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_38[43]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_38[42]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_38[41]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_38[40]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_38[39]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_38[38]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_38[37]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_38[36]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_38[35]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_38[34]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_38[33]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_38[32]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_38[31]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_38[30]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_38[29]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_38[28]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_38[27]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_38[26]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_38[25]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_38[24]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_38[23]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_38[22]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_38[21]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_38[20]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_38[19]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_38[18]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_38[17]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_38[16]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_38[15]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_38[14]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_38[13]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_38[12]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_38[11]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_38[10]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_38[9]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_38[8]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_38[7]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_38[6]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_38[5]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_38[4]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_38[3]))) | (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_38[2])));
  assign return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0
      = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_4_op1_mu_51_1_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_4_op2_mu_51_1_lpi_3_dfm_mx0, and_dcpl_225);
  assign return_add_generic_AC_RND_CONV_false_18_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_4_op_bigger_mux_3_cse
      & (~ (z_out_42[54]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_42[53]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_42[52]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_42[51]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_42[50]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_42[49]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_42[48]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_42[47]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_42[46]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_42[45]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_42[44]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_42[43]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_42[42]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_42[41]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_42[40]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_42[39]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_42[38]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_42[37]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_42[36]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_42[35]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_42[34]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_42[33]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_42[32]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_42[31]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_42[30]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_42[29]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_42[28]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_42[27]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_42[26]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_42[25]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_42[24]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_42[23]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_42[22]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_42[21]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_42[20]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_42[19]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_42[18]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_42[17]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_42[16]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_42[15]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_42[14]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_42[13]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_42[12]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_42[11]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_42[10]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_42[9]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_42[8]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_42[7]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_42[6]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_42[5]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_42[4]))) | ((return_add_generic_AC_RND_CONV_false_17_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_42[3]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_42[2])));
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_1 = MUX_v_10_2_2((stage_PE_1_tmp_im_d_1_sva_1_63_51[11:2]),
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w4_10_1, inverse_lpi_1_dfm_1);
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0 = MUX_s_1_2_2((stage_PE_1_tmp_im_d_1_sva_1_63_51[1]),
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w4_0, inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_17_not_3_nl = ~ (return_add_generic_AC_RND_CONV_false_17_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_17_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_17_res_rounded_acc_tmp[51:0]), return_add_generic_AC_RND_CONV_false_17_not_3_nl);
  assign return_add_generic_AC_RND_CONV_false_16_exception_sva_1 = return_add_generic_AC_RND_CONV_false_14_op1_inf_sva_1
      | return_mult_generic_AC_RND_CONV_false_op1_zero_sva_1 | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_3_mux_10_cse;
  assign return_add_generic_AC_RND_CONV_false_14_exception_sva_1 = return_add_generic_AC_RND_CONV_false_14_op1_inf_sva_1
      | return_mult_generic_AC_RND_CONV_false_op1_zero_sva_1 | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_1_mux_16_cse;
  assign nl_operator_6_false_39_acc_nl = ({1'b1 , (~ (leading_sign_57_0_1_0_18_out_3[5:1]))})
      + 6'b000001;
  assign operator_6_false_39_acc_nl = nl_operator_6_false_39_acc_nl[5:0];
  assign nl_operator_33_true_36_acc_psp_1_sva_1 = conv_s2s_7_12({operator_6_false_39_acc_nl
      , (~ (leading_sign_57_0_1_0_18_out_3[0]))}) + conv_u2s_10_12({reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1
      , reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2});
  assign operator_33_true_36_acc_psp_1_sva_1 = nl_operator_33_true_36_acc_psp_1_sva_1[11:0];
  assign nl_return_add_generic_AC_RND_CONV_false_18_acc_2_nl =  -(operator_33_true_36_acc_psp_1_sva_1[10:0]);
  assign return_add_generic_AC_RND_CONV_false_18_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_18_acc_2_nl[10:0];
  assign return_add_generic_AC_RND_CONV_false_18_acc_2_itm_10 = readslicef_11_1_10(return_add_generic_AC_RND_CONV_false_18_acc_2_nl);
  assign nl_operator_6_false_40_acc_psp_1_sva_1 = conv_u2s_10_11({reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1
      , reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2}) + conv_s2s_7_11({1'b1 , (~ leading_sign_57_0_1_0_18_out_3)})
      + 11'b00000000001;
  assign operator_6_false_40_acc_psp_1_sva_1 = nl_operator_6_false_40_acc_psp_1_sva_1[10:0];
  assign return_add_generic_AC_RND_CONV_false_18_res_rounded_and_cse = (z_out_38[3])
      & ((z_out_38[0]) | (z_out_38[1]) | (z_out_38[2]) | (z_out_38[4]));
  assign nl_return_add_generic_AC_RND_CONV_false_18_res_rounded_acc_tmp = conv_u2u_53_54(z_out_38[56:4])
      + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_18_res_rounded_and_cse);
  assign return_add_generic_AC_RND_CONV_false_18_res_rounded_acc_tmp = nl_return_add_generic_AC_RND_CONV_false_18_res_rounded_acc_tmp[53:0];
  assign return_add_generic_AC_RND_CONV_false_18_mux_4_itm = MUX_v_6_2_2(reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2,
      leading_sign_57_0_1_0_18_out_3, return_add_generic_AC_RND_CONV_false_18_acc_2_itm_10);
  assign nl_operator_6_false_37_acc_nl = ({1'b1 , (~ (leading_sign_57_0_1_0_17_out_3[5:1]))})
      + 6'b000001;
  assign operator_6_false_37_acc_nl = nl_operator_6_false_37_acc_nl[5:0];
  assign nl_operator_33_true_34_acc_psp_1_sva_1 = conv_s2s_7_12({operator_6_false_37_acc_nl
      , (~ (leading_sign_57_0_1_0_17_out_3[0]))}) + conv_u2s_10_12({reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1
      , reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2});
  assign operator_33_true_34_acc_psp_1_sva_1 = nl_operator_33_true_34_acc_psp_1_sva_1[11:0];
  assign nl_return_add_generic_AC_RND_CONV_false_17_acc_2_nl =  -(operator_33_true_34_acc_psp_1_sva_1[10:0]);
  assign return_add_generic_AC_RND_CONV_false_17_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_17_acc_2_nl[10:0];
  assign return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10 = readslicef_11_1_10(return_add_generic_AC_RND_CONV_false_17_acc_2_nl);
  assign return_add_generic_AC_RND_CONV_false_17_res_rounded_and_nl = (return_add_generic_AC_RND_CONV_false_17_res_rounded_asn_rndc_sva_1[3])
      & ((return_add_generic_AC_RND_CONV_false_17_res_rounded_asn_rndc_sva_1[0])
      | (return_add_generic_AC_RND_CONV_false_17_res_rounded_asn_rndc_sva_1[1]) |
      (return_add_generic_AC_RND_CONV_false_17_res_rounded_asn_rndc_sva_1[2]) | (return_add_generic_AC_RND_CONV_false_17_res_rounded_asn_rndc_sva_1[4]));
  assign nl_return_add_generic_AC_RND_CONV_false_17_res_rounded_acc_tmp = conv_u2u_53_54(return_add_generic_AC_RND_CONV_false_17_res_rounded_asn_rndc_sva_1[56:4])
      + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_17_res_rounded_and_nl);
  assign return_add_generic_AC_RND_CONV_false_17_res_rounded_acc_tmp = nl_return_add_generic_AC_RND_CONV_false_17_res_rounded_acc_tmp[53:0];
  assign nl_operator_32_false_1_acc_nl = (~ (BUTTERFLY_1_else_2_tmp2_1_sva[3:0]))
      + ({(BUTTERFLY_1_else_2_tmp2_1_sva[1:0]) , 2'b01});
  assign operator_32_false_1_acc_nl = nl_operator_32_false_1_acc_nl[3:0];
  assign nl_operator_32_false_1_mul_atp_sva_1 = ({operator_32_false_1_acc_nl , 12'b000000000001})
      + (~ (BUTTERFLY_1_else_2_tmp2_1_sva[15:0]));
  assign operator_32_false_1_mul_atp_sva_1 = nl_operator_32_false_1_mul_atp_sva_1[15:0];
  assign return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm, and_dcpl_224);
  assign return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0
      = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm_mx1,
      return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0, and_dcpl_224);
  assign return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1,
      and_dcpl_224);
  assign return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp = (in_f_d_rsci_q_d[62:52])
      == (stage_PE_1_tmp_im_d_1_sva_1_63_51[11:1]);
  assign return_add_generic_AC_RND_CONV_false_13_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_40[54]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_40[53]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_40[52]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_40[51]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_40[50]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_40[49]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_40[48]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_40[47]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_40[46]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_40[45]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_40[44]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_40[43]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_40[42]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_40[41]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_40[40]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_40[39]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_40[38]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_40[37]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_40[36]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_40[35]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_40[34]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_40[33]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_40[32]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_40[31]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_40[30]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_40[29]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_40[28]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_40[27]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_40[26]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_40[25]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_40[24]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_40[23]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_40[22]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_40[21]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_40[20]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_40[19]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_40[18]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_40[17]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_40[16]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_40[15]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_40[14]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_40[13]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_40[12]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_40[11]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_40[10]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_40[9]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_40[8]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_40[7]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_40[6]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_40[5]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_40[4]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_40[3]))) | (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_40[2])));
  assign return_add_generic_AC_RND_CONV_false_15_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_38[54]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_38[53]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_38[52]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_38[51]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_38[50]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_38[49]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_38[48]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_38[47]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_38[46]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_38[45]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_38[44]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_38[43]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_38[42]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_38[41]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_38[40]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_38[39]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_38[38]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_38[37]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_38[36]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_38[35]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_38[34]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_38[33]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_38[32]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_38[31]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_38[30]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_38[29]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_38[28]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_38[27]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_38[26]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_38[25]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_38[24]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_38[23]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_38[22]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_38[21]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_38[20]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_38[19]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_38[18]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_38[17]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_38[16]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_38[15]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_38[14]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_38[13]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_38[12]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_38[11]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_38[10]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_38[9]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_38[8]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_38[7]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_38[6]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_38[5]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_38[4]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_38[3]))) | (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_38[2])));
  assign return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_4_if_acc_1_itm_12_1) | (z_out_54[105]);
  assign return_mult_generic_AC_RND_CONV_false_4_e_incr_lpi_3_dfm_2 = ~((~(((z_out_54[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((z_out_54[51]) | return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_or_2))
      | (z_out_54[105]))) | (z_out_45[12]));
  assign return_mult_generic_AC_RND_CONV_false_4_zero_m_return_mult_generic_AC_RND_CONV_false_4_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_4_r_zero_return_mult_generic_AC_RND_CONV_false_4_r_zero_nor_mdf_sva_1
      = ~(return_mult_generic_AC_RND_CONV_false_4_op1_zero_sva_1 | return_mult_generic_AC_RND_CONV_false_4_op2_zero_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_4_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_4_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_4_else_1_sticky_bit_or_cse
      = ((z_out_26[105]) & (~ (z_out_41[52]))) | ((z_out_26[104]) & (~ (z_out_41[51])))
      | ((z_out_26[103]) & (~ (z_out_41[50]))) | ((z_out_26[102]) & (~ (z_out_41[49])))
      | ((z_out_26[101]) & (~ (z_out_41[48]))) | ((z_out_26[100]) & (~ (z_out_41[47])))
      | ((z_out_26[99]) & (~ (z_out_41[46]))) | ((z_out_26[98]) & (~ (z_out_41[45])))
      | ((z_out_26[97]) & (~ (z_out_41[44]))) | ((z_out_26[96]) & (~ (z_out_41[43])))
      | ((z_out_26[95]) & (~ (z_out_41[42]))) | ((z_out_26[94]) & (~ (z_out_41[41])))
      | ((z_out_26[93]) & (~ (z_out_41[40]))) | ((z_out_26[92]) & (~ (z_out_41[39])))
      | ((z_out_26[91]) & (~ (z_out_41[38]))) | ((z_out_26[90]) & (~ (z_out_41[37])))
      | ((z_out_26[89]) & (~ (z_out_41[36]))) | ((z_out_26[88]) & (~ (z_out_41[35])))
      | ((z_out_26[87]) & (~ (z_out_41[34]))) | ((z_out_26[86]) & (~ (z_out_41[33])))
      | ((z_out_26[85]) & (~ (z_out_41[32]))) | ((z_out_26[84]) & (~ (z_out_41[31])))
      | ((z_out_26[83]) & (~ (z_out_41[30]))) | ((z_out_26[82]) & (~ (z_out_41[29])))
      | ((z_out_26[81]) & (~ (z_out_41[28]))) | ((z_out_26[80]) & (~ (z_out_41[27])))
      | ((z_out_26[79]) & (~ (z_out_41[26]))) | ((z_out_26[78]) & (~ (z_out_41[25])))
      | ((z_out_26[77]) & (~ (z_out_41[24]))) | ((z_out_26[76]) & (~ (z_out_41[23])))
      | ((z_out_26[75]) & (~ (z_out_41[22]))) | ((z_out_26[74]) & (~ (z_out_41[21])))
      | ((z_out_26[73]) & (~ (z_out_41[20]))) | ((z_out_26[72]) & (~ (z_out_41[19])))
      | ((z_out_26[71]) & (~ (z_out_41[18]))) | ((z_out_26[70]) & (~ (z_out_41[17])))
      | ((z_out_26[69]) & (~ (z_out_41[16]))) | ((z_out_26[68]) & (~ (z_out_41[15])))
      | ((z_out_26[67]) & (~ (z_out_41[14]))) | ((z_out_26[66]) & (~ (z_out_41[13])))
      | ((z_out_26[65]) & (~ (z_out_41[12]))) | ((z_out_26[64]) & (~ (z_out_41[11])))
      | ((z_out_26[63]) & (~ (z_out_41[10]))) | ((z_out_26[62]) & (~ (z_out_41[9])))
      | ((z_out_26[61]) & (~ (z_out_41[8]))) | ((z_out_26[60]) & (~ (z_out_41[7])))
      | ((z_out_26[59]) & (~ (z_out_41[6]))) | ((z_out_26[58]) & (~ (z_out_41[5])))
      | ((z_out_26[57]) & (~ (z_out_41[4]))) | ((z_out_26[56]) & (~ (z_out_41[3])))
      | ((z_out_26[55]) & (~ (z_out_41[2]))) | ((z_out_26[54]) & (~ (z_out_41[1])))
      | ((z_out_26[53]) & (~ (z_out_41[0]))) | (z_out_26[52:0]!=53'b00000000000000000000000000000000000000000000000000000);
  assign return_mult_generic_AC_RND_CONV_false_4_if_1_or_nl = (z_out_54[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_or_2
      & (z_out_54[51]));
  assign return_mult_generic_AC_RND_CONV_false_4_mux_13_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_4_if_1_or_nl,
      return_mult_generic_AC_RND_CONV_false_4_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_4_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_4_else_1_sticky_bit_or_cse,
      z_out_45[12]);
  assign return_mult_generic_AC_RND_CONV_false_4_and_nl = (return_mult_generic_AC_RND_CONV_false_4_res_bef_rnd_3_53_1_lpi_3_dfm_1[0])
      & (return_mult_generic_AC_RND_CONV_false_4_mux_13_nl | (return_mult_generic_AC_RND_CONV_false_4_res_bef_rnd_3_53_1_lpi_3_dfm_1[1]));
  assign nl_r_rnd_dummy_4_51_0_sva_1 = (return_mult_generic_AC_RND_CONV_false_4_res_bef_rnd_3_53_1_lpi_3_dfm_1[52:1])
      + conv_u2u_1_52(return_mult_generic_AC_RND_CONV_false_4_and_nl);
  assign r_rnd_dummy_4_51_0_sva_1 = nl_r_rnd_dummy_4_51_0_sva_1[51:0];
  assign return_mult_generic_AC_RND_CONV_false_4_r_nan_sva_1 = return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1
      | (operator_11_true_49_operator_11_true_49_and_tmp & (~ return_extract_49_m_zero_return_extract_49_m_zero_nor_tmp))
      | (return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1 & return_mult_generic_AC_RND_CONV_false_4_op2_zero_sva_1)
      | (return_mult_generic_AC_RND_CONV_false_4_op1_zero_sva_1 & return_mult_generic_AC_RND_CONV_false_4_op2_inf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_4_exp_ovf_oif_aelse_nor_cse = ~((return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_1_cse[11])
      | (return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_1_cse[0]));
  assign return_mult_generic_AC_RND_CONV_false_4_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_4_exp_ovf_oif_aelse_and_tmp
      = (return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_1_cse[10:1]==10'b1111111111)
      & return_mult_generic_AC_RND_CONV_false_4_exp_ovf_oif_aelse_nor_cse & return_mult_generic_AC_RND_CONV_false_4_e_incr_lpi_3_dfm_2;
  assign return_mult_generic_AC_RND_CONV_false_4_lor_lpi_3_dfm_1 = return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1
      | return_mult_generic_AC_RND_CONV_false_4_op2_inf_sva_1 | return_mult_generic_AC_RND_CONV_false_4_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_4_exp_ovf_oif_aelse_and_tmp
      | (z_out_55[11]) | return_mult_generic_AC_RND_CONV_false_4_r_nan_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_4_return_mult_generic_AC_RND_CONV_false_4_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_4_if_1_and_1_tmp_1 | (z_out_45[12]));
  assign return_mult_generic_AC_RND_CONV_false_4_and_2_nl = return_mult_generic_AC_RND_CONV_false_4_if_1_and_1_tmp_1
      & (~ (z_out_45[12]));
  assign return_mult_generic_AC_RND_CONV_false_4_res_bef_rnd_3_53_1_lpi_3_dfm_1 =
      MUX1HOT_v_53_3_2((z_out_54[104:52]), (z_out_54[103:51]), (z_out_35[53:1]),
      {return_mult_generic_AC_RND_CONV_false_4_return_mult_generic_AC_RND_CONV_false_4_nor_nl
      , return_mult_generic_AC_RND_CONV_false_4_and_2_nl , (z_out_45[12])});
  assign return_mult_generic_AC_RND_CONV_false_4_op2_inf_sva_1 = operator_11_true_49_operator_11_true_49_and_tmp
      & return_extract_49_m_zero_return_extract_49_m_zero_nor_tmp;
  assign return_mult_generic_AC_RND_CONV_false_4_op1_zero_sva_1 = return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_cse_sva
      & return_extract_44_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_4_op2_zero_sva_1 = return_extract_49_return_extract_49_nor_tmp
      & return_extract_49_m_zero_return_extract_49_m_zero_nor_tmp;
  assign return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_mux_1_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_4_if_acc_1_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva, z_out_45[12]);
  assign return_mult_generic_AC_RND_CONV_false_4_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_mux_1_nl
      & (~ (z_out_54[105]));
  assign return_extract_49_return_extract_49_or_sva_1 = (return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1_9_1!=9'b000000000)
      | return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1_0 | return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm;
  assign return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_50 = reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd
      & (~ return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_4_if_7_not_7_nl = ~ return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0 = MUX_v_50_2_2(50'b00000000000000000000000000000000000000000000000000,
      reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1,
      return_add_generic_AC_RND_CONV_false_4_if_7_not_7_nl);
  assign return_extract_2_return_extract_2_return_extract_2_m_zero_not_7_nl = ~ return_extract_17_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1_9_1 = MUX_v_9_2_2(9'b000000000,
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0, return_extract_2_return_extract_2_return_extract_2_m_zero_not_7_nl);
  assign return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1_0 = reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1
      & (~ return_extract_17_m_zero_sva);
  assign return_extract_49_return_extract_49_nor_tmp = ~((return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1_9_1!=9'b000000000)
      | return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1_0 | return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm);
  assign operator_11_true_49_operator_11_true_49_and_tmp = (return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1_9_1==9'b111111111)
      & return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1_0 & return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm;
  assign return_extract_49_m_zero_return_extract_49_m_zero_nor_tmp = ~(drf_qr_lval_14_smx_0_lpi_3_dfm
      | return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_50 | (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0!=50'b00000000000000000000000000000000000000000000000000));
  assign nl_stage_u_add_9_acc_psp_sva_1 = conv_u2s_16_18({reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd
      , reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_2_1 , reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0
      , reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0 , reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1})
      - conv_s2s_17_18(z_out_58);
  assign stage_u_add_9_acc_psp_sva_1 = nl_stage_u_add_9_acc_psp_sva_1[17:0];
  assign return_add_generic_AC_RND_CONV_false_15_exception_sva_1 = return_add_generic_AC_RND_CONV_false_7_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_7_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_3_mux_10_cse;
  assign return_add_generic_AC_RND_CONV_false_13_exception_sva_1 = return_add_generic_AC_RND_CONV_false_7_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_7_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_1_mux_16_cse;
  assign return_add_generic_AC_RND_CONV_false_13_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_13_exception_sva_1
      | leading_sign_57_0_1_0_2_out_2;
  assign return_add_generic_AC_RND_CONV_false_19_op1_mu_0_lpi_3_dfm_1 = (stage_PE_1_tmp_im_d_1_sva_1_50_0[0])
      & (~ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_cse_sva);
  assign return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm,
      and_dcpl_312);
  assign return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_50_mx0
      = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50, and_dcpl_312);
  assign return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_19_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm,
      and_dcpl_312);
  assign return_add_generic_AC_RND_CONV_false_19_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[54]))) | (return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_50_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[53]))) | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_2_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_3_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_4_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_5_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_6_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_7_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_8_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_9_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_10_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_11_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_12_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_13_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_14_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_15_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_16_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_17_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_18_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_19_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_20_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_21_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_22_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_23_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_24_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_25_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_26_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_27_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_28_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_29_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_30_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_31_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_32_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_33_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_34_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_35_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_36_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_37_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_38_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_39_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_40_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_41_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_42_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_43_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_44_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_45_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_46_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_47_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_48_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_49_cse | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_50_cse
      | return_add_generic_AC_RND_CONV_false_6_sticky_bit_and_51_cse | (return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_19_lshift_1_itm[2])));
  assign return_mult_generic_AC_RND_CONV_false_3_zero_m_return_mult_generic_AC_RND_CONV_false_3_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_3_r_zero_return_mult_generic_AC_RND_CONV_false_3_r_zero_nor_mdf_sva_1
      = ~(return_mult_generic_AC_RND_CONV_false_4_op1_zero_sva_1 | return_mult_generic_AC_RND_CONV_false_3_op2_zero_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_3_r_nan_sva_1 = return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1
      | (operator_11_true_return_15_sva & (~ return_extract_17_m_zero_sva)) | (return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1
      & return_mult_generic_AC_RND_CONV_false_3_op2_zero_sva_1) | (return_mult_generic_AC_RND_CONV_false_4_op1_zero_sva_1
      & return_mult_generic_AC_RND_CONV_false_3_op2_inf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_3_lor_lpi_3_dfm_1 = return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1
      | return_mult_generic_AC_RND_CONV_false_3_op2_inf_sva_1 | return_mult_generic_AC_RND_CONV_false_3_exp_ovf_lor_lpi_3_dfm_2
      | return_mult_generic_AC_RND_CONV_false_3_r_nan_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_3_return_mult_generic_AC_RND_CONV_false_3_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_3_if_1_and_1_tmp_1 | (z_out_45[12]));
  assign return_mult_generic_AC_RND_CONV_false_3_and_2_nl = return_mult_generic_AC_RND_CONV_false_3_if_1_and_1_tmp_1
      & (~ (z_out_45[12]));
  assign return_mult_generic_AC_RND_CONV_false_3_res_bef_rnd_3_53_1_lpi_3_dfm_1 =
      MUX1HOT_v_53_3_2((return_mult_generic_AC_RND_CONV_false_3_p_sva_1[104:52]),
      (return_mult_generic_AC_RND_CONV_false_3_p_sva_1[103:51]), (z_out_35[53:1]),
      {return_mult_generic_AC_RND_CONV_false_3_return_mult_generic_AC_RND_CONV_false_3_nor_nl
      , return_mult_generic_AC_RND_CONV_false_3_and_2_nl , (z_out_45[12])});
  assign return_mult_generic_AC_RND_CONV_false_3_op2_inf_sva_1 = operator_11_true_return_15_sva
      & return_extract_17_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_3_op2_zero_sva_1 = return_extract_15_return_extract_15_nor_cse_sva
      & return_extract_17_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_3_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_3_if_acc_2_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva, z_out_45[12]);
  assign return_mult_generic_AC_RND_CONV_false_3_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_3_nl
      & (~ (return_mult_generic_AC_RND_CONV_false_3_p_sva_1[105]));
  assign return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      operator_33_true_15_acc_2, return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva);
  assign return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_5_if_acc_1_itm_12_1) | (return_mult_generic_AC_RND_CONV_false_5_p_sva_1[105]);
  assign return_mult_generic_AC_RND_CONV_false_5_if_if_not_nl = ~ (operator_6_false_45_acc_psp_sva_1[12]);
  assign return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      (operator_6_false_45_acc_psp_sva_1[11:0]), return_mult_generic_AC_RND_CONV_false_5_if_if_not_nl);
  assign return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1 = ({return_extract_41_return_extract_41_or_1_cse_sva
      , (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[51:0])}) * ({return_extract_51_return_extract_51_or_sva_1
      , return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1});
  assign nl_return_mult_generic_AC_RND_CONV_false_5_exp_acc_1_nl = conv_u2u_11_12({return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1
      , return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1}) + conv_u2u_1_12(~
      return_extract_41_return_extract_41_or_1_cse_sva) + 12'b000000000001;
  assign return_mult_generic_AC_RND_CONV_false_5_exp_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_5_exp_acc_1_nl[11:0];
  assign nl_return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp = conv_u2s_12_13(return_mult_generic_AC_RND_CONV_false_5_exp_acc_1_nl)
      + conv_s2s_11_13({1'b1 , (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[61:52])}) + conv_u2s_1_13(return_extract_51_return_extract_51_nor_tmp);
  assign return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp = nl_return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp[12:0];
  assign nl_operator_6_false_45_acc_psp_sva_1 = return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp
      + conv_s2s_7_13({1'b1 , (~ leading_sign_53_0_5_out_1)}) + 13'b0000000000001;
  assign operator_6_false_45_acc_psp_sva_1 = nl_operator_6_false_45_acc_psp_sva_1[12:0];
  assign return_mult_generic_AC_RND_CONV_false_5_if_nor_ovfl_sva_1 = ~((return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp[9:6]==4'b1111));
  assign return_mult_generic_AC_RND_CONV_false_5_e_incr_lpi_3_dfm_2 = ~((~(((return_mult_generic_AC_RND_CONV_false_5_p_sva_1[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((return_mult_generic_AC_RND_CONV_false_5_p_sva_1[51]) | return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_or_2))
      | (return_mult_generic_AC_RND_CONV_false_5_p_sva_1[105]))) | (return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp[12]));
  assign return_mult_generic_AC_RND_CONV_false_5_zero_m_return_mult_generic_AC_RND_CONV_false_5_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_5_r_zero_return_mult_generic_AC_RND_CONV_false_5_r_zero_nor_mdf_sva_1
      = ~(return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 | (return_extract_51_return_extract_51_nor_tmp
      & return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp));
  assign return_mult_generic_AC_RND_CONV_false_5_op2_inf_sva_1 = operator_11_true_51_operator_11_true_51_and_tmp
      & return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp;
  assign return_extract_51_return_extract_51_nor_tmp = ~((return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1);
  assign return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp = ~(return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_mux_1_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_5_if_acc_1_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva, return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp[12]);
  assign return_mult_generic_AC_RND_CONV_false_5_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_mux_1_nl
      & (~ (return_mult_generic_AC_RND_CONV_false_5_p_sva_1[105]));
  assign return_extract_51_return_extract_51_or_sva_1 = (return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_19_r_nan_or_1_nl = operator_11_true_return_15_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | (operator_11_true_return_13_sva
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva & return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign and_376_nl = (~((~((~ (stage_u_add_3_acc_itm_rsp_1[11])) & return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva)) & (~((return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[53])
      & return_add_generic_AC_RND_CONV_false_19_if_5_return_add_generic_AC_RND_CONV_false_19_if_5_and_tmp))
      & and_dcpl_314;
  assign return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_19_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_6_res_rounded_lpi_3_dfm_51_0_1[51]),
      and_376_nl);
  assign return_add_generic_AC_RND_CONV_false_19_if_7_return_add_generic_AC_RND_CONV_false_19_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_19_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_6_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_19_if_7_return_add_generic_AC_RND_CONV_false_19_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_19_mux_18_nl = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_and_9,
      (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_1[9:0]),
      return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_not_3_nl = ~ return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1;
  assign return_add_generic_AC_RND_CONV_false_19_e_r_qelse_return_add_generic_AC_RND_CONV_false_19_e_r_qelse_and_nl
      = MUX_v_10_2_2(10'b0000000000, return_add_generic_AC_RND_CONV_false_19_mux_18_nl,
      return_add_generic_AC_RND_CONV_false_6_e_r_qelse_not_3_nl);
  assign return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_19_e_r_qelse_return_add_generic_AC_RND_CONV_false_19_e_r_qelse_and_nl,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_19_exception_sva_1);
  assign return_add_generic_AC_RND_CONV_false_19_mux_19_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_and_11,
      return_add_generic_AC_RND_CONV_false_19_exp_plus_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[53]);
  assign or_241_nl = or_dcpl_212 | or_dcpl_183 | and_dcpl_129;
  assign return_add_generic_AC_RND_CONV_false_19_e_r_qelse_mux_2_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs, or_241_nl);
  assign return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_19_mux_19_nl
      & (~ return_add_generic_AC_RND_CONV_false_19_e_r_qelse_mux_2_nl)) | return_add_generic_AC_RND_CONV_false_19_exception_sva_1;
  assign operator_11_true_51_operator_11_true_51_and_tmp = (return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_19_if_5_return_add_generic_AC_RND_CONV_false_19_if_5_and_tmp
      = (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_19_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_19_if_5_or_nl = return_add_generic_AC_RND_CONV_false_19_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_19_if_5_return_add_generic_AC_RND_CONV_false_19_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_19_mux_16_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_19_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_19_if_5_or_nl, return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_19_exception_sva_1 = operator_11_true_return_13_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | operator_11_true_return_15_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_19_mux_16_nl;
  assign return_add_generic_AC_RND_CONV_false_19_exp_plus_1_0_lpi_3_dfm_1 = operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1
      | (~ return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva);
  assign return_add_generic_AC_RND_CONV_false_19_r_inf_lpi_3_dfm_2 = ((stage_u_add_3_acc_itm_rsp_1[11])
      | (~ return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva;
  assign return_mult_generic_AC_RND_CONV_false_5_shift_right_conc_3_5 = (~ (return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp[5]))
      | return_mult_generic_AC_RND_CONV_false_5_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_5_if_not_nl = ~ return_mult_generic_AC_RND_CONV_false_5_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_5_shift_right_conc_3_4_1 = ~(MUX_v_4_2_2(4'b0000,
      (return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp[4:1]), return_mult_generic_AC_RND_CONV_false_5_if_not_nl));
  assign return_mult_generic_AC_RND_CONV_false_5_shift_right_conc_3_0 = (~ (return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp[0]))
      | return_mult_generic_AC_RND_CONV_false_5_if_nor_ovfl_sva_1;
  assign drf_qr_lval_26_smx_lpi_3_dfm_mx0 = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1,
      BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0, and_dcpl_219);
  assign return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[0])
      & return_add_generic_AC_RND_CONV_false_11_mux_itm;
  assign return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1,
      and_dcpl_219);
  assign return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_51_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0,
      and_dcpl_219);
  assign return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2(reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_219);
  assign return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_219);
  assign return_add_generic_AC_RND_CONV_false_20_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[54]))) | (return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[53]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[52]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[51]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[50]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[49]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[48]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[47]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[46]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[45]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[44]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[43]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[42]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[41]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[40]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[39]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[38]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[37]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[36]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[35]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[34]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[33]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[32]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[31]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[30]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[29]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[28]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[27]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[26]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[25]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[24]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[23]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[22]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[21]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[20]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[19]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[18]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[17]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[16]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[15]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[14]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[13]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[12]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[11]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[10]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[9]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[8]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[7]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[6]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[5]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[4]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[3]))) | (return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_20_lshift_itm[2])));
  assign return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1 = (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm[0])
      & return_add_generic_AC_RND_CONV_false_21_unequal_tmp;
  assign return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(drf_qr_lval_14_smx_0_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1,
      and_dcpl_249);
  assign return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_51_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0,
      and_dcpl_249);
  assign return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_249);
  assign return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_249);
  assign nl_return_add_generic_AC_RND_CONV_false_21_ma1_lt_ma2_acc_1_nl = ({1'b1
      , return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm , return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm})
      + conv_u2u_52_53({(~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx1)
      , (~ return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1)}) + 53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_21_ma1_lt_ma2_acc_1_nl = nl_return_add_generic_AC_RND_CONV_false_21_ma1_lt_ma2_acc_1_nl[52:0];
  assign return_add_generic_AC_RND_CONV_false_21_ma1_lt_ma2_acc_1_itm_52 = readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_21_ma1_lt_ma2_acc_1_nl);
  assign return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_and_cse
      = return_add_generic_AC_RND_CONV_false_21_ma1_lt_ma2_acc_1_itm_52 & return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_21_op1_smaller_lor_lpi_3_dfm_2 = return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp[11]);
  assign return_add_generic_AC_RND_CONV_false_21_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_37[54]))) | (return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (z_out_37[53]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_37[52]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_37[51]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_37[50]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_37[49]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_37[48]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_37[47]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_37[46]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_37[45]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_37[44]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_37[43]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_37[42]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_37[41]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_37[40]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_37[39]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_37[38]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_37[37]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_37[36]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_37[35]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_37[34]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_37[33]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_37[32]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_37[31]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_37[30]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_37[29]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_37[28]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_37[27]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_37[26]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_37[25]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_37[24]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_37[23]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_37[22]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_37[21]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_37[20]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_37[19]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_37[18]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_37[17]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_37[16]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_37[15]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_37[14]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_37[13]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_37[12]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_37[11]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_37[10]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_37[9]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_37[8]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_37[7]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_37[6]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_37[5]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_37[4]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_37[3]))) | (return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_37[2])));
  assign return_add_generic_AC_RND_CONV_false_20_res_rounded_and_nl = (return_add_generic_AC_RND_CONV_false_20_res_rounded_asn_rndc_sva_1[3])
      & ((return_add_generic_AC_RND_CONV_false_20_res_rounded_asn_rndc_sva_1[0])
      | (return_add_generic_AC_RND_CONV_false_20_res_rounded_asn_rndc_sva_1[1]) |
      (return_add_generic_AC_RND_CONV_false_20_res_rounded_asn_rndc_sva_1[2]) | (return_add_generic_AC_RND_CONV_false_20_res_rounded_asn_rndc_sva_1[4]));
  assign nl_return_add_generic_AC_RND_CONV_false_20_res_rounded_acc_tmp = conv_u2u_53_54(return_add_generic_AC_RND_CONV_false_20_res_rounded_asn_rndc_sva_1[56:4])
      + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_20_res_rounded_and_nl);
  assign return_add_generic_AC_RND_CONV_false_20_res_rounded_acc_tmp = nl_return_add_generic_AC_RND_CONV_false_20_res_rounded_acc_tmp[53:0];
  assign return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 = operator_11_true_return_13_sva
      & (~ return_extract_17_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1 = operator_11_true_return_13_sva
      & return_extract_17_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_20_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_12_mux_itm);
  assign and_378_nl = or_dcpl_625 & (~(return_add_generic_AC_RND_CONV_false_20_if_5_return_add_generic_AC_RND_CONV_false_20_if_5_and_1_tmp
      & (return_add_generic_AC_RND_CONV_false_20_res_rounded_acc_tmp[53]))) & and_dcpl_316;
  assign return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_20_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_20_res_rounded_lpi_3_dfm_51_0_1[51]),
      and_378_nl);
  assign return_add_generic_AC_RND_CONV_false_20_not_3_nl = ~ (return_add_generic_AC_RND_CONV_false_20_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_20_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_20_res_rounded_acc_tmp[51:0]), return_add_generic_AC_RND_CONV_false_20_not_3_nl);
  assign nl_operator_33_true_43_acc_nl = conv_s2s_11_12({operator_6_false_49_acc_psp_sva_11_9
      , (operator_6_false_49_acc_psp_sva_8_0[8:1])}) + 12'b000000000001;
  assign operator_33_true_43_acc_nl = nl_operator_33_true_43_acc_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_21_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      operator_33_true_43_acc_nl, return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_21_res_rounded_and_cse = (z_out_39[3])
      & ((z_out_39[0]) | (z_out_39[1]) | (z_out_39[2]) | (z_out_39[4]));
  assign nl_return_add_generic_AC_RND_CONV_false_21_res_rounded_acc_tmp = conv_u2u_53_54(z_out_39[56:4])
      + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_21_res_rounded_and_cse);
  assign return_add_generic_AC_RND_CONV_false_21_res_rounded_acc_tmp = nl_return_add_generic_AC_RND_CONV_false_21_res_rounded_acc_tmp[53:0];
  assign return_add_generic_AC_RND_CONV_false_21_not_3_nl = ~ (return_add_generic_AC_RND_CONV_false_21_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_21_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_21_res_rounded_acc_tmp[51:0]), return_add_generic_AC_RND_CONV_false_21_not_3_nl);
  assign return_add_generic_AC_RND_CONV_false_21_op1_nan_sva_1 = operator_11_true_return_17_sva
      & (~ return_extract_1_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_21_op1_inf_sva_1 = operator_11_true_return_17_sva
      & return_extract_1_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_20_e_r_qelse_not_2_nl = ~ return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs_mx0w0;
  assign return_add_generic_AC_RND_CONV_false_20_e_r_qelse_return_add_generic_AC_RND_CONV_false_20_e_r_qelse_and_nl
      = MUX_v_10_2_2(10'b0000000000, z_out_44, return_add_generic_AC_RND_CONV_false_20_e_r_qelse_not_2_nl);
  assign return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_20_e_r_qelse_return_add_generic_AC_RND_CONV_false_20_e_r_qelse_and_nl,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_20_exception_sva_1);
  assign return_add_generic_AC_RND_CONV_false_20_mux_21_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_and_11,
      return_add_generic_AC_RND_CONV_false_7_exp_plus_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_20_res_rounded_acc_tmp[53]);
  assign or_245_nl = or_dcpl_193 | and_dcpl_131 | operator_11_true_return_13_sva;
  assign return_add_generic_AC_RND_CONV_false_20_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs, or_245_nl);
  assign return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_20_mux_21_nl
      & (~ return_add_generic_AC_RND_CONV_false_20_e_r_qelse_mux_1_nl)) | return_add_generic_AC_RND_CONV_false_20_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_20_if_7_return_add_generic_AC_RND_CONV_false_20_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_20_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_20_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_20_if_7_return_add_generic_AC_RND_CONV_false_20_if_7_nor_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0w0 = ({1'b1
      , return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1})
      + conv_u2s_11_12(~ (stage_PE_1_x_re_d_sva[62:52])) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0w0 = nl_return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0w0[11:0];
  assign nl_return_add_generic_AC_RND_CONV_false_22_e_dif1_acc_1_tmp = ({1'b1 , (stage_PE_1_x_re_d_sva[62:52])})
      + conv_u2s_11_12({(~ return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1)
      , (~ return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1)}) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_22_e_dif1_acc_1_tmp = nl_return_add_generic_AC_RND_CONV_false_22_e_dif1_acc_1_tmp[11:0];
  assign return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(return_add_generic_AC_RND_CONV_false_22_e_dif1_acc_1_tmp,
      return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0w0, return_add_generic_AC_RND_CONV_false_22_e_dif1_acc_1_tmp[11]);
  assign return_extract_57_return_extract_57_or_2_nl = (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_extract_57_return_extract_57_or_2_nl,
      return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1[50]), return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0 = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1[50:1]),
      (return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1[49:0]), return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1[0])
      & (~ return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0,
      and_dcpl_241);
  assign return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_51_lpi_3_dfm_mx0 =
      MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0[50]), return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0,
      and_dcpl_241);
  assign return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0[49:0]),
      return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_241);
  assign return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1,
      and_dcpl_241);
  assign return_add_generic_AC_RND_CONV_false_22_e1_eq_e2_equal_tmp = (stage_PE_1_x_re_d_sva[62:52])
      == ({return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1});
  assign return_add_generic_AC_RND_CONV_false_22_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_40[54]))) | (return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (z_out_40[53]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_40[52]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_40[51]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_40[50]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_40[49]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_40[48]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_40[47]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_40[46]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_40[45]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_40[44]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_40[43]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_40[42]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_40[41]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_40[40]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_40[39]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_40[38]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_40[37]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_40[36]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_40[35]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_40[34]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_40[33]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_40[32]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_40[31]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_40[30]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_40[29]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_40[28]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_40[27]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_40[26]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_40[25]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_40[24]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_40[23]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_40[22]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_40[21]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_40[20]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_40[19]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_40[18]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_40[17]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_40[16]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_40[15]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_40[14]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_40[13]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_40[12]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_40[11]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_40[10]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_40[9]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_40[8]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_40[7]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_40[6]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_40[5]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_40[4]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_40[3]))) | (return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_40[2])));
  assign nl_return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0w0 = ({1'b1
      , return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_mx1w0 , return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1})
      + conv_u2s_11_12(~ (stage_PE_1_x_im_d_sva[62:52])) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0w0 = nl_return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0w0[11:0];
  assign nl_return_add_generic_AC_RND_CONV_false_23_e_dif1_acc_1_tmp = ({1'b1 , (stage_PE_1_x_im_d_sva[62:52])})
      + conv_u2s_11_12({(~ return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_mx1w0)
      , (~ return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1)}) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_23_e_dif1_acc_1_tmp = nl_return_add_generic_AC_RND_CONV_false_23_e_dif1_acc_1_tmp[11:0];
  assign return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(return_add_generic_AC_RND_CONV_false_23_e_dif1_acc_1_tmp,
      return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0w0, return_add_generic_AC_RND_CONV_false_23_e_dif1_acc_1_tmp[11]);
  assign return_extract_59_return_extract_59_or_2_nl = (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_mx1w0!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_extract_59_return_extract_59_or_2_nl,
      return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm_mx2, return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm_mx2,
      (return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_mx0w6[50]), return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0 = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_mx0w6[50:1]),
      (return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_mx0w6[49:0]), return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_mx0w6[0])
      & (~ return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0, and_dcpl_196);
  assign return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_51_lpi_3_dfm_mx0 =
      MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[50]),
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0, and_dcpl_196);
  assign return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[49:0]),
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_196);
  assign return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1,
      and_dcpl_196);
  assign return_add_generic_AC_RND_CONV_false_23_e1_eq_e2_equal_tmp = (stage_PE_1_x_im_d_sva[62:52])
      == ({return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_mx1w0 ,
      return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1});
  assign return_add_generic_AC_RND_CONV_false_23_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[54]))) | (return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[53]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[52]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[51]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[50]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[49]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[48]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[47]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[46]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[45]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[44]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[43]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[42]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[41]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[40]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[39]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[38]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[37]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[36]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[35]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[34]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[33]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[32]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[31]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[30]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[29]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[28]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[27]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[26]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[25]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[24]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[23]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[22]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[21]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[20]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[19]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[18]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[17]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[16]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[15]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[14]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[13]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[12]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[11]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[10]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[9]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[8]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[7]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[6]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[5]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[4]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[3]))) | (return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (return_add_generic_AC_RND_CONV_false_23_lshift_itm[2])));
  assign return_add_generic_AC_RND_CONV_false_24_e_dif_qr_lpi_3_dfm_mx0_10_0 = MUX_v_11_2_2((return_add_generic_AC_RND_CONV_false_22_e_dif1_acc_1_tmp[10:0]),
      (return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0w0[10:0]), return_add_generic_AC_RND_CONV_false_22_e_dif1_acc_1_tmp[11]);
  assign return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0,
      and_dcpl_228);
  assign return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_51_lpi_3_dfm_mx0 =
      MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0[50]), return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0,
      and_dcpl_228);
  assign return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0[49:0]),
      return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_228);
  assign return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1,
      and_dcpl_228);
  assign return_add_generic_AC_RND_CONV_false_24_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_38[54]))) | (return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (z_out_38[53]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_38[52]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_38[51]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_38[50]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_38[49]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_38[48]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_38[47]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_38[46]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_38[45]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_38[44]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_38[43]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_38[42]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_38[41]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_38[40]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_38[39]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_38[38]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_38[37]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_38[36]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_38[35]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_38[34]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_38[33]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_38[32]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_38[31]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_38[30]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_38[29]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_38[28]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_38[27]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_38[26]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_38[25]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_38[24]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_38[23]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_38[22]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_38[21]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_38[20]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_38[19]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_38[18]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_38[17]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_38[16]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_38[15]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_38[14]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_38[13]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_38[12]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_38[11]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_38[10]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_38[9]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_38[8]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_38[7]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_38[6]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_38[5]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_38[4]))) | ((return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_38[3]))) | (return_add_generic_AC_RND_CONV_false_24_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_38[2])));
  assign return_add_generic_AC_RND_CONV_false_25_e_dif_qr_lpi_3_dfm_mx0_10_0 = MUX_v_11_2_2((return_add_generic_AC_RND_CONV_false_23_e_dif1_acc_1_tmp[10:0]),
      (return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0w0[10:0]), return_add_generic_AC_RND_CONV_false_23_e_dif1_acc_1_tmp[11]);
  assign return_add_generic_AC_RND_CONV_false_25_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_42[54]))) | (return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (z_out_42[53]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_42[52]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_42[51]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_42[50]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_42[49]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_42[48]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_42[47]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_42[46]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_42[45]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_42[44]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_42[43]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_42[42]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_42[41]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_42[40]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_42[39]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_42[38]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_42[37]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_42[36]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_42[35]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_42[34]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_42[33]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_42[32]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_42[31]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_42[30]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_42[29]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_42[28]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_42[27]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_42[26]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_42[25]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_42[24]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_42[23]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_42[22]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_42[21]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_42[20]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_42[19]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_42[18]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_42[17]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_42[16]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_42[15]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_42[14]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_42[13]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_42[12]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_42[11]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_42[10]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_42[9]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_42[8]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_42[7]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_42[6]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_42[5]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_42[4]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_42[3]))) | (return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_42[2])));
  assign return_add_generic_AC_RND_CONV_false_25_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_25_e_dif_qr_lpi_3_dfm_mx0_10_0[10:6]!=5'b00000)
      | ((return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0w0[11]) &
      (return_add_generic_AC_RND_CONV_false_23_e_dif1_acc_1_tmp[11]));
  assign return_add_generic_AC_RND_CONV_false_25_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_25_e_dif_qr_lpi_3_dfm_mx0_10_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_25_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_24_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_24_e_dif_qr_lpi_3_dfm_mx0_10_0[10:6]!=5'b00000)
      | ((return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0w0[11]) &
      (return_add_generic_AC_RND_CONV_false_22_e_dif1_acc_1_tmp[11]));
  assign return_add_generic_AC_RND_CONV_false_24_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_24_e_dif_qr_lpi_3_dfm_mx0_10_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_24_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_23_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_23_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_23_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp
      = ~((return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_mx1w0!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_22_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_22_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_22_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp
      = ~((return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_21_if_5_return_add_generic_AC_RND_CONV_false_21_if_5_and_tmp
      = (return_add_generic_AC_RND_CONV_false_21_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_21_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_21_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_21_if_5_or_nl = return_add_generic_AC_RND_CONV_false_8_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_21_if_5_return_add_generic_AC_RND_CONV_false_21_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_21_mux_14_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_21_if_5_or_nl, return_add_generic_AC_RND_CONV_false_21_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_21_exception_sva_1 = return_add_generic_AC_RND_CONV_false_21_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_21_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_21_mux_14_nl;
  assign return_add_generic_AC_RND_CONV_false_21_exp_plus_1_0_lpi_3_dfm_1 = (operator_6_false_49_acc_psp_sva_8_0[0])
      | (~ return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_21_mux_8_itm_3_0 = MUX_v_4_2_2((reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[3:0]),
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2, return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_20_mux_18_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_7_if_5_or_cse, return_add_generic_AC_RND_CONV_false_20_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_20_exception_sva_1 = return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_20_mux_18_nl;
  assign return_add_generic_AC_RND_CONV_false_22_op1_nan_sva_1 = operator_11_true_return_24_sva
      & (~ return_extract_12_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_22_op1_inf_sva_1 = operator_11_true_return_24_sva
      & return_extract_12_m_zero_sva;
  assign nl_operator_33_true_46_acc_tmp = conv_s2s_7_13({operator_6_false_6_operator_6_false_6_conc_2_6_1
      , (~ (leading_sign_57_0_1_0_15_out_3[0]))}) + conv_u2s_11_13({reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0
      , reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1 , drf_qr_lval_14_smx_0_lpi_3_dfm});
  assign operator_33_true_46_acc_tmp = nl_operator_33_true_46_acc_tmp[12:0];
  assign nl_return_add_generic_AC_RND_CONV_false_23_acc_2_nl =  -(operator_33_true_46_acc_tmp[11:0]);
  assign return_add_generic_AC_RND_CONV_false_23_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_23_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_23_acc_2_nl);
  assign nl_operator_33_true_47_acc_nl = conv_s2s_11_12(z_out_13[11:1]) + 12'b000000000001;
  assign operator_33_true_47_acc_nl = nl_operator_33_true_47_acc_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_23_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      operator_33_true_47_acc_nl, return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_23_res_rounded_and_nl = (z_out_41[3])
      & ((z_out_41[0]) | (z_out_41[1]) | (z_out_41[2]) | (z_out_41[4]));
  assign nl_return_add_generic_AC_RND_CONV_false_23_res_rounded_acc_tmp = conv_u2u_53_54(z_out_41[56:4])
      + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_23_res_rounded_and_nl);
  assign return_add_generic_AC_RND_CONV_false_23_res_rounded_acc_tmp = nl_return_add_generic_AC_RND_CONV_false_23_res_rounded_acc_tmp[53:0];
  assign return_add_generic_AC_RND_CONV_false_23_op1_nan_sva_1 = operator_11_true_return_26_sva
      & (~ return_extract_15_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_23_op1_inf_sva_1 = operator_11_true_return_26_sva
      & return_extract_15_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_23_not_3_nl = ~ (return_add_generic_AC_RND_CONV_false_23_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_23_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_23_res_rounded_acc_tmp[51:0]), return_add_generic_AC_RND_CONV_false_23_not_3_nl);
  assign nl_operator_6_false_54_acc_nl = ({1'b1 , (~ (leading_sign_57_0_1_0_24_out_3[5:1]))})
      + 6'b000001;
  assign operator_6_false_54_acc_nl = nl_operator_6_false_54_acc_nl[5:0];
  assign nl_operator_33_true_48_acc_tmp = conv_s2s_7_13({operator_6_false_54_acc_nl
      , (~ (leading_sign_57_0_1_0_24_out_3[0]))}) + conv_u2s_11_13({return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_itm
      , BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm});
  assign operator_33_true_48_acc_tmp = nl_operator_33_true_48_acc_tmp[12:0];
  assign nl_return_add_generic_AC_RND_CONV_false_24_acc_2_nl =  -(operator_33_true_48_acc_tmp[11:0]);
  assign return_add_generic_AC_RND_CONV_false_24_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_24_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_24_acc_2_nl);
  assign nl_operator_33_true_49_acc_nl = conv_s2s_11_12(operator_6_false_55_acc_psp_sva_1[11:1])
      + 12'b000000000001;
  assign operator_33_true_49_acc_nl = nl_operator_33_true_49_acc_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_24_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      operator_33_true_49_acc_nl, return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11);
  assign nl_return_add_generic_AC_RND_CONV_false_24_res_rounded_acc_tmp = conv_u2u_53_54(z_out_38[56:4])
      + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_18_res_rounded_and_cse);
  assign return_add_generic_AC_RND_CONV_false_24_res_rounded_acc_tmp = nl_return_add_generic_AC_RND_CONV_false_24_res_rounded_acc_tmp[53:0];
  assign return_add_generic_AC_RND_CONV_false_24_not_3_nl = ~ (return_add_generic_AC_RND_CONV_false_24_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_24_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_24_res_rounded_acc_tmp[51:0]), return_add_generic_AC_RND_CONV_false_24_not_3_nl);
  assign nl_operator_6_false_56_acc_nl = ({1'b1 , (~ (leading_sign_57_0_1_0_25_out_3[5:1]))})
      + 6'b000001;
  assign operator_6_false_56_acc_nl = nl_operator_6_false_56_acc_nl[5:0];
  assign nl_operator_33_true_50_acc_tmp = conv_s2s_7_13({operator_6_false_56_acc_nl
      , (~ (leading_sign_57_0_1_0_25_out_3[0]))}) + conv_u2s_11_13({in_u_rsc_merge_sva_rsp_1_rsp_0
      , in_u_rsc_merge_sva_rsp_1_rsp_1 , return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm});
  assign operator_33_true_50_acc_tmp = nl_operator_33_true_50_acc_tmp[12:0];
  assign nl_return_add_generic_AC_RND_CONV_false_25_acc_2_nl =  -(operator_33_true_50_acc_tmp[11:0]);
  assign return_add_generic_AC_RND_CONV_false_25_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_25_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_25_acc_2_nl);
  assign nl_operator_33_true_51_acc_nl = conv_s2s_11_12(z_out_52[11:1]) + 12'b000000000001;
  assign operator_33_true_51_acc_nl = nl_operator_33_true_51_acc_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_25_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      operator_33_true_51_acc_nl, return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11);
  assign return_add_generic_AC_RND_CONV_false_25_res_rounded_and_nl = (z_out_40[3])
      & ((z_out_40[0]) | (z_out_40[1]) | (z_out_40[2]) | (z_out_40[4]));
  assign nl_return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp = conv_u2u_53_54(z_out_40[56:4])
      + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_25_res_rounded_and_nl);
  assign return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp = nl_return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp[53:0];
  assign return_add_generic_AC_RND_CONV_false_25_not_3_nl = ~ (return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_25_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp[51:0]), return_add_generic_AC_RND_CONV_false_25_not_3_nl);
  assign return_add_generic_AC_RND_CONV_false_25_exp_plus_1_0_lpi_3_dfm_1 = (z_out_52[0])
      | (~ return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11);
  assign return_add_generic_AC_RND_CONV_false_25_r_inf_lpi_3_dfm_2 = ((operator_33_true_50_acc_tmp[11])
      | (~ return_add_generic_AC_RND_CONV_false_25_else_4_return_add_generic_AC_RND_CONV_false_25_else_4_nand_tmp))
      & return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11;
  assign return_add_generic_AC_RND_CONV_false_24_exp_plus_1_0_lpi_3_dfm_1 = (operator_6_false_55_acc_psp_sva_1[0])
      | (~ return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11);
  assign return_add_generic_AC_RND_CONV_false_24_r_inf_lpi_3_dfm_2 = ((operator_33_true_48_acc_tmp[11])
      | (~ return_add_generic_AC_RND_CONV_false_24_else_4_return_add_generic_AC_RND_CONV_false_24_else_4_nand_tmp))
      & return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11;
  assign nl_operator_6_false_55_acc_psp_sva_1 = conv_u2s_11_12({return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_itm
      , BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm}) + conv_s2s_7_12({1'b1
      , (~ leading_sign_57_0_1_0_24_out_3)}) + 12'b000000000001;
  assign operator_6_false_55_acc_psp_sva_1 = nl_operator_6_false_55_acc_psp_sva_1[11:0];
  assign return_add_generic_AC_RND_CONV_false_23_exp_plus_1_0_lpi_3_dfm_1 = (z_out_13[0])
      | (~ return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_23_if_5_return_add_generic_AC_RND_CONV_false_23_if_5_and_tmp
      = (return_add_generic_AC_RND_CONV_false_23_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_23_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_23_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_23_if_5_or_nl = return_add_generic_AC_RND_CONV_false_23_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_23_if_5_return_add_generic_AC_RND_CONV_false_23_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_23_mux_17_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_23_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_23_if_5_or_nl, return_add_generic_AC_RND_CONV_false_23_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_23_exception_sva_1 = return_add_generic_AC_RND_CONV_false_23_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_23_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_23_mux_17_nl;
  assign return_add_generic_AC_RND_CONV_false_23_r_inf_lpi_3_dfm_2 = ((operator_33_true_46_acc_tmp[11])
      | (~ return_add_generic_AC_RND_CONV_false_23_else_4_return_add_generic_AC_RND_CONV_false_23_else_4_nand_tmp))
      & return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_22_exception_sva_1 = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1 | return_add_generic_AC_RND_CONV_false_22_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_9_mux_17_cse;
  assign return_add_generic_AC_RND_CONV_false_22_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_22_exception_sva_1
      | leading_sign_57_0_1_0_2_out_2;
  assign return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1) | (z_out_54[105]);
  assign return_mult_generic_AC_RND_CONV_false_6_if_if_not_nl = ~ (operator_6_false_58_acc_psp_sva_1[11]);
  assign return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3 = MUX_v_11_2_2(11'b00000000000,
      (operator_6_false_58_acc_psp_sva_1[10:0]), return_mult_generic_AC_RND_CONV_false_6_if_if_not_nl);
  assign nl_operator_6_false_58_acc_psp_sva_1 = z_out_51 + conv_s2s_7_12({1'b1 ,
      (~ leading_sign_53_0_6_out_1)}) + 12'b000000000001;
  assign operator_6_false_58_acc_psp_sva_1 = nl_operator_6_false_58_acc_psp_sva_1[11:0];
  assign return_mult_generic_AC_RND_CONV_false_6_e_incr_lpi_2_dfm_2 = ~((~(((z_out_54[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((z_out_54[51]) | return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_or_2))
      | (z_out_54[105]))) | (z_out_51[11]));
  assign return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1
      = ~((out_f_d_rsci_q_d[62:52]==11'b00000000000) & return_extract_3_m_zero_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_6_lor_lpi_2_dfm_1 = (operator_11_true_return_3_sva_mx1w0
      & return_extract_3_m_zero_sva_1) | ((return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3==11'b11111111110)
      & return_mult_generic_AC_RND_CONV_false_6_e_incr_lpi_2_dfm_2) | return_mult_generic_AC_RND_CONV_false_6_op1_nan_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_6_op1_nan_sva_1 = operator_11_true_return_3_sva_mx1w0
      & (~ return_extract_3_m_zero_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1 = (~ return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_6_lor_lpi_2_dfm_1;
  assign return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_6_if_1_and_1_tmp_1 | (z_out_51[11]));
  assign return_mult_generic_AC_RND_CONV_false_6_and_2_nl = return_mult_generic_AC_RND_CONV_false_6_if_1_and_1_tmp_1
      & (~ (z_out_51[11]));
  assign return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1 =
      MUX1HOT_v_53_3_2((z_out_54[104:52]), (z_out_54[103:51]), (z_out_35[53:1]),
      {return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_nor_nl
      , return_mult_generic_AC_RND_CONV_false_6_and_2_nl , (z_out_51[11])});
  assign return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_mux_1_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1,
      return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva, z_out_51[11]);
  assign return_mult_generic_AC_RND_CONV_false_6_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_mux_1_nl
      & (~ (z_out_54[105]));
  assign nl_stage_monty_mul_acc_2_psp_sva_1 = z_out_48 + conv_u2s_14_15(signext_14_13({(z_out_48[14])
      , 11'b00000000000 , (z_out_48[14])}));
  assign stage_monty_mul_acc_2_psp_sva_1 = nl_stage_monty_mul_acc_2_psp_sva_1[14:0];
  assign nl_operator_32_false_2_mul_atp_sva_1 = (~ (in_u_rsci_q_d[9:0])) + 10'b0000000001;
  assign operator_32_false_2_mul_atp_sva_1 = nl_operator_32_false_2_mul_atp_sva_1[9:0];
  assign nl_operator_6_false_6_operator_6_false_6_conc_2_6_1 = ({1'b1 , (~ (leading_sign_57_0_1_0_15_out_3[5:1]))})
      + 6'b000001;
  assign operator_6_false_6_operator_6_false_6_conc_2_6_1 = nl_operator_6_false_6_operator_6_false_6_conc_2_6_1[5:0];
  assign nl_return_add_generic_AC_RND_CONV_false_15_acc_3_nl =  -(z_out_13[11:0]);
  assign return_add_generic_AC_RND_CONV_false_15_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_15_acc_3_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_15_acc_3_nl);
  assign return_add_generic_AC_RND_CONV_false_15_if_5_return_add_generic_AC_RND_CONV_false_15_if_5_and_1_tmp
      = (return_add_generic_AC_RND_CONV_false_3_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_3_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_3_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign nl_operator_6_false_2_operator_6_false_2_conc_2_6_1 = ({1'b1 , (~ (leading_sign_57_0_1_0_2_out_3[5:1]))})
      + 6'b000001;
  assign operator_6_false_2_operator_6_false_2_conc_2_6_1 = nl_operator_6_false_2_operator_6_false_2_conc_2_6_1[5:0];
  assign nl_return_add_generic_AC_RND_CONV_false_2_acc_3_nl =  -(operator_33_true_4_acc_tmp[11:0]);
  assign return_add_generic_AC_RND_CONV_false_2_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_2_acc_3_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_2_acc_3_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_2_acc_3_nl);
  assign return_add_generic_AC_RND_CONV_false_2_if_5_return_add_generic_AC_RND_CONV_false_2_if_5_and_1_tmp
      = (return_add_generic_AC_RND_CONV_false_1_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_1_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_1_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign nl_return_add_generic_AC_RND_CONV_false_22_acc_3_nl =  -(operator_33_true_44_acc_tmp[11:0]);
  assign return_add_generic_AC_RND_CONV_false_22_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_22_acc_3_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_22_acc_3_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_22_acc_3_nl);
  assign return_add_generic_AC_RND_CONV_false_22_if_5_return_add_generic_AC_RND_CONV_false_22_if_5_and_1_tmp
      = (return_add_generic_AC_RND_CONV_false_9_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_9_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_9_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign nl_operator_6_false_10_operator_6_false_10_conc_2_6_1 = ({1'b1 , (~ (return_add_generic_AC_RND_CONV_false_20_ls_sva[5:1]))})
      + 6'b000001;
  assign operator_6_false_10_operator_6_false_10_conc_2_6_1 = nl_operator_6_false_10_operator_6_false_10_conc_2_6_1[5:0];
  assign nl_operator_33_true_15_acc_2 = conv_s2s_11_12({operator_6_false_18_acc_psp_sva_11
      , operator_6_false_18_acc_psp_sva_10_0_rsp_0 , operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0})
      + 12'b000000000001;
  assign operator_33_true_15_acc_2 = nl_operator_33_true_15_acc_2[11:0];
  assign return_add_generic_AC_RND_CONV_false_6_r_sign_mux_2 = MUX_s_1_2_2(stage_PE_1_tmp_re_d_1_lpi_3_dfm_63,
      (~ stage_PE_1_tmp_im_d_1_lpi_3_dfm_63), return_add_generic_AC_RND_CONV_false_19_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_nor_2
      = ~(stage_PE_1_tmp_im_d_1_lpi_3_dfm_63 | (~ stage_PE_1_tmp_re_d_1_lpi_3_dfm_63));
  assign return_add_generic_AC_RND_CONV_false_3_return_add_generic_AC_RND_CONV_false_3_and_8_nl
      = (z_out_13[0]) & return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_3_mux_26 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_3_return_add_generic_AC_RND_CONV_false_3_and_8_nl,
      return_add_generic_AC_RND_CONV_false_3_exp_plus_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_10_nl
      = (operator_33_true_4_acc_tmp[0]) & return_add_generic_AC_RND_CONV_false_2_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_1_mux_32 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_10_nl,
      return_add_generic_AC_RND_CONV_false_1_exp_plus_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_2_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_and_10_nl
      = (operator_33_true_44_acc_tmp[0]) & return_add_generic_AC_RND_CONV_false_22_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_9_mux_35 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_and_10_nl,
      return_add_generic_AC_RND_CONV_false_9_exp_plus_1_0_lpi_3_dfm_1, z_out_47[53]);
  assign return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_and_9
      = MUX_v_10_2_2(10'b0000000000, (stage_u_add_3_acc_itm_rsp_1[10:1]), return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva);
  assign nl_return_add_generic_AC_RND_CONV_false_10_acc_3_nl =  -(stage_u_add_3_acc_itm_rsp_1[11:0]);
  assign return_add_generic_AC_RND_CONV_false_10_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_10_acc_3_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_10_acc_3_nl);
  assign return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_and_9
      = MUX_v_10_2_2(10'b0000000000, (stage_u_add_3_acc_itm_rsp_1[10:1]), return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_20_if_5_return_add_generic_AC_RND_CONV_false_20_if_5_and_1_tmp
      = (return_add_generic_AC_RND_CONV_false_7_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_7_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_7_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_7_if_5_return_add_generic_AC_RND_CONV_false_7_if_5_nor_2
      = ~((stage_u_add_3_acc_itm_rsp_1!=13'b0000000000000));
  assign return_add_generic_AC_RND_CONV_false_7_if_5_or_3 = return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1
      | return_add_generic_AC_RND_CONV_false_7_if_5_return_add_generic_AC_RND_CONV_false_7_if_5_nor_2;
  assign return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_and_11
      = (stage_u_add_3_acc_itm_rsp_1[0]) & return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_6_if_5_or_3 = return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva
      | return_add_generic_AC_RND_CONV_false_7_if_5_return_add_generic_AC_RND_CONV_false_7_if_5_nor_2;
  assign return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_and_11
      = (stage_u_add_3_acc_itm_rsp_1[0]) & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva;
  assign nl_return_mult_generic_AC_RND_CONV_false_3_if_acc_2_nl =  -z_out_63;
  assign return_mult_generic_AC_RND_CONV_false_3_if_acc_2_nl = nl_return_mult_generic_AC_RND_CONV_false_3_if_acc_2_nl[12:0];
  assign return_mult_generic_AC_RND_CONV_false_3_if_acc_2_itm_12_1 = readslicef_13_1_12(return_mult_generic_AC_RND_CONV_false_3_if_acc_2_nl);
  assign return_mult_generic_AC_RND_CONV_false_if_1_or_1_nl = (return_mult_generic_AC_RND_CONV_false_3_p_sva_1[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_if_1_aelse_return_mult_generic_AC_RND_CONV_false_if_1_aelse_or_2
      & (return_mult_generic_AC_RND_CONV_false_3_p_sva_1[51]));
  assign return_mult_generic_AC_RND_CONV_false_mux_15 = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_if_1_or_1_nl,
      return_mult_generic_AC_RND_CONV_false_4_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_4_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_4_else_1_sticky_bit_or_cse,
      z_out_45[12]);
  assign return_mult_generic_AC_RND_CONV_false_3_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_3_exp_ovf_oif_aelse_and_1_tmp
      = (return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_1_cse[10:1]==10'b1111111111)
      & return_mult_generic_AC_RND_CONV_false_4_exp_ovf_oif_aelse_nor_cse & return_mult_generic_AC_RND_CONV_false_3_e_incr_lpi_3_dfm_2;
  assign return_mult_generic_AC_RND_CONV_false_else_2_else_else_mux_2 = MUX_v_11_2_2((return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_1_cse[10:0]),
      (z_out_55[10:0]), return_mult_generic_AC_RND_CONV_false_3_e_incr_lpi_3_dfm_2);
  assign nl_return_add_generic_AC_RND_CONV_false_21_acc_3_nl = ({(~ (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_2_1[0]))
      , (~ reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0) , (~ reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0)
      , (~ reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1)}) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_21_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_21_acc_3_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_21_acc_3_nl);
  assign return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_and_8
      = reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1 & return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_8_if_5_or_3 = return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1
      | (~((reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_2_1!=2'b00) | reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0
      | (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0!=9'b000000000)
      | reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1));
  assign return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_and_10_9
      = reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0 & return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_and_10_8_0
      = MUX_v_9_2_2(9'b000000000, reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0,
      return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1);
  assign or_dcpl_3 = ~(mode_lpi_1_dfm & BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm);
  assign nor_tmp = BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm & mode_lpi_1_dfm;
  assign and_dcpl_1 = mode_lpi_1_dfm & (~ inverse_lpi_1_dfm_1);
  assign or_dcpl_25 = return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva;
  assign or_dcpl_35 = (fsm_output[7:6]!=2'b00);
  assign and_dcpl_35 = ~(mode_lpi_1_dfm | inverse_lpi_1_dfm_1);
  assign and_dcpl_42 = or_dcpl_3 & (~ (z_out_49[9]));
  assign and_dcpl_44 = or_dcpl_3 & (~ (BUTTERFLY_mux_5_itm_9_0[9]));
  assign nor_8_cse = ~((fsm_output[36:35]!=2'b00));
  assign nl_for_acc_nl = conv_u2s_3_4(z_out_13[3:1]) + 4'b1011;
  assign for_acc_nl = nl_for_acc_nl[3:0];
  assign or_dcpl_60 = ~((~(t_in_10_0_lpi_1_dfm_1_1 & (~(t_in_10_0_lpi_1_dfm_1_10
      | t_in_10_0_lpi_1_dfm_1_9 | t_in_10_0_lpi_1_dfm_1_8 | t_in_10_0_lpi_1_dfm_1_7
      | t_in_10_0_lpi_1_dfm_1_6 | t_in_10_0_lpi_1_dfm_1_5 | t_in_10_0_lpi_1_dfm_1_4
      | t_in_10_0_lpi_1_dfm_1_3 | t_in_10_0_lpi_1_dfm_1_2)))) & (readslicef_4_1_3(for_acc_nl)));
  assign and_dcpl_74 = (operator_16_false_io_read_mode1_rsc_cse_sva[6:3]==4'b0000);
  assign and_dcpl_80 = ~((operator_16_false_io_read_mode1_rsc_cse_sva[15:14]!=2'b00));
  assign and_dcpl_83 = and_dcpl_80 & (operator_16_false_io_read_mode1_rsc_cse_sva[13:7]==7'b0000000);
  assign or_dcpl_64 = (operator_16_false_io_read_mode1_rsc_cse_sva[1:0]!=2'b01);
  assign or_dcpl_65 = (operator_16_false_io_read_mode1_rsc_cse_sva[3:2]!=2'b00);
  assign or_dcpl_69 = (operator_16_false_io_read_mode1_rsc_cse_sva[7:4]!=4'b0000);
  assign or_dcpl_75 = (operator_16_false_io_read_mode1_rsc_cse_sva[15:14]!=2'b00);
  assign or_dcpl_77 = or_dcpl_75 | (operator_16_false_io_read_mode1_rsc_cse_sva[13:8]!=6'b000000);
  assign and_dcpl_85 = ~((~(or_dcpl_77 | or_dcpl_69 | or_dcpl_65 | or_dcpl_64)) |
      operator_16_false_operator_16_false_nor_cse_sva);
  assign and_dcpl_91 = ~((~(or_dcpl_77 | or_dcpl_69 | or_dcpl_65 | (~((operator_16_false_io_read_mode1_rsc_cse_sva[1])
      ^ (operator_16_false_io_read_mode1_rsc_cse_sva[0]))))) | operator_16_false_operator_16_false_nor_cse_sva);
  assign or_dcpl_82 = (fsm_output[5]) | (fsm_output[21]);
  assign or_dcpl_83 = (fsm_output[4]) | (fsm_output[20]);
  assign or_dcpl_85 = (fsm_output[5:4]!=2'b00);
  assign or_dcpl_86 = (fsm_output[21:20]!=2'b00);
  assign or_dcpl_87 = (fsm_output[23:22]!=2'b00);
  assign or_dcpl_88 = (fsm_output[7]) | (fsm_output[5]);
  assign or_dcpl_89 = (fsm_output[25:24]!=2'b00);
  assign or_dcpl_92 = (fsm_output[36:35]!=2'b00);
  assign or_dcpl_98 = (fsm_output[25]) | (fsm_output[29]);
  assign or_dcpl_99 = (fsm_output[27:26]!=2'b00);
  assign or_dcpl_101 = (and_dcpl_80 & (operator_16_false_io_read_mode1_rsc_cse_sva[13:0]==14'b00000000000001))
      | operator_16_false_operator_16_false_nor_cse_sva;
  assign or_dcpl_102 = (fsm_output[33:32]!=2'b00);
  assign or_dcpl_104 = (fsm_output[16]) | (fsm_output[14]);
  assign or_dcpl_106 = (fsm_output[10:9]!=2'b00);
  assign or_dcpl_107 = (fsm_output[13:12]!=2'b00);
  assign or_dcpl_109 = (fsm_output[20]) | (fsm_output[22]);
  assign or_dcpl_111 = (fsm_output[21]) | (fsm_output[14]);
  assign and_dcpl_110 = ~((fsm_output[0]) | (fsm_output[38]));
  assign or_dcpl_124 = (fsm_output[26:25]!=2'b00);
  assign or_dcpl_125 = or_dcpl_124 | (fsm_output[29]);
  assign or_dcpl_133 = (fsm_output[15:14]!=2'b00);
  assign or_dcpl_145 = (fsm_output[23]) | (fsm_output[9]);
  assign or_dcpl_147 = (fsm_output[16]) | (fsm_output[13]);
  assign or_dcpl_151 = ~(mode_lpi_1_dfm & inverse_lpi_1_dfm_1);
  assign and_dcpl_112 = (return_add_generic_AC_RND_CONV_false_2_res_rounded_acc_tmp[53])
      & return_add_generic_AC_RND_CONV_false_2_if_5_return_add_generic_AC_RND_CONV_false_2_if_5_and_1_tmp;
  assign or_dcpl_152 = and_dcpl_112 | or_dcpl_151;
  assign or_dcpl_153 = operator_11_true_return_1_sva | operator_11_true_return_13_sva;
  assign or_dcpl_158 = return_add_generic_AC_RND_CONV_false_1_r_inf_lpi_3_dfm_2 |
      operator_11_true_return_1_sva;
  assign or_dcpl_159 = or_dcpl_158 | and_dcpl_112 | operator_11_true_return_13_sva;
  assign and_dcpl_114 = return_add_generic_AC_RND_CONV_false_15_if_5_return_add_generic_AC_RND_CONV_false_15_if_5_and_1_tmp
      & (return_add_generic_AC_RND_CONV_false_res_rounded_acc_tmp[53]);
  assign or_dcpl_164 = return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2 |
      and_dcpl_114;
  assign or_dcpl_167 = return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2 |
      operator_11_true_return_1_sva;
  assign or_dcpl_168 = or_dcpl_167 | and_dcpl_114 | operator_11_true_return_13_sva;
  assign or_dcpl_172 = operator_11_true_return_1_sva | operator_11_true_return_24_sva;
  assign and_dcpl_118 = ~(return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva
      | operator_11_true_return_15_sva);
  assign and_dcpl_121 = (~((~((~ (stage_u_add_3_acc_itm_rsp_1[11])) & return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva)) & (~(return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm
      & (return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[53])));
  assign or_dcpl_183 = operator_11_true_return_15_sva | operator_11_true_return_13_sva;
  assign or_dcpl_190 = operator_11_true_return_13_sva | (~ mode_lpi_1_dfm);
  assign and_dcpl_125 = return_add_generic_AC_RND_CONV_false_20_if_5_return_add_generic_AC_RND_CONV_false_20_if_5_and_1_tmp
      & (return_add_generic_AC_RND_CONV_false_7_res_rounded_acc_tmp[53]);
  assign or_dcpl_193 = return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2 |
      operator_11_true_return_1_sva;
  assign or_dcpl_198 = operator_11_true_return_17_sva | (~ mode_lpi_1_dfm);
  assign and_dcpl_127 = (z_out_46[53]) & return_add_generic_AC_RND_CONV_false_8_if_5_return_add_generic_AC_RND_CONV_false_8_if_5_and_tmp;
  assign or_dcpl_201 = return_add_generic_AC_RND_CONV_false_8_r_inf_lpi_3_dfm_2 |
      operator_11_true_return_13_sva;
  assign and_dcpl_129 = (return_add_generic_AC_RND_CONV_false_19_res_rounded_acc_tmp[53])
      & return_add_generic_AC_RND_CONV_false_19_if_5_return_add_generic_AC_RND_CONV_false_19_if_5_and_tmp;
  assign or_dcpl_212 = return_add_generic_AC_RND_CONV_false_19_r_inf_lpi_3_dfm_2
      | or_dcpl_25;
  assign and_dcpl_131 = return_add_generic_AC_RND_CONV_false_20_if_5_return_add_generic_AC_RND_CONV_false_20_if_5_and_1_tmp
      & (return_add_generic_AC_RND_CONV_false_20_res_rounded_acc_tmp[53]);
  assign and_dcpl_132 = return_add_generic_AC_RND_CONV_false_21_if_5_return_add_generic_AC_RND_CONV_false_21_if_5_and_tmp
      & (return_add_generic_AC_RND_CONV_false_21_res_rounded_acc_tmp[53]);
  assign or_dcpl_238 = (~ mode_lpi_1_dfm) | inverse_lpi_1_dfm_1;
  assign and_dcpl_133 = return_add_generic_AC_RND_CONV_false_22_if_5_return_add_generic_AC_RND_CONV_false_22_if_5_and_1_tmp
      & (z_out_47[53]);
  assign or_dcpl_245 = return_add_generic_AC_RND_CONV_false_9_r_inf_lpi_3_dfm_2 |
      operator_11_true_return_1_sva | and_dcpl_133 | operator_11_true_return_24_sva;
  assign and_dcpl_135 = return_add_generic_AC_RND_CONV_false_10_if_5_return_add_generic_AC_RND_CONV_false_10_if_5_and_tmp
      & (z_out_46[53]);
  assign or_dcpl_250 = operator_11_true_return_13_sva | operator_11_true_return_26_sva;
  assign and_dcpl_136 = (z_out_46[53]) & return_add_generic_AC_RND_CONV_false_11_if_5_return_add_generic_AC_RND_CONV_false_11_if_5_and_tmp;
  assign and_dcpl_139 = return_add_generic_AC_RND_CONV_false_24_if_5_return_add_generic_AC_RND_CONV_false_24_if_5_and_tmp
      & (return_add_generic_AC_RND_CONV_false_24_res_rounded_acc_tmp[53]);
  assign and_dcpl_141 = return_add_generic_AC_RND_CONV_false_25_if_5_return_add_generic_AC_RND_CONV_false_25_if_5_and_tmp
      & (return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp[53]);
  assign and_dcpl_143 = return_add_generic_AC_RND_CONV_false_23_if_5_return_add_generic_AC_RND_CONV_false_23_if_5_and_tmp
      & (return_add_generic_AC_RND_CONV_false_23_res_rounded_acc_tmp[53]);
  assign and_dcpl_147 = ~((fsm_output[1]) | (fsm_output[18]) | (fsm_output[34]));
  assign and_dcpl_149 = ~((fsm_output[1]) | (fsm_output[36]) | (fsm_output[35]));
  assign and_dcpl_150 = and_dcpl_110 & (~ (fsm_output[37]));
  assign and_dcpl_164 = ~((fsm_output[3]) | (fsm_output[19]));
  assign or_dcpl_300 = (fsm_output[9:8]!=2'b00);
  assign or_dcpl_305 = (fsm_output[12:11]!=2'b00);
  assign and_dcpl_170 = ~((fsm_output[2]) | (fsm_output[0]));
  assign and_dcpl_179 = ~((fsm_output[37]) | (fsm_output[1]));
  assign or_dcpl_316 = (fsm_output[22]) | (fsm_output[10]) | return_add_generic_AC_RND_CONV_false_14_or_cse;
  assign or_dcpl_320 = (fsm_output[24]) | (fsm_output[27]);
  assign or_dcpl_325 = (fsm_output[29]) | (fsm_output[13]);
  assign or_dcpl_326 = (fsm_output[32]) | (fsm_output[30]);
  assign or_dcpl_328 = (fsm_output[6]) | (fsm_output[10]) | (fsm_output[7]);
  assign and_dcpl_196 = ~(return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_23_e_dif1_acc_1_tmp[11]));
  assign and_dcpl_197 = ~(operator_11_true_return_13_sva | operator_11_true_return_26_sva);
  assign or_dcpl_338 = (fsm_output[27]) | (fsm_output[11]);
  assign or_dcpl_340 = (fsm_output[31]) | (fsm_output[27]);
  assign or_dcpl_343 = (fsm_output[28]) | (fsm_output[30]);
  assign or_dcpl_352 = or_dcpl_305 | (fsm_output[25]);
  assign or_dcpl_353 = return_add_generic_AC_RND_CONV_false_15_res_mant_or_1_cse
      | (fsm_output[27]);
  assign or_dcpl_354 = or_dcpl_353 | or_dcpl_352;
  assign or_dcpl_356 = ~((({return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0 , return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_1_op2_mu_51_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1})) & return_add_generic_AC_RND_CONV_false_1_e1_eq_e2_equal_tmp);
  assign or_dcpl_357 = ~(return_add_generic_AC_RND_CONV_false_9_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1})));
  assign or_dcpl_358 = ~(return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva & return_add_generic_AC_RND_CONV_false_12_mux_itm);
  assign or_dcpl_359 = ~(return_add_generic_AC_RND_CONV_false_14_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0
      , return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm_1
      , return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm_mx1 , return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1})));
  assign or_dcpl_360 = ~(return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm_mx1
      , return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0 , return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1})));
  assign or_dcpl_361 = ~(return_add_generic_AC_RND_CONV_false_22_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm , return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0
      , return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1})));
  assign or_dcpl_365 = (fsm_output[14]) | (fsm_output[9]);
  assign or_dcpl_367 = (fsm_output[28:27]!=2'b00);
  assign or_dcpl_377 = (fsm_output[25]) | (fsm_output[13]);
  assign or_dcpl_380 = or_dcpl_338 | (fsm_output[12]);
  assign or_dcpl_385 = (fsm_output[24]) | (fsm_output[23]) | (fsm_output[21]);
  assign or_dcpl_387 = (fsm_output[13]) | (fsm_output[6]);
  assign or_dcpl_388 = (fsm_output[12]) | (fsm_output[25]);
  assign or_dcpl_390 = return_add_generic_AC_RND_CONV_false_15_res_mant_or_1_cse
      | (fsm_output[24]);
  assign or_dcpl_396 = (fsm_output[30]) | (fsm_output[24]);
  assign and_dcpl_214 = ~(and_272_cse | (z_out_17[11]));
  assign and_dcpl_215 = ~(and_277_cse | (z_out_18[11]));
  assign and_dcpl_216 = ~(return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_and_1_cse
      | (z_out_18[11]));
  assign and_dcpl_219 = ~(and_275_cse | (return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp[11]));
  assign and_dcpl_220 = ~(and_276_cse | (return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp[11]));
  assign and_dcpl_224 = ~(and_271_cse | (z_out_17[11]));
  assign or_dcpl_432 = (fsm_output[30:29]!=2'b00);
  assign and_dcpl_225 = ~(return_add_generic_AC_RND_CONV_false_4_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_4_op1_smaller_oelse_and_1_cse
      | (return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp[10]));
  assign or_dcpl_436 = (fsm_output[25]) | (fsm_output[15]);
  assign or_dcpl_437 = or_dcpl_99 | (fsm_output[11]);
  assign and_dcpl_226 = ~(return_add_generic_AC_RND_CONV_false_11_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_11_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_9_e_dif1_acc_1_tmp[11]));
  assign and_dcpl_227 = ~(return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_10_e_dif1_acc_1_tmp[11]));
  assign or_dcpl_441 = ~(return_add_generic_AC_RND_CONV_false_22_e1_eq_e2_equal_tmp
      & z_out_2_52);
  assign and_dcpl_228 = or_dcpl_441 & (~ (return_add_generic_AC_RND_CONV_false_22_e_dif1_acc_1_tmp[11]));
  assign or_dcpl_442 = return_add_generic_AC_RND_CONV_false_14_or_cse | or_dcpl_300;
  assign or_dcpl_443 = (fsm_output[25]) | (fsm_output[10]);
  assign and_dcpl_229 = ~((z_out_55[11]) | return_mult_generic_AC_RND_CONV_false_3_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_3_exp_ovf_oif_aelse_and_1_tmp);
  assign and_dcpl_231 = ~(operator_11_true_return_1_sva | operator_11_true_return_15_sva);
  assign or_dcpl_450 = ~(return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_cse_sva
      & return_extract_44_m_zero_sva);
  assign or_dcpl_454 = (fsm_output[25]) | (fsm_output[22]) | (fsm_output[10]);
  assign or_dcpl_456 = or_dcpl_390 | or_dcpl_380;
  assign and_dcpl_241 = ~(return_add_generic_AC_RND_CONV_false_24_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_24_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_22_e_dif1_acc_1_tmp[11]));
  assign or_dcpl_471 = (fsm_output[14:13]!=2'b00);
  assign or_dcpl_474 = ~(return_add_generic_AC_RND_CONV_false_17_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_4_op1_mu_52_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_4_op1_mu_51_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_4_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_4_op2_mu_52_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_4_op2_mu_51_1_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_4_op2_mu_0_lpi_3_dfm_1})));
  assign or_dcpl_475 = (fsm_output[31]) | (fsm_output[25]);
  assign or_dcpl_477 = or_dcpl_326 | (fsm_output[24]) | or_dcpl_475;
  assign or_dcpl_480 = ~(return_add_generic_AC_RND_CONV_false_23_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1})));
  assign or_dcpl_488 = ~(return_add_generic_AC_RND_CONV_false_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_1_op2_mu_51_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0 , return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1})));
  assign or_dcpl_505 = (fsm_output[10]) | (fsm_output[14]) | (fsm_output[15]);
  assign or_dcpl_511 = return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_2_cse
      | (fsm_output[8]);
  assign or_dcpl_523 = (fsm_output[11]) | (fsm_output[25]);
  assign and_dcpl_248 = ~(return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp[11]));
  assign and_dcpl_249 = ~(return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp[11]));
  assign and_dcpl_254 = ~(operator_11_true_return_1_sva | operator_11_true_return_13_sva);
  assign and_dcpl_281 = (~((~(return_add_generic_AC_RND_CONV_false_2_else_4_return_add_generic_AC_RND_CONV_false_2_else_4_nand_tmp
      & (~ (operator_33_true_4_acc_tmp[11])))) & return_add_generic_AC_RND_CONV_false_2_acc_3_itm_11_1))
      & (~((return_add_generic_AC_RND_CONV_false_2_res_rounded_acc_tmp[53]) & return_add_generic_AC_RND_CONV_false_2_if_5_return_add_generic_AC_RND_CONV_false_2_if_5_and_1_tmp));
  assign or_dcpl_551 = (fsm_output[15]) | (fsm_output[9]);
  assign or_dcpl_571 = return_add_generic_AC_RND_CONV_false_15_res_mant_or_1_cse
      | or_dcpl_338;
  assign and_dcpl_294 = ~(operator_11_true_return_1_sva | operator_11_true_return_24_sva);
  assign and_dcpl_300 = ~(operator_11_true_return_13_sva | operator_11_true_return_17_sva
      | return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva);
  assign or_dcpl_597 = ~((~((~ (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_2_1[0]))
      & return_add_generic_AC_RND_CONV_false_21_else_4_return_add_generic_AC_RND_CONV_false_21_else_4_nand_tmp))
      & return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1);
  assign and_dcpl_312 = ~(return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_and_1_cse
      | return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm);
  assign and_dcpl_314 = and_dcpl_118 & (~(operator_11_true_return_13_sva | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva));
  assign and_dcpl_316 = and_dcpl_254 & (~ return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign or_dcpl_625 = ~((~((~ (stage_u_add_3_acc_itm_rsp_1[11])) & return_add_generic_AC_RND_CONV_false_10_else_4_return_add_generic_AC_RND_CONV_false_10_else_4_nand_tmp))
      & return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1);
  assign or_tmp_26 = operator_16_false_operator_16_false_nor_cse_sva & (fsm_output[36]);
  assign and_392_cse = and_dcpl_91 & (fsm_output[36]);
  assign and_421_cse = and_dcpl_85 & or_dcpl_92;
  assign or_tmp_46 = (fsm_output[34]) | ((~ (for_i_3_0_sva[0])) & (fsm_output[2]));
  assign and_448_cse = inverse_lpi_1_dfm_1 & (fsm_output[24]);
  assign and_450_cse = (~ inverse_lpi_1_dfm_1) & (fsm_output[24]);
  assign and_475_cse = inverse_lpi_1_dfm_1 & (fsm_output[30]);
  assign and_477_cse = (~ inverse_lpi_1_dfm_1) & (fsm_output[30]);
  assign and_503_cse = and_dcpl_85 & (fsm_output[35]);
  assign and_537_cse = inverse_lpi_1_dfm_1 & (fsm_output[14]);
  assign and_539_cse = (~ inverse_lpi_1_dfm_1) & (fsm_output[14]);
  assign and_565_cse = return_add_generic_AC_RND_CONV_false_1_r_inf_lpi_3_dfm_2 |
      or_dcpl_153 | or_dcpl_152;
  assign and_569_cse = or_dcpl_164 | or_dcpl_153 | or_dcpl_151;
  assign and_573_cse = (z_out_45[12]) | (~ mode_lpi_1_dfm);
  assign and_631_cse = return_add_generic_AC_RND_CONV_false_9_r_inf_lpi_3_dfm_2 |
      or_dcpl_172 | and_dcpl_133 | or_dcpl_238;
  assign or_tmp_180 = inverse_lpi_1_dfm_1 & (fsm_output[2]);
  assign or_tmp_181 = (~ inverse_lpi_1_dfm_1) & (fsm_output[2]);
  assign or_tmp_388 = return_add_generic_AC_RND_CONV_false_17_op1_smaller_lor_lpi_3_dfm_2
      & (fsm_output[6]);
  assign or_tmp_389 = and_dcpl_225 & (fsm_output[6]);
  assign or_tmp_543 = or_dcpl_353 | or_dcpl_305 | or_dcpl_377 | or_dcpl_106;
  assign or_tmp_567 = (fsm_output[30]) | (fsm_output[14]);
  assign or_tmp_606 = or_dcpl_89 | or_dcpl_300;
  assign and_1747_cse = or_dcpl_436 | (fsm_output[9]);
  assign or_tmp_773 = inverse_lpi_1_dfm_1 & (fsm_output[25]);
  assign out1_rsci_idat_63_0_mx0c1 = and_dcpl_83 & and_dcpl_74 & (operator_16_false_io_read_mode1_rsc_cse_sva[2:0]==3'b001)
      & (~ operator_16_false_operator_16_false_nor_cse_sva) & (fsm_output[36]);
  assign out1_rsci_idat_63_0_mx0c2 = and_dcpl_85 & (fsm_output[36]);
  assign out1_rsci_idat_79_64_mx0c1 = and_dcpl_83 & and_dcpl_74 & (operator_16_false_io_read_mode1_rsc_cse_sva[2:1]==2'b01)
      & (~((operator_16_false_io_read_mode1_rsc_cse_sva[0]) | operator_16_false_operator_16_false_nor_cse_sva))
      & (fsm_output[36]);
  assign out_f_d_rsci_adr_d_mx0c2 = (fsm_output[32]) | (fsm_output[29]) | (fsm_output[6])
      | (fsm_output[35]);
  assign out_f_d_rsci_adr_d_mx0c3 = (fsm_output[25]) | (fsm_output[7]) | and_477_cse;
  assign out_f_d_rsci_adr_d_mx0c5 = (fsm_output[33]) | (fsm_output[31]) | and_475_cse;
  assign in_f_d_rsci_adr_d_mx0c2 = or_dcpl_147 | (fsm_output[22]) | (fsm_output[35]);
  assign BUTTERFLY_1_i_9_0_sva_mx0c3 = or_dcpl_326 | or_dcpl_104;
  assign BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c0 = (~ mode_lpi_1_dfm)
      & (fsm_output[6]);
  assign BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c4 = or_dcpl_432 | (fsm_output[15])
      | (mode_lpi_1_dfm & or_dcpl_35);
  assign BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c7 = (fsm_output[25])
      | and_2638_cse;
  assign drf_qr_lval_10_smx_lpi_3_dfm_mx0c0 = or_dcpl_432 | (fsm_output[16]) | or_dcpl_387
      | (fsm_output[22]) | (fsm_output[7]) | (fsm_output[23]) | or_dcpl_133;
  assign in_u_rsc_merge_sva_mx0c2 = or_dcpl_396 | or_dcpl_475 | or_dcpl_325 | or_dcpl_133
      | (mode_lpi_1_dfm & or_dcpl_300);
  assign or_1478_tmp = in_f_d_rsci_adr_d_mx0c2 | (fsm_output[21]);
  assign or_723_nl = or_dcpl_145 | and_539_cse;
  assign or_726_nl = (fsm_output[17]) | (fsm_output[15]) | and_537_cse;
  assign BUTTERFLY_1_i_mux1h_2_nl = MUX1HOT_s_1_6_2(reg_BUTTERFLY_1_i_9_0_ftd, (~
      reg_BUTTERFLY_1_i_9_0_ftd), (BUTTERFLY_1_fry_9_0_sva[9]), (~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm),
      (~ (BUTTERFLY_i_9_0_sva_1[9])), (~ (BUTTERFLY_1_fry_9_0_sva[9])), {or_723_nl
      , (fsm_output[10]) , in_f_d_rsci_adr_d_mx0c2 , or_726_nl , (fsm_output[20])
      , (fsm_output[21])});
  assign nor_129_nl = ~((fsm_output[20]) | or_1478_tmp);
  assign mux1h_4_nl = MUX1HOT_v_9_3_2(reg_BUTTERFLY_1_i_9_0_ftd_1, (BUTTERFLY_i_9_0_sva_1[8:0]),
      (BUTTERFLY_1_fry_9_0_sva[8:0]), {nor_129_nl , (fsm_output[20]) , or_1478_tmp});
  assign in_f_d_rsci_adr_d = {BUTTERFLY_1_i_mux1h_2_nl , mux1h_4_nl};
  assign BUTTERFLY_if_1_if_and_3_cse = return_add_generic_AC_RND_CONV_false_9_or_1_svs_1
      & and_539_cse;
  assign nor_113_m1c = ~(or_tmp_833 | or_tmp_834 | or_tmp_835);
  assign and_2106_cse = return_add_generic_AC_RND_CONV_false_or_1_svs_1 & (fsm_output[9]);
  assign and_2105_cse = return_add_generic_AC_RND_CONV_false_10_or_1_svs_1 & (fsm_output[15]);
  assign and_2108_cse = return_add_generic_AC_RND_CONV_false_11_or_1_svs_1 & (fsm_output[16]);
  assign and_2107_cse = return_add_generic_AC_RND_CONV_false_12_or_1_svs_1 & (fsm_output[17]);
  assign or_1482_tmp = BUTTERFLY_if_1_if_and_3_cse | and_2105_cse | and_2106_cse
      | and_2107_cse | and_2108_cse;
  assign return_add_generic_AC_RND_CONV_false_10_mux_20_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_and_11,
      return_add_generic_AC_RND_CONV_false_10_exp_plus_1_0_lpi_3_dfm_1, z_out_46[53]);
  assign BUTTERFLY_if_1_if_or_nl = (fsm_output[9]) | (fsm_output[17]);
  assign BUTTERFLY_if_1_if_or_1_nl = (fsm_output[10]) | and_539_cse | (fsm_output[15]);
  assign BUTTERFLY_if_1_if_mux1h_nl = MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_12_mux_itm,
      return_add_generic_AC_RND_CONV_false_10_mux_7_itm, return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1,
      operator_11_true_return_15_sva, return_add_generic_AC_RND_CONV_false_11_mux_itm,
      {BUTTERFLY_if_1_if_or_nl , BUTTERFLY_if_1_if_or_1_nl , (fsm_output[13]) , and_537_cse
      , (fsm_output[16])});
  assign and_2157_nl = (fsm_output[9]) & nor_113_m1c;
  assign and_2158_nl = (fsm_output[10]) & nor_113_m1c;
  assign and_2159_nl = (fsm_output[13]) & nor_113_m1c;
  assign and_2160_nl = and_537_cse & nor_113_m1c;
  assign and_2161_nl = and_539_cse & nor_113_m1c;
  assign or_1732_nl = ((fsm_output[15]) & nor_113_m1c) | ((fsm_output[17]) & nor_113_m1c);
  assign BUTTERFLY_if_1_if_and_10_nl = (~ (z_out_46[53])) & (fsm_output[16]) & nor_113_m1c;
  assign BUTTERFLY_if_1_if_and_11_nl = (z_out_46[53]) & (fsm_output[16]) & nor_113_m1c;
  assign mux1h_1_nl = MUX1HOT_v_10_9_2(return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_itm,
      return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1, ({in_u_rsc_merge_sva_rsp_1_rsp_0
      , in_u_rsc_merge_sva_rsp_1_rsp_1}), return_add_generic_AC_RND_CONV_false_9_e_r_return_add_generic_AC_RND_CONV_false_9_e_r_or_cse,
      (return_add_generic_AC_RND_CONV_false_10_exp_plus_1_12_1_lpi_3_dfm_1[9:0]),
      return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_and_9,
      (return_add_generic_AC_RND_CONV_false_11_exp_plus_1_12_1_lpi_3_dfm_1[9:0]),
      return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_and_9,
      {and_2157_nl , and_2158_nl , and_2159_nl , and_2160_nl , and_2161_nl , or_1732_nl
      , BUTTERFLY_if_1_if_and_10_nl , BUTTERFLY_if_1_if_and_11_nl , or_tmp_834});
  assign not_741_nl = ~ or_tmp_835;
  assign and_2164_nl = MUX_v_10_2_2(10'b0000000000, mux1h_1_nl, not_741_nl);
  assign or_1488_nl = MUX_v_10_2_2(and_2164_nl, 10'b1111111111, or_tmp_833);
  assign or_202_nl = or_dcpl_167 | and_dcpl_114 | operator_11_true_return_24_sva;
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_3_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs, or_202_nl);
  assign return_add_generic_AC_RND_CONV_false_e_r_return_add_generic_AC_RND_CONV_false_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_3_mux_26 & (~ return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_3_nl))
      | return_add_generic_AC_RND_CONV_false_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_22_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs, or_dcpl_245);
  assign return_add_generic_AC_RND_CONV_false_9_e_r_return_add_generic_AC_RND_CONV_false_9_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_9_mux_35 & (~ return_add_generic_AC_RND_CONV_false_22_e_r_qelse_mux_1_nl))
      | return_add_generic_AC_RND_CONV_false_9_exception_sva_1;
  assign or_281_nl = return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2 | operator_11_true_return_13_sva
      | and_dcpl_135 | operator_11_true_return_26_sva;
  assign return_add_generic_AC_RND_CONV_false_10_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs, or_281_nl);
  assign return_add_generic_AC_RND_CONV_false_10_e_r_return_add_generic_AC_RND_CONV_false_10_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_10_mux_20_cse & (~ return_add_generic_AC_RND_CONV_false_10_e_r_qelse_mux_1_nl))
      | return_add_generic_AC_RND_CONV_false_10_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_11_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_and_11,
      return_add_generic_AC_RND_CONV_false_11_exp_plus_1_0_lpi_3_dfm_1, z_out_46[53]);
  assign or_292_nl = return_add_generic_AC_RND_CONV_false_11_r_inf_lpi_3_dfm_2 |
      or_dcpl_172 | and_dcpl_136 | operator_11_true_return_17_sva | return_add_generic_AC_RND_CONV_false_15_do_sub_sva;
  assign return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs, or_292_nl);
  assign return_add_generic_AC_RND_CONV_false_11_e_r_return_add_generic_AC_RND_CONV_false_11_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_11_mux_13_nl & (~ return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_1_nl))
      | return_add_generic_AC_RND_CONV_false_11_exception_sva_1;
  assign or_300_nl = return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2 | or_dcpl_25
      | or_dcpl_183 | and_dcpl_135;
  assign return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs, or_300_nl);
  assign return_add_generic_AC_RND_CONV_false_12_e_r_return_add_generic_AC_RND_CONV_false_12_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_10_mux_20_cse & (~ return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_1_nl))
      | return_add_generic_AC_RND_CONV_false_12_exception_sva_1;
  assign BUTTERFLY_if_1_if_or_2_nl = (fsm_output[10]) | and_537_cse;
  assign BUTTERFLY_if_1_if_mux1h_2_nl = MUX1HOT_s_1_7_2(return_add_generic_AC_RND_CONV_false_e_r_return_add_generic_AC_RND_CONV_false_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm,
      return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_9_e_r_return_add_generic_AC_RND_CONV_false_9_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_10_e_r_return_add_generic_AC_RND_CONV_false_10_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_11_e_r_return_add_generic_AC_RND_CONV_false_11_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_12_e_r_return_add_generic_AC_RND_CONV_false_12_e_r_or_1_nl,
      {(fsm_output[9]) , BUTTERFLY_if_1_if_or_2_nl , (fsm_output[13]) , and_539_cse
      , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
  assign return_add_generic_AC_RND_CONV_false_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_15_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_9_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_9_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op1_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_9_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_7_op1_inf_sva_1 & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva);
  assign return_add_generic_AC_RND_CONV_false_10_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_10_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_11_r_nan_or_nl = operator_11_true_return_17_sva
      | return_add_generic_AC_RND_CONV_false_15_do_sub_sva | (operator_11_true_return_1_sva
      & operator_11_true_return_24_sva & return_add_generic_AC_RND_CONV_false_13_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_12_r_nan_or_nl = operator_11_true_return_15_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | (operator_11_true_return_13_sva
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva & return_add_generic_AC_RND_CONV_false_12_do_sub_sva);
  assign BUTTERFLY_if_1_if_and_nl = (~ return_add_generic_AC_RND_CONV_false_or_1_svs_1)
      & (fsm_output[9]);
  assign BUTTERFLY_if_1_if_and_2_nl = (~ return_add_generic_AC_RND_CONV_false_9_or_1_svs_1)
      & and_539_cse;
  assign BUTTERFLY_if_1_if_or_3_nl = ((~ return_add_generic_AC_RND_CONV_false_10_or_1_svs_1)
      & (fsm_output[15])) | ((~ return_add_generic_AC_RND_CONV_false_11_or_1_svs_1)
      & (fsm_output[16])) | ((~ return_add_generic_AC_RND_CONV_false_12_or_1_svs_1)
      & (fsm_output[17]));
  assign BUTTERFLY_if_1_if_mux1h_3_nl = MUX1HOT_s_1_11_2((return_add_generic_AC_RND_CONV_false_3_res_rounded_lpi_3_dfm_51_0_1[51]),
      return_add_generic_AC_RND_CONV_false_r_nan_or_nl, drf_qr_lval_12_smx_0_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm,
      (return_add_generic_AC_RND_CONV_false_4_res_rounded_lpi_3_dfm_51_0_1[51]),
      return_add_generic_AC_RND_CONV_false_9_r_nan_or_nl, (return_add_generic_AC_RND_CONV_false_5_res_rounded_lpi_3_dfm_51_0_1[51]),
      return_add_generic_AC_RND_CONV_false_10_r_nan_or_nl, return_add_generic_AC_RND_CONV_false_11_r_nan_or_nl,
      return_add_generic_AC_RND_CONV_false_12_r_nan_or_nl, {BUTTERFLY_if_1_if_and_nl
      , and_2106_cse , (fsm_output[10]) , (fsm_output[13]) , and_537_cse , BUTTERFLY_if_1_if_and_2_nl
      , BUTTERFLY_if_1_if_and_3_cse , BUTTERFLY_if_1_if_or_3_nl , and_2105_cse ,
      and_2108_cse , and_2107_cse});
  assign and_2166_nl = (fsm_output[9]) & (~ or_1482_tmp);
  assign and_2167_nl = (fsm_output[10]) & (~ or_1482_tmp);
  assign and_2168_nl = (fsm_output[13]) & (~ or_1482_tmp);
  assign and_2169_nl = and_537_cse & (~ or_1482_tmp);
  assign and_2170_nl = and_539_cse & (~ or_1482_tmp);
  assign or_1733_nl = ((fsm_output[15]) & (~ or_1482_tmp)) | ((fsm_output[16]) &
      (~ or_1482_tmp)) | ((fsm_output[17]) & (~ or_1482_tmp));
  assign mux1h_5_nl = MUX1HOT_v_51_6_2((return_add_generic_AC_RND_CONV_false_3_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm,
      return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0,
      (return_add_generic_AC_RND_CONV_false_4_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      (return_add_generic_AC_RND_CONV_false_5_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      {and_2166_nl , and_2167_nl , and_2168_nl , and_2169_nl , and_2170_nl , or_1733_nl});
  assign not_742_nl = ~ or_1482_tmp;
  assign and_2165_nl = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      mux1h_5_nl, not_742_nl);
  assign in_f_d_rsci_d_d = {BUTTERFLY_if_1_if_mux1h_nl , or_1488_nl , BUTTERFLY_if_1_if_mux1h_2_nl
      , BUTTERFLY_if_1_if_mux1h_3_nl , and_2165_nl};
  assign in_f_d_rsci_we_d_pff = (and_dcpl_1 & ((fsm_output[17:15]!=3'b000))) | (stage_PE_1_and_1_tmp
      & ((fsm_output[13]) | (fsm_output[10]) | (fsm_output[9]))) | (mode_lpi_1_dfm
      & (fsm_output[14]));
  assign in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = (mode_lpi_1_dfm & (or_dcpl_109
      | (fsm_output[23]) | (fsm_output[21]))) | and_503_cse;
  assign BUTTERFLY_1_i_or_3_cse = (inverse_lpi_1_dfm_1 & (fsm_output[20])) | ((~
      inverse_lpi_1_dfm_1) & (fsm_output[20]));
  assign BUTTERFLY_1_i_mux1h_1_nl = MUX1HOT_s_1_3_2(reg_BUTTERFLY_1_i_9_0_ftd, (BUTTERFLY_1_fry_9_0_sva[9]),
      (z_out_27[9]), {or_709_ssc , or_710_ssc , BUTTERFLY_1_i_or_3_cse});
  assign BUTTERFLY_1_i_mux1h_7_nl = MUX1HOT_v_9_3_2(reg_BUTTERFLY_1_i_9_0_ftd_1,
      (BUTTERFLY_1_fry_9_0_sva[8:0]), (z_out_27[8:0]), {or_709_ssc , or_710_ssc ,
      BUTTERFLY_1_i_or_3_cse});
  assign in_u_rsci_adr_d = {BUTTERFLY_1_i_mux1h_1_nl , BUTTERFLY_1_i_mux1h_7_nl};
  assign BUTTERFLY_else_1_if_or_nl = (fsm_output[9]) | (fsm_output[14]) | (fsm_output[15]);
  assign in_u_rsci_d_d = MUX1HOT_v_16_3_2(z_out_59, (z_out_58[15:0]), ({{1{stage_monty_mul_acc_2_psp_sva_1[14]}},
      stage_monty_mul_acc_2_psp_sva_1}), {BUTTERFLY_else_1_if_or_nl , (fsm_output[12])
      , (fsm_output[36])});
  assign in_u_rsci_we_d_pff = (and_dcpl_35 & or_dcpl_133) | (stage_PE_1_and_cse &
      ((fsm_output[12]) | (fsm_output[9]))) | and_392_cse;
  assign in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = and_503_cse | ((~ mode_lpi_1_dfm)
      & or_dcpl_86);
  assign or_1483_tmp = out_f_d_rsci_adr_d_mx0c2 | (fsm_output[5]);
  assign BUTTERFLY_if_1_or_9_tmp = out_f_d_rsci_adr_d_mx0c3 | (fsm_output[26]) |
      out_f_d_rsci_adr_d_mx0c5;
  assign BUTTERFLY_if_1_mux1h_2_nl = MUX1HOT_s_1_6_2((~ (BUTTERFLY_i_9_0_sva_1[9])),
      (~ (BUTTERFLY_1_fry_9_0_sva[9])), (BUTTERFLY_1_fry_9_0_sva[9]), reg_BUTTERFLY_1_i_9_0_ftd,
      (~ reg_BUTTERFLY_1_i_9_0_ftd), (~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm),
      {(fsm_output[4]) , (fsm_output[5]) , out_f_d_rsci_adr_d_mx0c2 , out_f_d_rsci_adr_d_mx0c3
      , (fsm_output[26]) , out_f_d_rsci_adr_d_mx0c5});
  assign nor_130_nl = ~(BUTTERFLY_if_1_or_9_tmp | or_1483_tmp);
  assign mux1h_6_nl = MUX1HOT_v_9_3_2((BUTTERFLY_i_9_0_sva_1[8:0]), reg_BUTTERFLY_1_i_9_0_ftd_1,
      (BUTTERFLY_1_fry_9_0_sva[8:0]), {nor_130_nl , BUTTERFLY_if_1_or_9_tmp , or_1483_tmp});
  assign out_f_d_rsci_adr_d = {BUTTERFLY_if_1_mux1h_2_nl , mux1h_6_nl};
  assign BUTTERFLY_if_1_and_5_cse = return_add_generic_AC_RND_CONV_false_22_or_1_svs_1
      & and_477_cse;
  assign or_1484_tmp = (and_477_cse & return_add_generic_AC_RND_CONV_false_22_exception_sva_1)
      | (return_add_generic_AC_RND_CONV_false_13_exception_sva_1 & (fsm_output[25]));
  assign and_2114_cse = return_add_generic_AC_RND_CONV_false_13_or_1_svs_1 & (fsm_output[25]);
  assign or_1485_tmp = BUTTERFLY_if_1_and_5_cse | and_2114_cse;
  assign BUTTERFLY_if_1_or_nl = (fsm_output[25]) | and_477_cse;
  assign BUTTERFLY_if_1_mux1h_1_nl = MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_10_mux_7_itm,
      return_add_generic_AC_RND_CONV_false_11_mux_itm, return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1,
      operator_11_true_return_15_sva, return_add_generic_AC_RND_CONV_false_12_mux_itm,
      return_add_generic_AC_RND_CONV_false_17_mux_6_itm, {BUTTERFLY_if_1_or_nl ,
      BUTTERFLY_if_1_or_1_cse , (fsm_output[29]) , and_475_cse , (fsm_output[32])
      , (fsm_output[33])});
  assign and_2176_nl = (fsm_output[25]) & (~ or_1484_tmp);
  assign or_1491_nl = (fsm_output[26]) | and_475_cse | (fsm_output[33]);
  assign and_2179_nl = and_477_cse & (~ or_1484_tmp);
  assign mux1h_7_nl = MUX1HOT_v_10_5_2(return_add_generic_AC_RND_CONV_false_1_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_itm,
      return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_9_e_r_return_add_generic_AC_RND_CONV_false_9_e_r_or_cse,
      ({in_u_rsc_merge_sva_rsp_1_rsp_0 , in_u_rsc_merge_sva_rsp_1_rsp_1}), {and_2176_nl
      , or_1491_nl , (fsm_output[29]) , and_2179_nl , BUTTERFLY_if_1_or_3_cse});
  assign or_1489_nl = MUX_v_10_2_2(mux1h_7_nl, 10'b1111111111, or_1484_tmp);
  assign return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_7_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs, or_dcpl_159);
  assign return_add_generic_AC_RND_CONV_false_13_e_r_return_add_generic_AC_RND_CONV_false_13_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_32 & (~ return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_7_nl))
      | return_add_generic_AC_RND_CONV_false_13_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_22_e_r_qelse_mux_3_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs, or_dcpl_245);
  assign return_add_generic_AC_RND_CONV_false_22_e_r_return_add_generic_AC_RND_CONV_false_22_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_9_mux_35 & (~ return_add_generic_AC_RND_CONV_false_22_e_r_qelse_mux_3_nl))
      | return_add_generic_AC_RND_CONV_false_22_exception_sva_1;
  assign BUTTERFLY_if_1_or_4_nl = (fsm_output[26]) | and_475_cse;
  assign BUTTERFLY_if_1_mux1h_7_nl = MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_13_e_r_return_add_generic_AC_RND_CONV_false_13_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm,
      return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_22_e_r_return_add_generic_AC_RND_CONV_false_22_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_and_1_itm,
      return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm,
      {(fsm_output[25]) , BUTTERFLY_if_1_or_4_nl , (fsm_output[29]) , and_477_cse
      , BUTTERFLY_if_1_or_3_cse , (fsm_output[33])});
  assign return_add_generic_AC_RND_CONV_false_13_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_7_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_7_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_13_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_22_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_22_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_22_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1 & return_add_generic_AC_RND_CONV_false_15_do_sub_sva);
  assign BUTTERFLY_if_1_and_2_nl = (~ return_add_generic_AC_RND_CONV_false_13_or_1_svs_1)
      & (fsm_output[25]);
  assign BUTTERFLY_if_1_and_4_nl = (~ return_add_generic_AC_RND_CONV_false_22_or_1_svs_1)
      & and_477_cse;
  assign BUTTERFLY_if_1_mux1h_8_nl = MUX1HOT_s_1_9_2((return_add_generic_AC_RND_CONV_false_1_res_rounded_lpi_3_dfm_51_0_1[51]),
      return_add_generic_AC_RND_CONV_false_13_r_nan_or_nl, drf_qr_lval_12_smx_0_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm,
      (return_add_generic_AC_RND_CONV_false_4_res_rounded_lpi_3_dfm_51_0_1[51]),
      return_add_generic_AC_RND_CONV_false_22_r_nan_or_nl, drf_qr_lval_14_smx_0_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm, {BUTTERFLY_if_1_and_2_nl
      , and_2114_cse , BUTTERFLY_if_1_or_1_cse , (fsm_output[29]) , and_475_cse ,
      BUTTERFLY_if_1_and_4_nl , BUTTERFLY_if_1_and_5_cse , (fsm_output[32]) , (fsm_output[33])});
  assign and_2182_nl = (fsm_output[25]) & (~ or_1485_tmp);
  assign or_1492_nl = and_475_cse | (fsm_output[33]);
  assign and_2186_nl = and_477_cse & (~ or_1485_tmp);
  assign mux1h_8_nl = MUX1HOT_v_51_6_2((return_add_generic_AC_RND_CONV_false_1_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm,
      return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0,
      (return_add_generic_AC_RND_CONV_false_4_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0, {and_2182_nl , BUTTERFLY_if_1_or_1_cse
      , (fsm_output[29]) , or_1492_nl , and_2186_nl , (fsm_output[32])});
  assign not_746_nl = ~ or_1485_tmp;
  assign and_2181_nl = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      mux1h_8_nl, not_746_nl);
  assign out_f_d_rsci_d_d = {BUTTERFLY_if_1_mux1h_1_nl , or_1489_nl , BUTTERFLY_if_1_mux1h_7_nl
      , BUTTERFLY_if_1_mux1h_8_nl , and_2181_nl};
  assign out_f_d_rsci_we_d_pff = (and_dcpl_1 & (or_dcpl_102 | (fsm_output[31])))
      | (stage_PE_1_and_1_tmp & or_dcpl_125) | (mode_lpi_1_dfm & (fsm_output[30]));
  assign out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = (mode_lpi_1_dfm & ((fsm_output[4])
      | (fsm_output[6]) | or_dcpl_88)) | (or_dcpl_101 & (fsm_output[35]));
  assign BUTTERFLY_1_i_mux1h_nl = MUX1HOT_s_1_3_2(reg_BUTTERFLY_1_i_9_0_ftd, (BUTTERFLY_mux_5_itm_9_0[9]),
      (BUTTERFLY_1_fry_9_0_sva[9]), {or_683_ssc , (fsm_output[6]) , or_685_ssc});
  assign BUTTERFLY_1_i_mux1h_8_nl = MUX1HOT_v_9_3_2(reg_BUTTERFLY_1_i_9_0_ftd_1,
      (BUTTERFLY_mux_5_itm_9_0[8:0]), (BUTTERFLY_1_fry_9_0_sva[8:0]), {or_683_ssc
      , (fsm_output[6]) , or_685_ssc});
  assign out_u_rsci_adr_d = {BUTTERFLY_1_i_mux1h_nl , BUTTERFLY_1_i_mux1h_8_nl};
  assign BUTTERFLY_else_1_if_mux1h_1_nl = MUX1HOT_v_3_4_2((BUTTERFLY_1_else_1_if_acc_1_sdt[15:13]),
      (z_out_58[15:13]), (z_out_59[15:13]), reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd,
      {(fsm_output[22]) , and_448_cse , and_450_cse , (fsm_output[25])});
  assign BUTTERFLY_else_1_if_mux1h_7_nl = MUX1HOT_v_2_4_2((BUTTERFLY_1_else_1_if_acc_1_sdt[12:11]),
      (z_out_58[12:11]), (z_out_59[12:11]), reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_2_1,
      {(fsm_output[22]) , and_448_cse , and_450_cse , (fsm_output[25])});
  assign BUTTERFLY_else_1_if_mux1h_8_nl = MUX1HOT_s_1_4_2((BUTTERFLY_1_else_1_if_acc_1_sdt[10]),
      (z_out_58[10]), (z_out_59[10]), reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0,
      {(fsm_output[22]) , and_448_cse , and_450_cse , (fsm_output[25])});
  assign BUTTERFLY_else_1_if_mux1h_9_nl = MUX1HOT_v_10_4_2((BUTTERFLY_1_else_1_if_acc_1_sdt[9:0]),
      (z_out_58[9:0]), (z_out_59[9:0]), ({reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0
      , reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1}), {(fsm_output[22])
      , and_448_cse , and_450_cse , (fsm_output[25])});
  assign out_u_rsci_d_d = {BUTTERFLY_else_1_if_mux1h_1_nl , BUTTERFLY_else_1_if_mux1h_7_nl
      , BUTTERFLY_else_1_if_mux1h_8_nl , BUTTERFLY_else_1_if_mux1h_9_nl};
  assign out_u_rsci_we_d_pff = (and_dcpl_35 & (fsm_output[25])) | (stage_PE_1_and_cse
      & (fsm_output[22])) | ((~ mode_lpi_1_dfm) & (fsm_output[24]));
  assign out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = (operator_16_false_operator_16_false_nor_cse_sva
      & (fsm_output[35])) | (~(mode_lpi_1_dfm | (~((fsm_output[6:5]!=2'b00)))));
  assign or_dcpl_629 = (~((~(and_1143_ssc | and_1141_ssc)) | return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10))
      | (and_1149_ssc & (~ return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11));
  assign or_tmp = ((~ return_add_generic_AC_RND_CONV_false_21_unequal_tmp) & return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs
      & (fsm_output[31])) | ((~((~ return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs_mx0w0)
      | return_add_generic_AC_RND_CONV_false_23_exception_sva_1)) & (fsm_output[30]));
  assign or_tmp_829 = (return_add_generic_AC_RND_CONV_false_21_unequal_tmp & (fsm_output[31]))
      | (return_add_generic_AC_RND_CONV_false_23_exception_sva_1 & (fsm_output[30]));
  assign or_tmp_830 = ((~ return_mult_generic_AC_RND_CONV_false_5_zero_m_return_mult_generic_AC_RND_CONV_false_5_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_5_r_zero_return_mult_generic_AC_RND_CONV_false_5_r_zero_nor_mdf_sva_1)
      & (fsm_output[27])) | ((~ return_mult_generic_AC_RND_CONV_false_2_zero_m_return_mult_generic_AC_RND_CONV_false_2_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_2_r_zero_return_mult_generic_AC_RND_CONV_false_2_r_zero_nor_mdf_sva_1)
      & (fsm_output[11]));
  assign or_tmp_833 = (and_539_cse & return_add_generic_AC_RND_CONV_false_9_exception_sva_1)
      | (return_add_generic_AC_RND_CONV_false_10_exception_sva_1 & (fsm_output[15]))
      | (return_add_generic_AC_RND_CONV_false_exception_sva_1 & (fsm_output[9]))
      | (return_add_generic_AC_RND_CONV_false_12_exception_sva_1 & (fsm_output[17]))
      | (return_add_generic_AC_RND_CONV_false_11_exception_sva_1 & (fsm_output[16]));
  assign or_tmp_834 = ((~(return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs_mx0w0
      | (z_out_46[53]) | return_add_generic_AC_RND_CONV_false_10_exception_sva_1))
      & (fsm_output[15])) | ((~(return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs_mx0w0
      | (z_out_46[53]) | return_add_generic_AC_RND_CONV_false_12_exception_sva_1))
      & (fsm_output[17]));
  assign or_tmp_835 = (return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs_mx0w0
      & (~ return_add_generic_AC_RND_CONV_false_10_exception_sva_1) & (fsm_output[15]))
      | (return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs_mx0w0 & (~ return_add_generic_AC_RND_CONV_false_12_exception_sva_1)
      & (fsm_output[17])) | ((~ return_add_generic_AC_RND_CONV_false_11_exception_sva_1)
      & return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w0 & (fsm_output[16]));
  assign or_1342_ssc = and_1747_cse | and_1804_cse;
  assign or_1344_ssc = and_1808_cse | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_11_cse;
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_and_cse = (~ (return_add_generic_AC_RND_CONV_false_23_res_rounded_acc_tmp[53]))
      & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_and_1_cse = (return_add_generic_AC_RND_CONV_false_23_res_rounded_acc_tmp[53])
      & (fsm_output[30]);
  assign stage_PE_tmp_im_d_and_cse = (~ return_mult_generic_AC_RND_CONV_false_2_e_incr_lpi_3_dfm_2)
      & (fsm_output[11]);
  assign stage_PE_tmp_im_d_and_2_cse = (~ return_mult_generic_AC_RND_CONV_false_5_e_incr_lpi_3_dfm_2)
      & (fsm_output[27]);
  assign and_2189_nl = (z_out_47[53]) & (~ return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs_mx0w0);
  assign mux_18_nl = MUX_v_10_2_2((operator_33_true_44_acc_tmp[10:1]), (return_add_generic_AC_RND_CONV_false_9_exp_plus_1_12_1_lpi_3_dfm_1[9:0]),
      and_2189_nl);
  assign not_748_nl = ~ return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs_mx0w0;
  assign return_add_generic_AC_RND_CONV_false_9_e_r_return_add_generic_AC_RND_CONV_false_9_e_r_or_cse
      = MUX_v_10_2_2(10'b0000000000, mux_18_nl, not_748_nl);
  assign or_1495_cse_1 = (fsm_output[8]) | (fsm_output[24]);
  assign or_1531_cse = (fsm_output[7]) | (fsm_output[9]) | (fsm_output[25]) | (fsm_output[23]);
  assign or_1556_cse = (fsm_output[26]) | (fsm_output[10]);
  assign or_tmp_900 = return_add_generic_AC_RND_CONV_false_12_do_sub_sva & or_1556_cse;
  assign or_tmp_920 = inverse_lpi_1_dfm_1 & or_dcpl_83;
  assign or_tmp_1003 = (fsm_output[19:18]!=2'b00);
  assign or_tmp_1041 = ~(inverse_lpi_1_dfm_1 | (~((fsm_output[4]) | (fsm_output[20]))));
  assign return_add_generic_AC_RND_CONV_false_10_e_dif_sat_conc_4_itm_4_1 = MUX_v_4_2_2((reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0[3:0]),
      (return_add_generic_AC_RND_CONV_false_20_ls_sva[5:2]), return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_10_res_mant_or_9_cse = return_add_generic_AC_RND_CONV_false_15_res_mant_or_cse
      | or_dcpl_325;
  assign in_u_and_ssc = run_wen & ((fsm_output[7]) | (fsm_output[10]) | in_u_rsc_merge_sva_mx0c2
      | (fsm_output[21]) | (fsm_output[23]));
  assign stage_PE_tmp_im_d_or_cse = (return_mult_generic_AC_RND_CONV_false_2_e_incr_lpi_3_dfm_2
      & (fsm_output[11])) | (return_mult_generic_AC_RND_CONV_false_5_e_incr_lpi_3_dfm_2
      & (fsm_output[27]));
  assign operator_6_false_18_and_1_ssc = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_1_cse
      & (~ or_tmp_606);
  assign stage_u_add_3_and_ssc = run_wen & (~ (fsm_output[23]));
  assign stage_u_add_3_or_1_cse = (fsm_output[13]) | or_1367_cse;
  assign return_add_generic_AC_RND_CONV_false_4_res_mant_conc_2_itm_56_1 = MUX_v_56_2_2((z_out_31[56:1]),
      (~ (z_out_31[56:1])), return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign nl_operator_6_false_8_operator_6_false_8_conc_itm_6_1 = ({1'b1 , (~ return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_0)
      , (~ return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_1) , (~ (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2[3:1]))})
      + 6'b000001;
  assign operator_6_false_8_operator_6_false_8_conc_itm_6_1 = nl_operator_6_false_8_operator_6_false_8_conc_itm_6_1[5:0];
  assign return_add_generic_AC_RND_CONV_false_10_exp_conc_5_itm_10_7 = MUX_v_4_2_2(in_u_rsc_merge_sva_rsp_1_rsp_0,
      (stage_PE_1_x_im_d_sva[62:59]), and_dcpl_227);
  assign return_add_generic_AC_RND_CONV_false_10_exp_conc_5_itm_6_1 = MUX_v_6_2_2(in_u_rsc_merge_sva_rsp_1_rsp_1,
      (stage_PE_1_x_im_d_sva[58:53]), and_dcpl_227);
  assign return_add_generic_AC_RND_CONV_false_24_mux_4_itm_5_1 = MUX_v_5_2_2((return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_itm[4:0]),
      (leading_sign_57_0_1_0_24_out_3[5:1]), return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11);
  assign return_add_generic_AC_RND_CONV_false_23_mux_11_itm_5_2 = MUX_v_4_2_2((reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0[3:0]),
      (leading_sign_57_0_1_0_15_out_3[5:2]), return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1);
  assign for_or_4_cse = (fsm_output[8]) | (fsm_output[16]);
  assign for_or_10_cse_1 = (fsm_output[15]) | (fsm_output[17]);
  assign return_mult_generic_AC_RND_CONV_false_2_else_1_nor_cse = ~((fsm_output[11])
      | (fsm_output[27]));
  assign return_add_generic_AC_RND_CONV_false_5_res_rounded_or_1_cse = (fsm_output[13])
      | (fsm_output[15]) | (fsm_output[16]) | (fsm_output[17]);
  assign for_or_5_cse = (fsm_output[16]) | (fsm_output[30]);
  assign BUTTERFLY_else_2_mux_1_cse = MUX_s_1_2_2((stage_u_add_3_acc_itm_rsp_0[3]),
      (z_out_1[16]), fsm_output[24]);
  assign BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_1_cse = MUX_s_1_2_2((z_out_60[17]),
      (z_out_61[17]), or_dcpl_551);
  assign BUTTERFLY_else_1_if_mux_4_cse = MUX_v_3_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd,
      (in_u_rsci_q_d[15:13]), fsm_output[22]);
  assign BUTTERFLY_else_1_if_mux_5_cse = MUX_v_2_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_2_1,
      (in_u_rsci_q_d[12:11]), fsm_output[22]);
  assign BUTTERFLY_else_1_if_mux_6_cse = MUX_s_1_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0,
      (in_u_rsci_q_d[10]), fsm_output[22]);
  assign BUTTERFLY_else_1_if_mux_7_cse_9_1 = MUX_v_9_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0,
      (in_u_rsci_q_d[9:1]), fsm_output[22]);
  assign BUTTERFLY_else_1_if_mux_7_cse_0 = MUX_s_1_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1,
      (in_u_rsci_q_d[0]), fsm_output[22]);
  assign return_add_generic_AC_RND_CONV_false_3_and_20_cse = (~ return_add_generic_AC_RND_CONV_false_25_op1_smaller_return_add_generic_AC_RND_CONV_false_25_op1_smaller_or_cse)
      & (fsm_output[29]);
  assign return_mult_generic_AC_RND_CONV_false_1_else_1_or_cse = (fsm_output[24])
      | or_1556_cse;
  assign return_add_generic_AC_RND_CONV_false_3_and_cse = (~ return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1)
      & (fsm_output[6]);
  assign return_add_generic_AC_RND_CONV_false_3_and_1_cse = return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1
      & (fsm_output[6]);
  assign return_add_generic_AC_RND_CONV_false_3_and_2_cse = (~ return_add_generic_AC_RND_CONV_false_do_sub_sva_1)
      & (fsm_output[8]);
  assign return_add_generic_AC_RND_CONV_false_3_and_3_cse = return_add_generic_AC_RND_CONV_false_do_sub_sva_1
      & (fsm_output[8]);
  assign return_add_generic_AC_RND_CONV_false_3_and_4_cse = (~ return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1)
      & (fsm_output[22]);
  assign return_add_generic_AC_RND_CONV_false_3_and_5_cse = return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1
      & (fsm_output[22]);
  assign return_add_generic_AC_RND_CONV_false_3_and_6_cse = (~ return_add_generic_AC_RND_CONV_false_13_do_sub_sva_1)
      & (fsm_output[24]);
  assign return_add_generic_AC_RND_CONV_false_3_and_7_cse = return_add_generic_AC_RND_CONV_false_13_do_sub_sva_1
      & (fsm_output[24]);
  assign return_add_generic_AC_RND_CONV_false_3_and_8_cse = (~ return_add_generic_AC_RND_CONV_false_10_op2_inf_sva)
      & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_3_and_9_cse = return_add_generic_AC_RND_CONV_false_10_op2_inf_sva
      & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_1_and_8_cse = (~ return_add_generic_AC_RND_CONV_false_10_op2_inf_sva)
      & (fsm_output[13]);
  assign return_add_generic_AC_RND_CONV_false_1_and_9_cse = return_add_generic_AC_RND_CONV_false_10_op2_inf_sva
      & (fsm_output[13]);
  assign return_add_generic_AC_RND_CONV_false_1_and_14_cse = (~ return_add_generic_AC_RND_CONV_false_15_do_sub_sva)
      & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_1_and_15_cse = return_add_generic_AC_RND_CONV_false_15_do_sub_sva
      & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_1_and_28_cse = (~ return_add_generic_AC_RND_CONV_false_11_op1_smaller_return_add_generic_AC_RND_CONV_false_11_op1_smaller_or_cse)
      & (fsm_output[13]);
  assign return_add_generic_AC_RND_CONV_false_1_and_30_cse = (~ return_add_generic_AC_RND_CONV_false_24_op1_smaller_return_add_generic_AC_RND_CONV_false_24_op1_smaller_or_cse)
      & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_11_and_1_cse = (~ return_add_generic_AC_RND_CONV_false_10_do_sub_sva)
      & (fsm_output[26]);
  assign return_add_generic_AC_RND_CONV_false_11_and_2_cse = return_add_generic_AC_RND_CONV_false_10_do_sub_sva
      & (fsm_output[26]);
  assign return_add_generic_AC_RND_CONV_false_11_and_3_cse = (~ return_add_generic_AC_RND_CONV_false_12_mux_itm)
      & (fsm_output[28]);
  assign return_add_generic_AC_RND_CONV_false_11_and_4_cse = return_add_generic_AC_RND_CONV_false_12_mux_itm
      & (fsm_output[28]);
  assign return_add_generic_AC_RND_CONV_false_11_and_11_cse = (~ return_add_generic_AC_RND_CONV_false_19_op1_smaller_lor_lpi_3_dfm_2)
      & (fsm_output[26]);
  assign return_add_generic_AC_RND_CONV_false_11_and_13_cse = (~ or_450_cse) & (fsm_output[28]);
  assign return_add_generic_AC_RND_CONV_false_11_or_cse = return_add_generic_AC_RND_CONV_false_11_and_11_cse
      | return_add_generic_AC_RND_CONV_false_11_and_13_cse;
  assign return_add_generic_AC_RND_CONV_false_11_and_12_cse = return_add_generic_AC_RND_CONV_false_19_op1_smaller_lor_lpi_3_dfm_2
      & (fsm_output[26]);
  assign return_add_generic_AC_RND_CONV_false_3_or_4_cse = return_add_generic_AC_RND_CONV_false_3_and_cse
      | return_add_generic_AC_RND_CONV_false_3_and_3_cse | return_add_generic_AC_RND_CONV_false_3_and_4_cse
      | return_add_generic_AC_RND_CONV_false_3_and_6_cse;
  assign return_add_generic_AC_RND_CONV_false_3_or_5_cse = return_add_generic_AC_RND_CONV_false_3_and_1_cse
      | return_add_generic_AC_RND_CONV_false_3_and_2_cse | return_add_generic_AC_RND_CONV_false_3_and_5_cse
      | return_add_generic_AC_RND_CONV_false_3_and_7_cse;
  assign return_add_generic_AC_RND_CONV_false_3_and_30_cse = (~ return_add_generic_AC_RND_CONV_false_1_op1_smaller_lor_lpi_3_dfm_2)
      & (fsm_output[6]);
  assign return_add_generic_AC_RND_CONV_false_3_and_32_cse = (~ or_452_cse) & (fsm_output[22]);
  assign return_add_generic_AC_RND_CONV_false_5_and_7_cse = return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1
      & (fsm_output[15]);
  assign return_add_generic_AC_RND_CONV_false_5_and_9_cse = return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1
      & (fsm_output[17]);
  assign return_add_generic_AC_RND_CONV_false_5_or_4_cse = return_add_generic_AC_RND_CONV_false_20_ls_or_cse
      | return_add_generic_AC_RND_CONV_false_5_and_7_cse | return_add_generic_AC_RND_CONV_false_5_and_9_cse
      | (return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1 & (fsm_output[29]));
  assign return_add_generic_AC_RND_CONV_false_5_and_6_cse = (~ return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1)
      & (fsm_output[15]);
  assign return_add_generic_AC_RND_CONV_false_5_and_8_cse = (~ return_add_generic_AC_RND_CONV_false_10_acc_3_itm_11_1)
      & (fsm_output[17]);
  assign return_add_generic_AC_RND_CONV_false_5_and_10_cse = (~ return_add_generic_AC_RND_CONV_false_21_acc_3_itm_11_1)
      & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_3_or_14_cse = and_1014_cse | ((~ or_446_cse)
      & (fsm_output[8]));
  assign return_add_generic_AC_RND_CONV_false_3_or_16_cse = and_1032_cse | ((~ or_445_cse)
      & (fsm_output[24]));
  assign return_add_generic_AC_RND_CONV_false_5_or_6_cse = return_add_generic_AC_RND_CONV_false_20_ls_or_cse
      | return_add_generic_AC_RND_CONV_false_5_and_7_cse | return_add_generic_AC_RND_CONV_false_5_and_9_cse;
  assign stage_PE_qif_qelse_mux_12_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_rsp_0_9,
      m_in_15_1_lpi_1_dfm_1_rsp_0_10, mode_lpi_1_dfm);
  assign stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_0 = stage_PE_qif_qelse_mux_12_nl
      & inverse_lpi_1_dfm_1;
  assign stage_PE_qif_qelse_mux_16_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_rsp_0_10,
      m_in_15_1_lpi_1_dfm_1_rsp_0_11, mode_lpi_1_dfm);
  assign stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_1 = stage_PE_qif_qelse_mux_16_nl
      & inverse_lpi_1_dfm_1;
  assign stage_PE_qif_qelse_mux_1_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_rsp_0_12,
      m_in_15_1_lpi_1_dfm_1_rsp_0_13, mode_lpi_1_dfm);
  assign stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_3 = stage_PE_qif_qelse_mux_1_nl
      & inverse_lpi_1_dfm_1;
  assign stage_PE_qif_qelse_mux_17_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_rsp_0_11,
      m_in_15_1_lpi_1_dfm_1_rsp_0_12, mode_lpi_1_dfm);
  assign stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_2 = stage_PE_qif_qelse_mux_17_nl
      & inverse_lpi_1_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_11_and_45_cse = (~ return_add_generic_AC_RND_CONV_false_13_do_sub_sva)
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_11_and_46_cse = return_add_generic_AC_RND_CONV_false_13_do_sub_sva
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_1_and_itm = (~ return_add_generic_AC_RND_CONV_false_2_acc_3_itm_11_1)
      & or_1531_cse;
  assign return_add_generic_AC_RND_CONV_false_1_and_1_itm = return_add_generic_AC_RND_CONV_false_2_acc_3_itm_11_1
      & or_1531_cse;
  assign return_add_generic_AC_RND_CONV_false_1_and_2_itm = (~ return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1)
      & (fsm_output[8]);
  assign return_add_generic_AC_RND_CONV_false_1_and_3_itm = return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1
      & (fsm_output[8]);
  assign return_add_generic_AC_RND_CONV_false_5_or_1_itm = (fsm_output[15]) | (fsm_output[17])
      | (fsm_output[29]);
  assign or_1746_nl = (fsm_output[9]) | (fsm_output[23]) | (fsm_output[13]) | (fsm_output[12]);
  assign mux_nl = MUX_s_1_2_2((fsm_output[9]), or_1746_nl, BUTTERFLY_1_else_1_if_nor_cse);
  assign and_2619_nl = mode_lpi_1_dfm & mux_nl;
  assign or_1743_nl = and_2638_cse | (fsm_output[23]) | (fsm_output[13]) | (fsm_output[12]);
  assign mux_19_nl = MUX_s_1_2_2(and_2619_nl, or_1743_nl, fsm_output[15]);
  assign and_2620_ssc = (mux_19_nl | (fsm_output[29]) | (fsm_output[30]) | (fsm_output[6])
      | (fsm_output[28]) | (fsm_output[24]) | (fsm_output[22]) | (fsm_output[25]))
      & run_wen;
  assign BUTTERFLY_else_1_if_and_5_cse = or_tmp_773 & BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c7;
  assign return_add_generic_AC_RND_CONV_false_9_conc_59_itm_5_1 = MUX_v_5_2_2((reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[4:0]),
      (leading_sign_57_0_1_0_2_out_3[5:1]), return_add_generic_AC_RND_CONV_false_22_acc_3_itm_11_1);
  assign BUTTERFLY_1_nor_1_cse = ~(or_tmp_1003 | (fsm_output[8]));
  assign return_mult_generic_AC_RND_CONV_false_1_else_1_and_1_cse = (z_out_26[105])
      & (~ (fsm_output[36]));
  assign return_mult_generic_AC_RND_CONV_false_1_else_1_return_mult_generic_AC_RND_CONV_false_1_else_1_mux_2_cse
      = MUX_s_1_2_2((z_out_26[104]), return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp,
      fsm_output[36]);
  assign return_add_generic_AC_RND_CONV_false_1_and_54_cse = (~ return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11)
      & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_1_and_55_cse = return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11
      & (fsm_output[30]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      out1_rsci_idat_63 <= 1'b0;
      out1_rsci_idat_62_52 <= 11'b00000000000;
      out1_rsci_idat_51 <= 1'b0;
      out1_rsci_idat_50_0 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      out1_rsci_idat_63 <= 1'b0;
      out1_rsci_idat_62_52 <= 11'b00000000000;
      out1_rsci_idat_51 <= 1'b0;
      out1_rsci_idat_50_0 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( for_1_if_and_ssc ) begin
      out1_rsci_idat_63 <= MUX_s_1_2_2((out_f_d_rsci_q_d[63]), (in_f_d_rsci_q_d[63]),
          out1_rsci_idat_63_0_mx0c2);
      out1_rsci_idat_62_52 <= MUX1HOT_v_11_3_2((out_f_d_rsci_q_d[62:52]), return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_or_nl,
          (in_f_d_rsci_q_d[62:52]), {or_tmp_26 , out1_rsci_idat_63_0_mx0c1 , out1_rsci_idat_63_0_mx0c2});
      out1_rsci_idat_51 <= MUX1HOT_s_1_4_2((out_f_d_rsci_q_d[51]), (z_out[51]), return_mult_generic_AC_RND_CONV_false_6_op1_nan_sva_1,
          (in_f_d_rsci_q_d[51]), {or_tmp_26 , BUTTERFLY_if_1_and_nl , BUTTERFLY_if_1_and_1_nl
          , out1_rsci_idat_63_0_mx0c2});
      out1_rsci_idat_50_0 <= MUX1HOT_v_51_3_2((out_f_d_rsci_q_d[50:0]), return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_and_1_nl,
          (in_f_d_rsci_q_d[50:0]), {or_tmp_26 , out1_rsci_idat_63_0_mx0c1 , out1_rsci_idat_63_0_mx0c2});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      out1_rsci_idat_79_64 <= 16'b0000000000000000;
    end
    else if ( rst ) begin
      out1_rsci_idat_79_64 <= 16'b0000000000000000;
    end
    else if ( run_wen & (or_tmp_26 | out1_rsci_idat_79_64_mx0c1 | and_392_cse) )
        begin
      out1_rsci_idat_79_64 <= MUX1HOT_v_16_3_2(out_u_rsci_q_d, in_u_rsci_q_d, ({{1{stage_monty_mul_acc_2_psp_sva_1[14]}},
          stage_monty_mul_acc_2_psp_sva_1}), {or_tmp_26 , out1_rsci_idat_79_64_mx0c1
          , and_392_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_cgo_cse <= 1'b0;
      BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo <= 1'b0;
      BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo <= 1'b0;
      BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo <= 1'b0;
      BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo <= 1'b0;
      reg_out_u_triosy_obj_iswt0_cse <= 1'b0;
      reg_out1_rsci_iswt0_cse <= 1'b0;
      reg_out_u_rsci_cgo_ir_cse <= 1'b0;
      reg_out_f_d_rsci_cgo_ir_cse <= 1'b0;
      reg_in_u_rsci_cgo_ir_cse <= 1'b0;
      reg_in_f_d_rsci_cgo_ir_cse <= 1'b0;
      reg_ap_start_rsci_iswt0_cse <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_1_ftd <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_1_ftd_4 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_1_ftd_3 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_1_ftd_1 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_2 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_3 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_4 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_5 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_5 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_4 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_3 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_2 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_1 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_0 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_7 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_a_reg <= 9'b000000000;
      reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_addr_cse <= 10'b0000000000;
      return_add_generic_AC_RND_CONV_false_17_mux_7_itm_55_51 <= 5'b00000;
      return_add_generic_AC_RND_CONV_false_18_mux_1_itm_55_51 <= 5'b00000;
      return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva <= 1'b0;
      return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm <= 51'b000000000000000000000000000000000000000000000000000;
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_51 <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_0 <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_1 <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2 <= 4'b0000;
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_0 <= 4'b0000;
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_1 <= 2'b00;
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_2 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_cgo_cse <= 1'b0;
      BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo <= 1'b0;
      BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo <= 1'b0;
      BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo <= 1'b0;
      BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo <= 1'b0;
      reg_out_u_triosy_obj_iswt0_cse <= 1'b0;
      reg_out1_rsci_iswt0_cse <= 1'b0;
      reg_out_u_rsci_cgo_ir_cse <= 1'b0;
      reg_out_f_d_rsci_cgo_ir_cse <= 1'b0;
      reg_in_u_rsci_cgo_ir_cse <= 1'b0;
      reg_in_f_d_rsci_cgo_ir_cse <= 1'b0;
      reg_ap_start_rsci_iswt0_cse <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_1_ftd <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_1_ftd_4 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_1_ftd_3 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_1_ftd_1 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_2 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_3 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_4 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_5 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_5 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_4 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_3 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_2 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_1 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_0 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_b_ftd_7 <= 1'b0;
      reg_BUTTERFLY_i_div_cmp_a_reg <= 9'b000000000;
      reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_addr_cse <= 10'b0000000000;
      return_add_generic_AC_RND_CONV_false_17_mux_7_itm_55_51 <= 5'b00000;
      return_add_generic_AC_RND_CONV_false_18_mux_1_itm_55_51 <= 5'b00000;
      return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva <= 1'b0;
      return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm <= 51'b000000000000000000000000000000000000000000000000000;
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_51 <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_0 <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_1 <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2 <= 4'b0000;
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_0 <= 4'b0000;
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_1 <= 2'b00;
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_2 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen ) begin
      reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_cgo_cse <= or_dcpl_83 |
          or_dcpl_82;
      BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo <= inverse_lpi_1_dfm_1 & or_dcpl_85;
      BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo <= (~ inverse_lpi_1_dfm_1) &
          or_dcpl_85;
      BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo <= inverse_lpi_1_dfm_1 & or_dcpl_86;
      BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo <= (~ inverse_lpi_1_dfm_1)
          & or_dcpl_86;
      reg_out_u_triosy_obj_iswt0_cse <= (z_out_55[10]) & (fsm_output[37]);
      reg_out1_rsci_iswt0_cse <= fsm_output[36];
      reg_out_u_rsci_cgo_ir_cse <= or_670_rmff;
      reg_out_f_d_rsci_cgo_ir_cse <= or_671_rmff;
      reg_in_u_rsci_cgo_ir_cse <= or_672_rmff;
      reg_in_f_d_rsci_cgo_ir_cse <= or_673_rmff;
      reg_ap_start_rsci_iswt0_cse <= ~ and_dcpl_110;
      reg_BUTTERFLY_i_div_cmp_b_ftd <= MUX_s_1_2_2(stage_PE_index_const_mux_nl, stage_PE_index_const_mux_3_nl,
          or_tmp_46);
      reg_BUTTERFLY_i_div_cmp_b_1_ftd <= MUX_s_1_2_2(stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_3,
          stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_0_rsp_0, BUTTERFLY_i_or_3_cse);
      reg_BUTTERFLY_i_div_cmp_b_1_ftd_4 <= MUX_s_1_2_2(stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_2,
          stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_0_rsp_1, BUTTERFLY_i_or_3_cse);
      reg_BUTTERFLY_i_div_cmp_b_1_ftd_3 <= MUX_s_1_2_2(stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_1,
          stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_1, BUTTERFLY_i_or_3_cse);
      reg_BUTTERFLY_i_div_cmp_b_1_ftd_1 <= MUX_s_1_2_2(stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_0,
          stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_1, BUTTERFLY_i_or_3_cse);
      reg_BUTTERFLY_i_div_cmp_b_ftd_2 <= MUX_s_1_2_2(stage_PE_index_const_mux_2_nl,
          stage_PE_index_const_mux_7_nl, or_tmp_46);
      reg_BUTTERFLY_i_div_cmp_b_ftd_3 <= MUX_s_1_2_2(stage_PE_mux1h_nl, stage_PE_mux1h_7_nl,
          or_tmp_46);
      reg_BUTTERFLY_i_div_cmp_b_ftd_4 <= MUX_s_1_2_2(stage_PE_mux1h_1_nl, stage_PE_mux1h_9_nl,
          or_tmp_46);
      reg_BUTTERFLY_i_div_cmp_b_ftd_5 <= MUX_s_1_2_2(stage_PE_mux1h_2_nl, stage_PE_mux1h_11_nl,
          or_tmp_46);
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_5 <= MUX1HOT_s_1_3_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_5,
          t_in_10_0_lpi_1_dfm_1_7, stage_PE_1_index_const_9_1_lpi_2_dfm_5, {BUTTERFLY_i_or_4_ssc
          , BUTTERFLY_i_or_5_ssc , BUTTERFLY_i_or_3_cse});
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_4 <= MUX1HOT_s_1_3_2(stage_PE_qif_qelse_mux_15_itm,
          t_in_10_0_lpi_1_dfm_1_6, stage_PE_1_index_const_9_1_lpi_2_dfm_4, {BUTTERFLY_i_or_4_ssc
          , BUTTERFLY_i_or_5_ssc , BUTTERFLY_i_or_3_cse});
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_3 <= MUX1HOT_s_1_3_2(t_in_10_0_lpi_1_dfm_1_6,
          t_in_10_0_lpi_1_dfm_1_5, stage_PE_1_index_const_9_1_lpi_2_dfm_3, {BUTTERFLY_i_and_14_nl
          , BUTTERFLY_i_or_7_nl , BUTTERFLY_i_or_3_cse});
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_2 <= MUX1HOT_s_1_3_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_2,
          t_in_10_0_lpi_1_dfm_1_4, stage_PE_1_index_const_9_1_lpi_2_dfm_2, {BUTTERFLY_i_or_4_ssc
          , BUTTERFLY_i_or_5_ssc , BUTTERFLY_i_or_3_cse});
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_1 <= MUX1HOT_s_1_3_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_1,
          t_in_10_0_lpi_1_dfm_1_3, stage_PE_1_index_const_9_1_lpi_2_dfm_1, {BUTTERFLY_i_or_4_ssc
          , BUTTERFLY_i_or_5_ssc , BUTTERFLY_i_or_3_cse});
      reg_BUTTERFLY_i_div_cmp_b_ftd_6_0 <= MUX1HOT_s_1_3_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_0,
          t_in_10_0_lpi_1_dfm_1_2, stage_PE_1_index_const_9_1_lpi_2_dfm_0, {BUTTERFLY_i_or_4_ssc
          , BUTTERFLY_i_or_5_ssc , BUTTERFLY_i_or_3_cse});
      reg_BUTTERFLY_i_div_cmp_b_ftd_7 <= MUX_s_1_2_2(stage_PE_mux1h_3_nl, stage_PE_mux1h_13_nl,
          or_tmp_46);
      reg_BUTTERFLY_i_div_cmp_a_reg <= MUX_v_9_2_2(9'b000000000, BUTTERFLY_i_mux_1_nl,
          t_in_not_nl);
      reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_addr_cse <= nl_reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_addr_cse[9:0];
      return_add_generic_AC_RND_CONV_false_17_mux_7_itm_55_51 <= MUX_v_5_2_2((z_out_34[56:52]),
          (~ (z_out_34[56:52])), return_add_generic_AC_RND_CONV_false_17_or_nl);
      return_add_generic_AC_RND_CONV_false_18_mux_1_itm_55_51 <= MUX1HOT_v_5_4_2((z_out_34[56:52]),
          (~ (z_out_34[56:52])), (~ (return_add_generic_AC_RND_CONV_false_25_rshift_itm[56:52])),
          (return_add_generic_AC_RND_CONV_false_25_rshift_itm[56:52]), {return_add_generic_AC_RND_CONV_false_18_return_add_generic_AC_RND_CONV_false_18_nor_nl
          , return_add_generic_AC_RND_CONV_false_18_and_2_nl , return_add_generic_AC_RND_CONV_false_18_and_3_nl
          , return_add_generic_AC_RND_CONV_false_18_and_4_cse});
      return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva <= MUX1HOT_s_1_10_2(all_same_out,
          return_mult_generic_AC_RND_CONV_false_1_if_3_return_mult_generic_AC_RND_CONV_false_1_if_3_or_1_nl,
          leading_sign_57_0_1_0_6_out_2, return_mult_generic_AC_RND_CONV_false_2_if_3_return_mult_generic_AC_RND_CONV_false_2_if_3_or_1_nl,
          all_same_out_1, leading_sign_57_0_1_0_10_out_2, leading_sign_57_0_1_0_17_out_2,
          leading_sign_57_0_1_0_19_out_2, return_mult_generic_AC_RND_CONV_false_5_if_3_return_mult_generic_AC_RND_CONV_false_5_if_3_or_1_nl,
          leading_sign_57_0_1_0_20_out_2, {(fsm_output[7]) , (fsm_output[9]) , (fsm_output[10])
          , (fsm_output[11]) , return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse
          , (fsm_output[14]) , (fsm_output[23]) , (fsm_output[26]) , (fsm_output[27])
          , (fsm_output[28])});
      return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva <= MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp,
          (({stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_1 , stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0})
          == ({operator_6_false_18_acc_psp_sva_10_0_rsp_0 , operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0
          , operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1})), return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1,
          ((stage_PE_1_x_im_d_sva[62:52]) == ({return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_mx0w2
          , return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1})), return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1,
          return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp,
          (({stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx1_10_1 , stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx1_0})
          == ({operator_6_false_18_acc_psp_sva_10_0_rsp_0 , operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0
          , operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1})), return_add_generic_AC_RND_CONV_false_19_acc_2_itm_11_1,
          {(fsm_output[7]) , (fsm_output[9]) , (fsm_output[10]) , (fsm_output[13])
          , (fsm_output[15]) , (fsm_output[23]) , (fsm_output[25]) , (fsm_output[26])});
      return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm <= MUX1HOT_v_51_4_2(return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1,
          stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0, return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0,
          stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1, {(fsm_output[8]) , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_18_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_5_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_24_cse});
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_51 <= MUX_s_1_2_2(stage_PE_tmp_re_d_1_lpi_3_dfm_51_mx0,
          stage_PE_1_tmp_re_d_1_lpi_3_dfm_51_mx1, fsm_output[25]);
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_0 <= MUX1HOT_s_1_8_2((return_add_generic_AC_RND_CONV_false_4_e_dif_sat_or_cse[5]),
          (leading_sign_57_0_1_0_4_out_3[5]), (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_3_itm[5]),
          (rtn_out_1[5]), (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_5_itm[5]),
          (leading_sign_57_0_1_0_10_out_3[5]), (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_9_itm[5]),
          (leading_sign_57_0_1_0_21_out_3[5]), {(fsm_output[6]) , (fsm_output[7])
          , (fsm_output[10]) , return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse
          , (fsm_output[13]) , (fsm_output[14]) , (fsm_output[26]) , (fsm_output[28])});
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_1 <= MUX1HOT_s_1_9_2((return_add_generic_AC_RND_CONV_false_4_e_dif_sat_or_cse[4]),
          (leading_sign_57_0_1_0_4_out_3[4]), (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_3_itm[4]),
          (rtn_out_1[4]), (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_5_itm[4]),
          (leading_sign_57_0_1_0_10_out_3[4]), (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_conc_4_itm_4_1[3]),
          (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_9_itm[4]), (leading_sign_57_0_1_0_21_out_3[4]),
          {(fsm_output[6]) , (fsm_output[7]) , (fsm_output[10]) , return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse
          , (fsm_output[13]) , (fsm_output[14]) , (fsm_output[15]) , (fsm_output[26])
          , (fsm_output[28])});
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2 <= MUX1HOT_v_4_10_2((return_add_generic_AC_RND_CONV_false_4_e_dif_sat_or_cse[3:0]),
          (leading_sign_57_0_1_0_4_out_3[3:0]), return_mult_generic_AC_RND_CONV_false_1_if_nand_1_nl,
          (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_3_itm[3:0]), (rtn_out_1[3:0]),
          (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_5_itm[3:0]), (leading_sign_57_0_1_0_10_out_3[3:0]),
          ({(return_add_generic_AC_RND_CONV_false_10_e_dif_sat_conc_4_itm_4_1[2:0])
          , return_add_generic_AC_RND_CONV_false_11_mux_23_nl}), (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_mux1h_9_itm[3:0]),
          (leading_sign_57_0_1_0_21_out_3[3:0]), {(fsm_output[6]) , (fsm_output[7])
          , (fsm_output[8]) , (fsm_output[10]) , return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse
          , (fsm_output[13]) , (fsm_output[14]) , (fsm_output[15]) , (fsm_output[26])
          , (fsm_output[28])});
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_0 <= MUX1HOT_v_4_5_2((z_out_7[56:53]),
          (return_add_generic_AC_RND_CONV_false_4_res_mant_4_sva_1[56:53]), (z_out_8[56:53]),
          (return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_2[56:53]), (return_add_generic_AC_RND_CONV_false_21_res_mant_4_sva_1[56:53]),
          {return_add_generic_AC_RND_CONV_false_10_res_mant_or_9_cse , (fsm_output[7])
          , return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse , (fsm_output[14])
          , (fsm_output[28])});
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_1 <= MUX1HOT_v_2_6_2((z_out_7[52:51]),
          (return_add_generic_AC_RND_CONV_false_4_res_mant_4_sva_1[52:51]), (z_out_53[52:51]),
          (z_out_8[52:51]), (return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_2[52:51]),
          (return_add_generic_AC_RND_CONV_false_21_res_mant_4_sva_1[52:51]), {return_add_generic_AC_RND_CONV_false_10_res_mant_or_9_cse
          , (fsm_output[7]) , or_1143_itm , return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse
          , (fsm_output[14]) , (fsm_output[28])});
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_rsp_2 <= MUX1HOT_v_51_7_2((z_out_7[50:0]),
          (return_add_generic_AC_RND_CONV_false_4_res_mant_4_sva_1[50:0]), (z_out_53[50:0]),
          (z_out_8[50:0]), (return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva_2[50:0]),
          (return_add_generic_AC_RND_CONV_false_17_res_rounded_lpi_3_dfm_51_0_1[50:0]),
          (return_add_generic_AC_RND_CONV_false_21_res_mant_4_sva_1[50:0]), {return_add_generic_AC_RND_CONV_false_10_res_mant_or_9_cse
          , (fsm_output[7]) , or_1143_itm , return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse
          , (fsm_output[14]) , (fsm_output[23]) , (fsm_output[28])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[11])) | (~ mode_lpi_1_dfm) | (return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp[12])))
        ) begin
      return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_2_if_acc_1_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & mode_lpi_1_dfm & (~ (stage_u_add_3_acc_itm_rsp_1[12])) &
        (fsm_output[9]) ) begin
      return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_1_if_acc_1_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[7])) | and_565_cse)) ) begin
      return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[7])) | and_569_cse)) ) begin
      return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[10])) | and_573_cse)) ) begin
      return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_3_if_acc_2_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[9])) | or_dcpl_164 | or_dcpl_172 | or_dcpl_151))
        ) begin
      return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[9])) | return_add_generic_AC_RND_CONV_false_1_r_inf_lpi_3_dfm_2
        | or_dcpl_172 | or_dcpl_152)) ) begin
      return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & and_dcpl_121 & and_dcpl_118 & (~ operator_11_true_return_13_sva)
        & mode_lpi_1_dfm & (fsm_output[11]) ) begin
      return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (fsm_output[10]) & return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1
        & mode_lpi_1_dfm ) begin
      return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp <= ~((operator_33_true_12_acc_tmp[11:0]==12'b011111111111));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[13])) | or_dcpl_193 | and_dcpl_125 | or_dcpl_190))
        ) begin
      return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[13])) | or_dcpl_201 | and_dcpl_127 | or_dcpl_198))
        ) begin
      return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[27])) | (return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp[12])
        | (~ mode_lpi_1_dfm))) ) begin
      return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_5_if_acc_1_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[24])) | (z_out_45[12]) | (~ mode_lpi_1_dfm)))
        ) begin
      return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_4_if_acc_1_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[23])) | and_565_cse)) ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[23])) | and_569_cse)) ) begin
      return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[26])) | and_573_cse)) ) begin
      return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_3_if_acc_2_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[25])) | and_565_cse)) ) begin
      return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[25])) | and_569_cse)) ) begin
      return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (fsm_output[26]) & return_add_generic_AC_RND_CONV_false_19_acc_2_itm_11_1
        & mode_lpi_1_dfm ) begin
      return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp <= ~((z_out_16[11:0]==12'b011111111111));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[27])) | or_dcpl_212 | and_dcpl_129 | operator_11_true_return_15_sva
        | or_dcpl_190)) ) begin
      return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[29])) | or_dcpl_193 | and_dcpl_131 | or_dcpl_190))
        ) begin
      return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[29])) | or_dcpl_201 | and_dcpl_132 | or_dcpl_198))
        ) begin
      return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[36])) | or_dcpl_75 | (operator_16_false_io_read_mode1_rsc_cse_sva[13:4]!=10'b0000000000)
        | or_dcpl_65 | or_dcpl_64 | operator_16_false_operator_16_false_nor_cse_sva
        | (z_out_51[11]))) ) begin
      return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[14])) | and_631_cse)) ) begin
      return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[15])) | or_dcpl_238 | (~ return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1)))
        ) begin
      return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp <= ~((z_out_48[11:0]==12'b011111111111));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[15])) | return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2
        | or_dcpl_250 | and_dcpl_135 | or_dcpl_238)) ) begin
      return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[16])) | or_dcpl_172 | operator_11_true_return_17_sva
        | return_add_generic_AC_RND_CONV_false_11_r_inf_lpi_3_dfm_2 | and_dcpl_136
        | return_add_generic_AC_RND_CONV_false_15_do_sub_sva | or_dcpl_238)) ) begin
      return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[17])) | or_dcpl_25 | operator_11_true_return_15_sva
        | return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2 | and_dcpl_135
        | operator_11_true_return_13_sva | or_dcpl_238)) ) begin
      return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[30])) | return_add_generic_AC_RND_CONV_false_24_r_inf_lpi_3_dfm_2
        | or_dcpl_172 | and_dcpl_139 | or_dcpl_238)) ) begin
      return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[30])) | return_add_generic_AC_RND_CONV_false_25_r_inf_lpi_3_dfm_2
        | or_dcpl_250 | and_dcpl_141 | or_dcpl_238)) ) begin
      return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[30])) | and_631_cse)) ) begin
      return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[30])) | return_add_generic_AC_RND_CONV_false_23_r_inf_lpi_3_dfm_2
        | or_dcpl_250 | and_dcpl_143 | or_dcpl_238)) ) begin
      return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_16_false_io_read_mode1_rsc_cse_sva <= 16'b0000000000000000;
    end
    else if ( rst ) begin
      operator_16_false_io_read_mode1_rsc_cse_sva <= 16'b0000000000000000;
    end
    else if ( operator_16_false_and_cse & (~ operator_16_false_operator_16_false_nor_tmp)
        ) begin
      operator_16_false_io_read_mode1_rsc_cse_sva <= mode1_rsci_idat;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_16_false_operator_16_false_nor_cse_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_16_false_operator_16_false_nor_cse_sva <= 1'b0;
    end
    else if ( operator_16_false_and_cse ) begin
      operator_16_false_operator_16_false_nor_cse_sva <= operator_16_false_operator_16_false_nor_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      t_in_10_0_lpi_1_dfm_1_8 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_7 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_6 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_5 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_4 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_3 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_2 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_1 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_0 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_10 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_9 <= 1'b0;
      for_i_3_0_sva <= 4'b0000;
      m_in_15_1_lpi_1_dfm_1_rsp_0_9 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_rsp_0_10 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_rsp_0_11 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_rsp_0_13 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_rsp_0_12 <= 1'b0;
    end
    else if ( rst ) begin
      t_in_10_0_lpi_1_dfm_1_8 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_7 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_6 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_5 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_4 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_3 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_2 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_1 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_0 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_10 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_9 <= 1'b0;
      for_i_3_0_sva <= 4'b0000;
      m_in_15_1_lpi_1_dfm_1_rsp_0_9 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_rsp_0_10 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_rsp_0_11 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_rsp_0_13 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_rsp_0_12 <= 1'b0;
    end
    else if ( t_in_and_cse ) begin
      t_in_10_0_lpi_1_dfm_1_8 <= t_in_10_0_lpi_1_dfm_1_9 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_7 <= t_in_10_0_lpi_1_dfm_1_8 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_6 <= t_in_10_0_lpi_1_dfm_1_7 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_5 <= t_in_10_0_lpi_1_dfm_1_6 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_4 <= t_in_10_0_lpi_1_dfm_1_5 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_3 <= t_in_10_0_lpi_1_dfm_1_4 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_2 <= t_in_10_0_lpi_1_dfm_1_3 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_1 <= t_in_10_0_lpi_1_dfm_1_2 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_0 <= t_in_10_0_lpi_1_dfm_1_1 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_10 <= (~(operator_16_false_1_operator_16_false_1_and_mdf_sva_1
          | operator_16_false_operator_16_false_nor_tmp)) & nor_155_cse;
      t_in_10_0_lpi_1_dfm_1_9 <= MUX_s_1_2_2(mode_lpi_1_dfm_mx0w0, t_in_10_0_lpi_1_dfm_1_10,
          mode_or_cse);
      for_i_3_0_sva <= MUX_v_4_2_2(4'b0000, (z_out_13[3:0]), not_681_nl);
      m_in_15_1_lpi_1_dfm_1_rsp_0_9 <= t_in_10_0_lpi_1_dfm_1_0 & (~ (fsm_output[1]));
      m_in_15_1_lpi_1_dfm_1_rsp_0_10 <= m_in_15_1_lpi_1_dfm_1_rsp_0_9 & (~ (fsm_output[1]));
      m_in_15_1_lpi_1_dfm_1_rsp_0_11 <= m_in_15_1_lpi_1_dfm_1_rsp_0_10 & (~ (fsm_output[1]));
      m_in_15_1_lpi_1_dfm_1_rsp_0_13 <= m_in_15_1_lpi_1_dfm_1_rsp_0_12 & (~ (fsm_output[1]));
      m_in_15_1_lpi_1_dfm_1_rsp_0_12 <= m_in_15_1_lpi_1_dfm_1_rsp_0_11 & (~ (fsm_output[1]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      mode_lpi_1_dfm <= 1'b0;
      inverse_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( rst ) begin
      mode_lpi_1_dfm <= 1'b0;
      inverse_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( mode_and_cse ) begin
      mode_lpi_1_dfm <= mode_lpi_1_dfm_mx0w0;
      inverse_lpi_1_dfm_1 <= ~(((mode1_rsci_idat==16'b0000000000000010)) | operator_16_false_operator_16_false_nor_tmp);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_qr_1_10_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_qr_1_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_qr_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_index_const_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_15_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_10_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_1 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_1 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_0_rsp_0 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_0_rsp_1 <= 1'b0;
    end
    else if ( rst ) begin
      stage_PE_1_qr_1_10_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_qr_1_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_qr_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_index_const_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_15_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_10_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_1 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_1 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_0_rsp_0 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_0_rsp_1 <= 1'b0;
    end
    else if ( stage_PE_1_and_2_cse ) begin
      stage_PE_1_qr_1_10_1_lpi_2_dfm_8 <= MUX1HOT_s_1_3_2(t_in_10_0_lpi_1_dfm_1_1,
          t_in_10_0_lpi_1_dfm_1_9, t_in_10_0_lpi_1_dfm_1_8, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_7 <= MUX1HOT_s_1_3_2(t_in_10_0_lpi_1_dfm_1_2,
          t_in_10_0_lpi_1_dfm_1_8, t_in_10_0_lpi_1_dfm_1_7, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_6 <= MUX1HOT_s_1_3_2(t_in_10_0_lpi_1_dfm_1_3,
          t_in_10_0_lpi_1_dfm_1_7, t_in_10_0_lpi_1_dfm_1_6, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_5 <= MUX1HOT_s_1_3_2(t_in_10_0_lpi_1_dfm_1_4,
          t_in_10_0_lpi_1_dfm_1_6, t_in_10_0_lpi_1_dfm_1_5, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_4 <= MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_5, t_in_10_0_lpi_1_dfm_1_4,
          stage_PE_1_and_1_tmp);
      stage_PE_1_qr_1_10_1_lpi_2_dfm_3 <= MUX1HOT_s_1_3_2(t_in_10_0_lpi_1_dfm_1_6,
          t_in_10_0_lpi_1_dfm_1_4, t_in_10_0_lpi_1_dfm_1_3, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_2 <= MUX1HOT_s_1_3_2(t_in_10_0_lpi_1_dfm_1_7,
          t_in_10_0_lpi_1_dfm_1_3, t_in_10_0_lpi_1_dfm_1_2, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_1 <= MUX1HOT_s_1_3_2(t_in_10_0_lpi_1_dfm_1_8,
          t_in_10_0_lpi_1_dfm_1_2, t_in_10_0_lpi_1_dfm_1_1, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_0 <= MUX1HOT_s_1_3_2(t_in_10_0_lpi_1_dfm_1_9,
          t_in_10_0_lpi_1_dfm_1_1, t_in_10_0_lpi_1_dfm_1_0, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_0_lpi_2_dfm <= t_in_10_0_lpi_1_dfm_1_10;
      stage_PE_1_qr_10_1_lpi_2_dfm_8 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_8,
          t_in_10_0_lpi_1_dfm_1_9, or_tmp_181);
      stage_PE_1_qr_10_1_lpi_2_dfm_7 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_7,
          t_in_10_0_lpi_1_dfm_1_8, or_tmp_181);
      stage_PE_1_qr_10_1_lpi_2_dfm_6 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_6,
          t_in_10_0_lpi_1_dfm_1_7, or_tmp_181);
      stage_PE_1_qr_10_1_lpi_2_dfm_5 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_5,
          t_in_10_0_lpi_1_dfm_1_6, or_tmp_181);
      stage_PE_1_qr_10_1_lpi_2_dfm_4 <= MUX_s_1_2_2(stage_PE_qif_qelse_mux_18_nl,
          t_in_10_0_lpi_1_dfm_1_5, or_tmp_181);
      stage_PE_1_qr_10_1_lpi_2_dfm_3 <= MUX_s_1_2_2(stage_PE_qif_qelse_mux_5_nl,
          t_in_10_0_lpi_1_dfm_1_4, or_tmp_181);
      stage_PE_1_qr_10_1_lpi_2_dfm_2 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_2,
          t_in_10_0_lpi_1_dfm_1_3, or_tmp_181);
      stage_PE_1_qr_10_1_lpi_2_dfm_1 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_1,
          t_in_10_0_lpi_1_dfm_1_2, or_tmp_181);
      stage_PE_1_qr_10_1_lpi_2_dfm_0 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_0,
          t_in_10_0_lpi_1_dfm_1_1, or_tmp_181);
      stage_PE_1_qr_0_lpi_2_dfm <= MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_9, t_in_10_0_lpi_1_dfm_1_10,
          stage_PE_qif_qelse_or_nl);
      stage_PE_1_index_const_9_1_lpi_2_dfm_8 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_8,
          t_in_10_0_lpi_1_dfm_1_10, or_tmp_181);
      stage_PE_1_index_const_9_1_lpi_2_dfm_7 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_7,
          t_in_10_0_lpi_1_dfm_1_9, or_tmp_181);
      stage_PE_1_index_const_9_1_lpi_2_dfm_6 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_6,
          t_in_10_0_lpi_1_dfm_1_8, or_tmp_181);
      stage_PE_1_index_const_9_1_lpi_2_dfm_5 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_5,
          t_in_10_0_lpi_1_dfm_1_7, or_tmp_181);
      stage_PE_1_index_const_9_1_lpi_2_dfm_4 <= MUX_s_1_2_2(stage_PE_qif_qelse_mux_15_itm,
          t_in_10_0_lpi_1_dfm_1_6, or_tmp_181);
      stage_PE_1_index_const_9_1_lpi_2_dfm_3 <= MUX_s_1_2_2(stage_PE_qif_qelse_mux_19_nl,
          t_in_10_0_lpi_1_dfm_1_5, or_tmp_181);
      stage_PE_1_index_const_9_1_lpi_2_dfm_2 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_2,
          t_in_10_0_lpi_1_dfm_1_4, or_tmp_181);
      stage_PE_1_index_const_9_1_lpi_2_dfm_1 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_1,
          t_in_10_0_lpi_1_dfm_1_3, or_tmp_181);
      stage_PE_1_index_const_9_1_lpi_2_dfm_0 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_0,
          t_in_10_0_lpi_1_dfm_1_2, or_tmp_181);
      stage_PE_1_index_const_0_lpi_2_dfm <= MUX_s_1_2_2(stage_PE_asn_13_mx0w0, t_in_10_0_lpi_1_dfm_1_1,
          or_tmp_181);
      stage_PE_1_index_const_15_lpi_2_dfm <= stage_PE_index_const_15_lpi_2_dfm_mx0w0;
      stage_PE_1_index_const_10_lpi_2_dfm <= stage_PE_index_const_10_lpi_2_dfm_mx0w0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_1 <= stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_1 <= stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_1;
      stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_0_rsp_0 <= stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_3;
      stage_PE_1_index_const_14_11_lpi_2_dfm_rsp_0_rsp_0_rsp_1 <= stage_PE_index_const_14_11_lpi_2_dfm_mx0w0_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_fry_9_0_sva <= 10'b0000000000;
    end
    else if ( rst ) begin
      BUTTERFLY_1_fry_9_0_sva <= 10'b0000000000;
    end
    else if ( run_wen & (~((~((fsm_output[33]) | (fsm_output[2]))) & and_dcpl_164
        & and_dcpl_110 & and_dcpl_179 & nor_90_cse & (~((fsm_output[32]) | (fsm_output[20])))
        & (~((fsm_output[18]) | (fsm_output[34]) | (fsm_output[16]))))) ) begin
      BUTTERFLY_1_fry_9_0_sva <= MUX_v_10_2_2(10'b0000000000, BUTTERFLY_fry_BUTTERFLY_fry_mux_nl,
          nor_155_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_26_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_26_sva <= 1'b0;
    end
    else if ( run_wen & ((~(inverse_lpi_1_dfm_1 | (and_dcpl_170 & (~ (fsm_output[38]))
        & and_dcpl_179 & nor_8_cse & (~((fsm_output[5]) | (fsm_output[21])))))) |
        (fsm_output[2])) ) begin
      operator_11_true_return_26_sva <= MUX1HOT_s_1_3_2(stage_PE_1_and_1_tmp, operator_11_true_return_3_sva_mx1w0,
          operator_11_true_return_26_sva_2, {(fsm_output[2]) , (fsm_output[5]) ,
          (fsm_output[21])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_6_false_49_acc_psp_sva_11_9 <= 3'b000;
    end
    else if ( rst ) begin
      operator_6_false_49_acc_psp_sva_11_9 <= 3'b000;
    end
    else if ( run_wen & mode_lpi_1_dfm ) begin
      operator_6_false_49_acc_psp_sva_11_9 <= operator_6_false_49_acc_sdt[11:9];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_6_false_49_acc_psp_sva_8_0 <= 9'b000000000;
    end
    else if ( rst ) begin
      operator_6_false_49_acc_psp_sva_8_0 <= 9'b000000000;
    end
    else if ( nor_88_cse & nor_87_cse & (~((fsm_output[5]) | (fsm_output[10]))) &
        (~((fsm_output[13:12]!=2'b00))) & nor_90_cse & nor_145_cse & (~((fsm_output[16])
        | (fsm_output[11]))) & (~((fsm_output[3]) | (fsm_output[7]))) & run_wen )
        begin
      operator_6_false_49_acc_psp_sva_8_0 <= MUX_v_9_2_2(BUTTERFLY_n_and_nl, (operator_6_false_49_acc_sdt[8:0]),
          fsm_output[28]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm <= 1'b0;
    end
    else if ( rst ) begin
      BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm <= 1'b0;
    end
    else if ( run_wen & (~((~((fsm_output[2]) | (fsm_output[3]) | (fsm_output[19])))
        & and_dcpl_150 & and_dcpl_147 & nor_8_cse)) & mode_lpi_1_dfm ) begin
      BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm <= (operator_6_false_49_acc_psp_sva_8_0==9'b011111111);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_BUTTERFLY_1_i_9_0_ftd <= 1'b0;
    end
    else if ( rst ) begin
      reg_BUTTERFLY_1_i_9_0_ftd <= 1'b0;
    end
    else if ( BUTTERFLY_1_i_and_ssc ) begin
      reg_BUTTERFLY_1_i_9_0_ftd <= BUTTERFLY_i_9_0_sva_1[9];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_BUTTERFLY_1_i_9_0_ftd_1 <= 9'b000000000;
    end
    else if ( rst ) begin
      reg_BUTTERFLY_1_i_9_0_ftd_1 <= 9'b000000000;
    end
    else if ( BUTTERFLY_1_i_and_ssc & (~ or_tmp_567) ) begin
      reg_BUTTERFLY_1_i_9_0_ftd_1 <= MUX_v_9_2_2((BUTTERFLY_i_9_0_sva_1[8:0]), (BUTTERFLY_1_fry_9_0_sva[8:0]),
          BUTTERFLY_i_or_2_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & (~(BUTTERFLY_if_1_or_3_cse | (fsm_output[27]) | or_dcpl_305
        | (fsm_output[13]) | or_dcpl_328 | or_dcpl_300)) ) begin
      return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm <= MUX1HOT_s_1_7_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1,
          return_extract_44_return_extract_44_or_1_tmp, stage_PE_1_tmp_re_d_1_lpi_3_dfm_51_mx1,
          return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_3_nl,
          return_add_generic_AC_RND_CONV_false_10_op1_mu_mux1h_3_cse, return_add_generic_AC_RND_CONV_false_25_r_nan_or_1_nl,
          (return_add_generic_AC_RND_CONV_false_25_res_rounded_lpi_3_dfm_51_0_1[51]),
          {(fsm_output[5]) , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_1_cse
          , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_2_cse , (fsm_output[26])
          , (fsm_output[29]) , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_3_nl
          , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_4_nl});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm <= 1'b0;
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_63 <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm <= 1'b0;
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_63 <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_14_op1_mu_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm <= MUX1HOT_s_1_11_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1,
          stage_PE_tmp_re_d_1_lpi_3_dfm_51_mx0, stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx1_50,
          (return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1[50]), return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2,
          return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm_1,
          stage_PE_1_tmp_re_d_1_lpi_3_dfm_51_mx1, stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx2_50,
          (return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1[50]), BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx3,
          {(fsm_output[5]) , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_5_cse
          , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_6_cse , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_7_cse
          , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_8_cse , (fsm_output[13])
          , (fsm_output[21]) , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_1_cse
          , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_2_cse , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_11_cse
          , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_12_cse});
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_63 <= MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_11_mux_19_cse,
          stage_d_mul_return_d_63_sva_1, stage_PE_1_tmp_re_d_1_lpi_3_dfm_63_mx1,
          stage_d_mul_return_d_1_63_sva_1, {(fsm_output[9]) , (fsm_output[10]) ,
          (fsm_output[25]) , (fsm_output[26])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_mux_7_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_mux_7_itm <= 1'b0;
    end
    else if ( run_wen & ((inverse_lpi_1_dfm_1 & (~(or_dcpl_354 | (fsm_output[10])
        | (fsm_output[7]) | (fsm_output[23]) | or_dcpl_300))) | (fsm_output[5]) |
        (fsm_output[13]) | (fsm_output[14]) | (fsm_output[21]) | (fsm_output[29]))
        ) begin
      return_add_generic_AC_RND_CONV_false_10_mux_7_itm <= MUX1HOT_s_1_15_2(return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp,
          return_add_generic_AC_RND_CONV_false_1_if_2_return_add_generic_AC_RND_CONV_false_1_if_2_and_2_nl,
          (stage_PE_1_x_im_d_sva[63]), (out_f_d_rsci_q_d[63]), return_add_generic_AC_RND_CONV_false_9_if_2_return_add_generic_AC_RND_CONV_false_9_if_2_and_2_nl,
          (stage_PE_1_x_re_d_sva[63]), return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_10_if_2_return_add_generic_AC_RND_CONV_false_10_if_2_and_1_mx3w0,
          operator_11_true_return_15_sva, return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp,
          return_add_generic_AC_RND_CONV_false_16_if_2_return_add_generic_AC_RND_CONV_false_16_if_2_nor_1_nl,
          (~ (in_f_d_rsci_q_d[63])), return_add_generic_AC_RND_CONV_false_13_if_2_return_add_generic_AC_RND_CONV_false_13_if_2_and_2_nl,
          (in_f_d_rsci_q_d[63]), (stage_PE_1_tmp_im_d_1_sva_1_63_51[12]), {(fsm_output[5])
          , return_add_generic_AC_RND_CONV_false_10_and_2_nl , return_add_generic_AC_RND_CONV_false_10_or_5_nl
          , return_add_generic_AC_RND_CONV_false_10_and_15_nl , return_add_generic_AC_RND_CONV_false_10_or_nl
          , return_add_generic_AC_RND_CONV_false_10_or_6_nl , return_add_generic_AC_RND_CONV_false_10_or_7_nl
          , return_add_generic_AC_RND_CONV_false_10_and_6_cse , return_add_generic_AC_RND_CONV_false_10_and_19_cse
          , (fsm_output[21]) , return_add_generic_AC_RND_CONV_false_10_and_8_nl ,
          return_add_generic_AC_RND_CONV_false_10_and_21_nl , return_add_generic_AC_RND_CONV_false_10_and_10_nl
          , return_add_generic_AC_RND_CONV_false_10_and_22_nl , return_add_generic_AC_RND_CONV_false_10_and_23_nl});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_17_m_zero_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_17_m_zero_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_352 | return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse))
        ) begin
      return_extract_17_m_zero_sva <= MUX1HOT_s_1_7_2(return_extract_3_m_zero_sva_1,
          return_extract_17_m_zero_return_extract_17_m_zero_nor_nl, return_extract_17_m_zero_sva_mx0w3,
          return_extract_15_m_zero_mux1h_3_cse, return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_svs_1,
          return_extract_47_m_zero_return_extract_47_m_zero_nor_nl, return_extract_59_m_zero_return_extract_59_m_zero_nor_nl,
          {(fsm_output[5]) , (fsm_output[8]) , or_916_nl , (fsm_output[21]) , (fsm_output[23])
          , (fsm_output[24]) , (fsm_output[29])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_44_m_zero_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_44_m_zero_sva <= 1'b0;
    end
    else if ( run_wen & ((inverse_lpi_1_dfm_1 & (~(or_dcpl_367 | (fsm_output[11])
        | or_dcpl_107 | or_dcpl_328 | or_dcpl_365))) | (fsm_output[5]) | (fsm_output[23])
        | (fsm_output[25]) | (fsm_output[26]) | (fsm_output[29])) ) begin
      return_extract_44_m_zero_sva <= MUX1HOT_s_1_5_2(return_extract_3_m_zero_sva_1,
          return_extract_45_m_zero_return_extract_45_m_zero_nor_nl, return_extract_44_m_zero_return_extract_44_m_zero_nor_nl,
          return_extract_52_m_zero_return_extract_52_m_zero_nor_nl, return_extract_57_m_zero_return_extract_57_m_zero_nor_nl,
          {return_extract_17_m_zero_or_1_nl , (fsm_output[23]) , (fsm_output[25])
          , (fsm_output[26]) , (fsm_output[29])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_1_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_367 | or_dcpl_305 | return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
        | (fsm_output[15]) | (fsm_output[8]))) ) begin
      operator_11_true_return_1_sva <= MUX1HOT_s_1_10_2(operator_11_true_return_3_sva_mx1w0,
          operator_11_true_12_operator_11_true_12_and_nl, operator_11_true_20_operator_11_true_20_and_nl,
          operator_11_true_25_operator_11_true_25_and_nl, return_add_generic_AC_RND_CONV_false_9_op1_inf_sva_1,
          operator_11_true_return_26_sva_2, operator_11_true_45_operator_11_true_45_and_nl,
          operator_11_true_44_operator_11_true_44_and_nl, operator_11_true_52_operator_11_true_52_and_nl,
          operator_11_true_57_operator_11_true_57_and_nl, {or_dcpl_88 , (fsm_output[9])
          , (fsm_output[10]) , (fsm_output[13]) , (fsm_output[14]) , or_934_nl ,
          (fsm_output[23]) , (fsm_output[25]) , (fsm_output[26]) , (fsm_output[29])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_x_im_d_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      stage_PE_1_x_im_d_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_390 | or_dcpl_338 | or_dcpl_388 | or_dcpl_387
        | or_dcpl_316 | or_dcpl_133 | or_dcpl_300)) ) begin
      stage_PE_1_x_im_d_sva <= MUX_v_64_2_2(out_f_d_rsci_q_d, in_f_d_rsci_q_d, fsm_output[21]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_mux_5_itm_13_10 <= 4'b0000;
    end
    else if ( rst ) begin
      BUTTERFLY_mux_5_itm_13_10 <= 4'b0000;
    end
    else if ( BUTTERFLY_and_ssc & (~ mode_lpi_1_dfm) ) begin
      BUTTERFLY_mux_5_itm_13_10 <= MUX_v_4_2_2((BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out[13:10]),
          (BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out[13:10]), inverse_lpi_1_dfm_1);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_mux_5_itm_9_0 <= 10'b0000000000;
    end
    else if ( rst ) begin
      BUTTERFLY_mux_5_itm_9_0 <= 10'b0000000000;
    end
    else if ( BUTTERFLY_and_ssc & (~(or_dcpl_102 | (fsm_output[26]) | (fsm_output[20])
        | or_dcpl_343 | (fsm_output[24]) | or_dcpl_340 | or_dcpl_98 | or_dcpl_87
        | (fsm_output[21]))) ) begin
      BUTTERFLY_mux_5_itm_9_0 <= MUX1HOT_v_10_4_2(BUTTERFLY_1_fry_9_0_sva, (z_out_49[9:0]),
          (BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out[9:0]), (BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out[9:0]),
          {nor_145_cse , (fsm_output[19]) , BUTTERFLY_and_5_nl , BUTTERFLY_and_6_nl});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_15_res_mant_or_1_cse
        | (fsm_output[31]) | or_dcpl_380 | or_dcpl_377 | (fsm_output[6]) | or_dcpl_106
        | (fsm_output[8]) | ((~ inverse_lpi_1_dfm_1) & (fsm_output[7])))) ) begin
      return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0 <= MUX1HOT_v_51_7_2((out_f_d_rsci_q_d[51:1]),
          (out_f_d_rsci_q_d[50:0]), (in_f_d_rsci_q_d[51:1]), (in_f_d_rsci_q_d[50:0]),
          return_add_generic_AC_RND_CONV_false_24_return_add_generic_AC_RND_CONV_false_24_and_4_nl,
          (z_out_34[51:1]), (~ (z_out_34[51:1])), {or_939_nl , or_940_nl , and_990_nl
          , and_992_nl , (fsm_output[30]) , return_add_generic_AC_RND_CONV_false_17_or_4_nl
          , return_add_generic_AC_RND_CONV_false_17_or_5_nl});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd <= 3'b000;
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_2_1 <= 2'b00;
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0 <= 1'b0;
    end
    else if ( rst ) begin
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd <= 3'b000;
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_2_1 <= 2'b00;
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0 <= 1'b0;
    end
    else if ( BUTTERFLY_1_else_1_if_and_ssc ) begin
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd <= MUX1HOT_v_3_3_2((out_u_rsci_q_d[15:13]),
          (in_u_rsci_q_d[15:13]), (BUTTERFLY_1_else_3_else_acc_4_sdt[15:13]), {BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c0
          , (fsm_output[22]) , (fsm_output[24])});
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_2_1 <= MUX1HOT_v_2_4_2((out_u_rsci_q_d[12:11]),
          (z_out_15[12:11]), (in_u_rsci_q_d[12:11]), (BUTTERFLY_1_else_3_else_acc_4_sdt[12:11]),
          {BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c0 , BUTTERFLY_else_1_if_or_3_cse
          , (fsm_output[22]) , (fsm_output[24])});
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0 <= MUX1HOT_s_1_7_2((out_u_rsci_q_d[10]),
          (z_out_15[10]), (in_u_rsci_q_d[10]), (BUTTERFLY_1_else_3_else_acc_4_sdt[10]),
          (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w0_10_1[9]), (stage_PE_1_tmp_im_d_1_sva_1_63_51[11]),
          (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w2_10_1[9]), {BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c0
          , BUTTERFLY_else_1_if_or_3_cse , (fsm_output[22]) , (fsm_output[24]) ,
          BUTTERFLY_else_1_if_and_cse , BUTTERFLY_else_1_if_and_1_cse , or_tmp_773});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_11_op_bigger_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm <= MUX1HOT_s_1_13_2(return_add_generic_AC_RND_CONV_false_4_op2_mu_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_4_op1_mu_0_lpi_3_dfm_1, return_mult_generic_AC_RND_CONV_false_1_if_nor_ovfl_sva_1,
          return_extract_12_return_extract_12_or_1_tmp, stage_PE_tmp_re_d_1_lpi_3_dfm_51_mx0,
          return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_3_nl,
          return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[50]),
          return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50, (return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0[50]),
          (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[50]), return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx6,
          return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0, {return_add_generic_AC_RND_CONV_false_11_op_bigger_and_4_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_5_cse , (fsm_output[8])
          , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_5_cse , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_6_cse
          , (fsm_output[10]) , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_13_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse});
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm <= MUX1HOT_s_1_9_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2,
          return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_2_cse, return_add_generic_AC_RND_CONV_false_14_op1_mu_mux_1_cse,
          return_add_generic_AC_RND_CONV_false_18_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_18_res_mant_3_0_sva_1),
          return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx6,
          return_add_generic_AC_RND_CONV_false_25_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_25_res_mant_3_0_sva_1),
          {(fsm_output[6]) , (fsm_output[10]) , (fsm_output[13]) , (fsm_output[14])
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse
          , (fsm_output[24]) , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_nl
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_nl});
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm <= MUX1HOT_v_50_8_2((return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1[49:0]),
          (return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1[50:1]), return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_1_cse_1,
          return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_2_cse, (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[49:0]),
          (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[50:1]), return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0,
          (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[49:0]),
          {return_add_generic_AC_RND_CONV_false_11_exp_and_1_cse , return_add_generic_AC_RND_CONV_false_11_exp_and_2_cse
          , (fsm_output[13]) , (fsm_output[14]) , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_13_cse , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_13_cse
          , and_1808_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_15_res_mant_4_sva <= 57'b000000000000000000000000000000000000000000000000000000000;
      return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_20_ls_sva <= 6'b000000;
      operator_6_false_18_acc_psp_sva_11 <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_15_res_mant_4_sva <= 57'b000000000000000000000000000000000000000000000000000000000;
      return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_20_ls_sva <= 6'b000000;
      operator_6_false_18_acc_psp_sva_11 <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_11_op_bigger_and_1_cse ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm <= MUX1HOT_s_1_10_2(return_add_generic_AC_RND_CONV_false_4_op2_mu_52_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_4_op1_mu_52_lpi_3_dfm_1, stage_PE_tmp_re_d_1_lpi_3_dfm_51_mx0,
          return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm,
          return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm, stage_PE_1_tmp_re_d_1_lpi_3_dfm_51_mx1,
          return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1, {return_add_generic_AC_RND_CONV_false_11_op_bigger_and_4_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_5_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_18_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_5_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_nl , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_11_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_24_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse});
      return_add_generic_AC_RND_CONV_false_15_res_mant_4_sva <= MUX1HOT_v_57_5_2((readslicef_58_57_1(acc_4_nl)),
          return_add_generic_AC_RND_CONV_false_5_res_mant_4_sva_1, return_add_generic_AC_RND_CONV_false_6_res_mant_4_sva_1,
          return_add_generic_AC_RND_CONV_false_8_res_mant_4_sva_1, z_out_9, {return_add_generic_AC_RND_CONV_false_15_res_mant_or_4_nl
          , (fsm_output[7]) , (fsm_output[10]) , (fsm_output[12]) , return_add_generic_AC_RND_CONV_false_15_res_mant_or_5_nl});
      return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva <= MUX1HOT_s_1_6_2(leading_sign_57_0_1_0_4_out_2,
          leading_sign_57_0_1_0_8_out_2, all_same_out, leading_sign_57_0_1_0_18_out_2,
          leading_sign_57_0_1_0_21_out_2, return_add_generic_AC_RND_CONV_false_25_exception_sva_1,
          {(fsm_output[7]) , (fsm_output[12]) , (fsm_output[14]) , (fsm_output[23])
          , (fsm_output[28]) , (fsm_output[30])});
      return_add_generic_AC_RND_CONV_false_20_ls_sva <= MUX1HOT_v_6_4_2(rtn_out,
          leading_sign_53_0_1_out_1, leading_sign_57_0_1_0_8_out_3, leading_sign_57_0_1_0_20_out_3,
          {return_add_generic_AC_RND_CONV_false_20_ls_or_cse , (fsm_output[8]) ,
          (fsm_output[12]) , (fsm_output[28])});
      operator_6_false_18_acc_psp_sva_11 <= MUX1HOT_s_1_3_2((z_out_50[11]), (return_add_generic_AC_RND_CONV_false_9_e_dif1_acc_1_tmp[11]),
          (return_add_generic_AC_RND_CONV_false_10_e_dif1_acc_1_tmp[11]), {operator_6_false_18_or_cse
          , (fsm_output[13]) , (fsm_output[14])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_41_return_extract_41_or_1_cse_sva <= 1'b0;
      stage_PE_1_gm_im_d_61_0_lpi_3_dfm <= 62'b00000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_extract_41_return_extract_41_or_1_cse_sva <= 1'b0;
      stage_PE_1_gm_im_d_61_0_lpi_3_dfm <= 62'b00000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( return_extract_41_and_1_cse ) begin
      return_extract_41_return_extract_41_or_1_cse_sva <= return_extract_41_return_extract_41_or_1_cse_sva_1;
      stage_PE_1_gm_im_d_61_0_lpi_3_dfm <= r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & ((~(and_dcpl_196 | or_dcpl_456 | or_dcpl_454 | (fsm_output[23])
        | (fsm_output[15]) | (fsm_output[9]))) | (fsm_output[6]) | (fsm_output[8])
        | (fsm_output[13]) | (fsm_output[14]) | (fsm_output[21])) ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm <= MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_4_op_bigger_mux_3_cse,
          return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_cse,
          return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_cse, return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0, {(fsm_output[6])
          , (fsm_output[8]) , (fsm_output[13]) , (fsm_output[14]) , (fsm_output[21])
          , (fsm_output[29])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_do_sub_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_do_sub_sva <= 1'b0;
    end
    else if ( run_wen & (~((fsm_output[26]) | (fsm_output[29]) | or_dcpl_471)) )
        begin
      return_add_generic_AC_RND_CONV_false_10_do_sub_sva <= MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_4_do_sub_sva_1,
          return_mult_generic_AC_RND_CONV_false_1_r_nan_sva_1, return_mult_generic_AC_RND_CONV_false_2_r_nan_sva_1,
          return_add_generic_AC_RND_CONV_false_10_do_sub_return_add_generic_AC_RND_CONV_false_10_do_sub_xor_nl,
          return_add_generic_AC_RND_CONV_false_5_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_19_do_sub_return_add_generic_AC_RND_CONV_false_19_do_sub_return_add_generic_AC_RND_CONV_false_19_do_sub_xnor_nl,
          return_mult_generic_AC_RND_CONV_false_5_r_nan_sva_1, return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_xnor_nl,
          {(fsm_output[6]) , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[12])
          , (fsm_output[22]) , (fsm_output[25]) , (fsm_output[27]) , (fsm_output[28])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_17_mux_6_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_17_mux_6_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_477 | or_dcpl_442)) ) begin
      return_add_generic_AC_RND_CONV_false_17_mux_6_itm <= MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_4_if_2_mux_nl,
          return_add_generic_AC_RND_CONV_false_12_if_2_mux_nl, fsm_output[29]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_89 | (fsm_output[7]) | or_dcpl_145 | (fsm_output[8])))
        & mode_lpi_1_dfm ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_itm <= MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_5_if_2_return_add_generic_AC_RND_CONV_false_5_if_2_and_2_nl,
          return_add_generic_AC_RND_CONV_false_5_r_sign_mux_1_nl, or_dcpl_474);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_mux_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_mux_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_396 | or_dcpl_338 | (fsm_output[25]) | (fsm_output[23])
        | or_dcpl_133)) ) begin
      return_add_generic_AC_RND_CONV_false_11_mux_itm <= MUX1HOT_s_1_15_2(return_add_generic_AC_RND_CONV_false_3_if_2_return_add_generic_AC_RND_CONV_false_3_if_2_nor_1_nl,
          (stage_PE_1_x_im_d_sva[63]), (~ (out_f_d_rsci_q_d[63])), return_add_generic_AC_RND_CONV_false_2_if_2_return_add_generic_AC_RND_CONV_false_2_if_2_nor_1_nl,
          (out_f_d_rsci_q_d[63]), (~ (stage_PE_1_tmp_im_d_1_sva_1_63_51[12])), return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_tmp,
          return_add_generic_AC_RND_CONV_false_11_if_2_return_add_generic_AC_RND_CONV_false_11_if_2_nor_mx3w0,
          (stage_PE_1_x_re_d_sva[63]), (~ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1),
          return_add_generic_AC_RND_CONV_false_14_if_2_return_add_generic_AC_RND_CONV_false_14_if_2_and_2_nl,
          (in_f_d_rsci_q_d[63]), return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp,
          return_add_generic_AC_RND_CONV_false_10_if_2_return_add_generic_AC_RND_CONV_false_10_if_2_and_1_mx3w0,
          operator_11_true_return_15_sva, {return_add_generic_AC_RND_CONV_false_11_and_25_nl
          , return_add_generic_AC_RND_CONV_false_11_or_4_nl , return_add_generic_AC_RND_CONV_false_11_and_36_nl
          , return_add_generic_AC_RND_CONV_false_11_and_27_cse , return_add_generic_AC_RND_CONV_false_11_and_37_cse
          , return_add_generic_AC_RND_CONV_false_11_and_38_cse , (fsm_output[10])
          , return_add_generic_AC_RND_CONV_false_10_and_4_cse , return_add_generic_AC_RND_CONV_false_10_and_16_cse
          , return_add_generic_AC_RND_CONV_false_10_and_17_cse , return_add_generic_AC_RND_CONV_false_11_and_31_nl
          , return_add_generic_AC_RND_CONV_false_11_and_42_nl , (fsm_output[26])
          , return_add_generic_AC_RND_CONV_false_11_and_33_nl , return_add_generic_AC_RND_CONV_false_11_and_44_nl});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_mux_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_mux_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_343 | or_dcpl_340 | or_dcpl_305 | (fsm_output[16:15]!=2'b00)))
        ) begin
      return_add_generic_AC_RND_CONV_false_12_mux_itm <= MUX1HOT_s_1_16_2(return_add_generic_AC_RND_CONV_false_5_do_sub_sva_1,
          return_add_generic_AC_RND_CONV_false_if_2_return_add_generic_AC_RND_CONV_false_if_2_and_2_nl,
          (out_f_d_rsci_q_d[63]), (stage_PE_1_tmp_im_d_1_sva_1_63_51[12]), return_add_generic_AC_RND_CONV_false_7_do_sub_return_add_generic_AC_RND_CONV_false_7_do_sub_xor_nl,
          (({return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0
          , return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx1
          , return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50_mx2
          , return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0_mx2
          , return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1})), return_add_generic_AC_RND_CONV_false_12_if_2_return_add_generic_AC_RND_CONV_false_12_if_2_nor_mx3w0,
          (stage_PE_1_x_im_d_sva[63]), (~ operator_11_true_return_15_sva), return_add_generic_AC_RND_CONV_false_15_if_2_return_add_generic_AC_RND_CONV_false_15_if_2_nor_1_nl,
          (in_f_d_rsci_q_d[63]), (~ (stage_PE_1_tmp_im_d_1_sva_1_63_51[12])), return_add_generic_AC_RND_CONV_false_20_do_sub_return_add_generic_AC_RND_CONV_false_20_do_sub_xor_nl,
          return_add_generic_AC_RND_CONV_false_11_if_2_return_add_generic_AC_RND_CONV_false_11_if_2_nor_mx3w0,
          (stage_PE_1_x_re_d_sva[63]), (~ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1),
          {(fsm_output[6]) , return_add_generic_AC_RND_CONV_false_11_and_27_cse ,
          return_add_generic_AC_RND_CONV_false_11_and_37_cse , return_add_generic_AC_RND_CONV_false_11_and_38_cse
          , (fsm_output[10]) , (fsm_output[13]) , return_add_generic_AC_RND_CONV_false_10_and_6_cse
          , return_add_generic_AC_RND_CONV_false_10_and_18_cse , return_add_generic_AC_RND_CONV_false_10_and_19_cse
          , return_add_generic_AC_RND_CONV_false_12_and_5_nl , return_add_generic_AC_RND_CONV_false_12_and_13_nl
          , return_add_generic_AC_RND_CONV_false_12_and_14_nl , (fsm_output[26])
          , return_add_generic_AC_RND_CONV_false_10_and_12_cse , return_add_generic_AC_RND_CONV_false_10_and_24_cse
          , return_add_generic_AC_RND_CONV_false_10_and_25_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 <= 1'b0;
    end
    else if ( return_extract_41_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 <= MUX1HOT_s_1_3_2(return_extract_50_and_nl,
          return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1, return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2,
          {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , (fsm_output[12])
          , (fsm_output[28])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_15_m_zero_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_15_m_zero_sva <= 1'b0;
    end
    else if ( run_wen & ((inverse_lpi_1_dfm_1 & (~(or_dcpl_390 | (fsm_output[27])
        | (fsm_output[25]) | (fsm_output[29]) | (fsm_output[22]) | or_dcpl_365)))
        | (fsm_output[6]) | (fsm_output[8]) | (fsm_output[12]) | (fsm_output[13])
        | (fsm_output[21])) ) begin
      return_extract_15_m_zero_sva <= MUX1HOT_s_1_5_2(return_extract_3_m_zero_sva_1,
          return_extract_15_m_zero_return_extract_15_m_zero_nor_nl, return_extract_17_m_zero_sva_mx0w3,
          return_extract_27_m_zero_return_extract_27_m_zero_nor_nl, return_extract_15_m_zero_mux1h_3_cse,
          {(fsm_output[6]) , (fsm_output[8]) , (fsm_output[12]) , (fsm_output[13])
          , return_extract_17_m_zero_or_2_nl});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_13_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_13_sva <= 1'b0;
    end
    else if ( run_wen & (~((fsm_output[24]) | (fsm_output[16]) | (fsm_output[14])
        | (fsm_output[8]))) ) begin
      operator_11_true_return_13_sva <= MUX1HOT_s_1_12_2(operator_11_true_return_3_sva_mx1w0,
          operator_11_true_13_operator_11_true_13_and_nl, return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp,
          return_add_generic_AC_RND_CONV_false_7_op1_inf_sva_1, return_mult_generic_AC_RND_CONV_false_2_lor_lpi_3_dfm_1,
          operator_11_true_53_operator_11_true_53_and_nl, operator_11_true_27_operator_11_true_27_and_nl,
          return_add_generic_AC_RND_CONV_false_10_op1_inf_sva_1, operator_11_true_return_26_sva_2,
          return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1, return_mult_generic_AC_RND_CONV_false_5_lor_lpi_3_dfm_1,
          operator_11_true_59_operator_11_true_59_and_nl, {(fsm_output[6]) , (fsm_output[7])
          , (fsm_output[9]) , (fsm_output[10]) , (fsm_output[11]) , BUTTERFLY_else_1_if_or_3_cse
          , (fsm_output[13]) , (fsm_output[15]) , or_dcpl_87 , (fsm_output[26]) ,
          (fsm_output[27]) , (fsm_output[29])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_13_do_sub_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_13_do_sub_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_367 | (fsm_output[13]) | or_dcpl_505)) ) begin
      return_add_generic_AC_RND_CONV_false_13_do_sub_sva <= MUX1HOT_s_1_7_2(return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1,
          return_add_generic_AC_RND_CONV_false_2_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_6_do_sub_return_add_generic_AC_RND_CONV_false_6_do_sub_return_add_generic_AC_RND_CONV_false_6_do_sub_xnor_nl,
          return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_xnor_nl,
          return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_13_do_sub_sva_1,
          return_add_generic_AC_RND_CONV_false_21_do_sub_return_add_generic_AC_RND_CONV_false_21_do_sub_xor_nl,
          {(fsm_output[6]) , (fsm_output[8]) , (fsm_output[9]) , (fsm_output[12])
          , (fsm_output[22]) , (fsm_output[24]) , (fsm_output[26])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_15_do_sub_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_15_do_sub_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_305 | (fsm_output[29]) | (fsm_output[15]))) )
        begin
      return_add_generic_AC_RND_CONV_false_15_do_sub_sva <= MUX1HOT_s_1_7_2(return_add_generic_AC_RND_CONV_false_3_do_sub_sva_1,
          return_add_generic_AC_RND_CONV_false_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_8_do_sub_return_add_generic_AC_RND_CONV_false_8_do_sub_xor_nl,
          return_add_generic_AC_RND_CONV_false_7_op1_nan_sva_1, return_add_generic_AC_RND_CONV_false_16_do_sub_sva_1,
          return_add_generic_AC_RND_CONV_false_15_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_22_do_sub_return_add_generic_AC_RND_CONV_false_22_do_sub_xor_nl,
          {(fsm_output[6]) , (fsm_output[8]) , (fsm_output[10]) , (fsm_output[14])
          , (fsm_output[22]) , (fsm_output[24]) , (fsm_output[28])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm
          <= 51'b000000000000000000000000000000000000000000000000000;
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_63 <= 1'b0;
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_51 <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm
          <= 51'b000000000000000000000000000000000000000000000000000;
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_63 <= 1'b0;
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_51 <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_14_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm
          <= MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
          return_add_generic_AC_RND_CONV_false_14_mux1h_8_nl, nor_157_nl);
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_63 <= MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_11_mux_19_cse,
          stage_d_mul_return_d_2_63_sva_1, (stage_PE_1_tmp_im_d_1_sva_1_63_51[12]),
          return_add_generic_AC_RND_CONV_false_10_mux_7_itm, stage_d_mul_return_d_5_63_sva_1,
          {(fsm_output[7]) , (fsm_output[10]) , stage_PE_1_tmp_im_d_and_5_nl , stage_PE_1_tmp_im_d_and_6_cse
          , (fsm_output[26])});
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_51 <= MUX1HOT_s_1_4_2(stage_PE_tmp_im_d_1_lpi_3_dfm_51_mx0,
          stage_d_mul_return_d_1_63_sva_1, stage_PE_1_tmp_im_d_1_lpi_3_dfm_51_mx1,
          stage_d_mul_return_d_63_sva_1, {(fsm_output[7]) , (fsm_output[10]) , (fsm_output[23])
          , (fsm_output[26])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_tmp_im_d_1_sva_1_63_51 <= 13'b0000000000000;
    end
    else if ( rst ) begin
      stage_PE_1_tmp_im_d_1_sva_1_63_51 <= 13'b0000000000000;
    end
    else if ( stage_PE_1_tmp_im_d_and_ssc ) begin
      stage_PE_1_tmp_im_d_1_sva_1_63_51 <= MUX_v_13_2_2((out_f_d_rsci_q_d[63:51]),
          (in_f_d_rsci_q_d[63:51]), or_dcpl_87);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_tmp_im_d_1_sva_1_50_0 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      stage_PE_1_tmp_im_d_1_sva_1_50_0 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( stage_PE_1_tmp_im_d_and_ssc & (inverse_lpi_1_dfm_1 | or_dcpl_35 | or_dcpl_87)
        ) begin
      stage_PE_1_tmp_im_d_1_sva_1_50_0 <= MUX1HOT_v_51_4_2((out_f_d_rsci_q_d[50:0]),
          stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0w0, stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx0w2,
          (in_f_d_rsci_q_d[50:0]), {or_dcpl_35 , stage_PE_1_x_im_d_and_1_nl , or_tmp_773
          , or_dcpl_87});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd <= 1'b0;
      return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd <= 1'b0;
      return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_7_exp_and_ssc ) begin
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd <= MUX_s_1_2_2((return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
          (return_mult_generic_AC_RND_CONV_false_4_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
          fsm_output[24]);
      return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm <= MUX_v_51_2_2(return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1,
          return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1, fsm_output[24]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1 <= 4'b0000;
    end
    else if ( rst ) begin
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1 <= 4'b0000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_7_exp_and_ssc & (~((fsm_output[16])
        | (fsm_output[7]) | (fsm_output[15]))) ) begin
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1 <= MUX1HOT_v_4_3_2(and_2119_nl, (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1[9:6]),
          (return_mult_generic_AC_RND_CONV_false_4_exp_1_11_0_lpi_3_dfm_3_10_0_1[9:6]),
          {drf_qr_lval_10_smx_lpi_3_dfm_mx0c0 , (fsm_output[10]) , (fsm_output[24])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2 <= 6'b000000;
    end
    else if ( rst ) begin
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2 <= 6'b000000;
    end
    else if ( (mux_22_nl | (fsm_output[30]) | (fsm_output[29]) | (fsm_output[14])
        | (fsm_output[13]) | (fsm_output[22]) | (fsm_output[6]) | (fsm_output[23])
        | (fsm_output[24]) | (fsm_output[10])) & run_wen ) begin
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2 <= MUX1HOT_v_6_5_2(and_2131_nl, (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1[5:0]),
          drf_qr_lval_10_smx_lpi_3_dfm_mx1_5_0, (return_mult_generic_AC_RND_CONV_false_4_exp_1_11_0_lpi_3_dfm_3_10_0_1[5:0]),
          drf_qr_lval_10_smx_lpi_3_dfm_mx2_5_0, {drf_qr_lval_10_smx_lpi_3_dfm_mx0c0
          , (fsm_output[10]) , (fsm_output[12]) , (fsm_output[24]) , (fsm_output[28])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_else_2_acc_1_psp_16_0_sva_16_11 <= 6'b000000;
    end
    else if ( rst ) begin
      BUTTERFLY_else_2_acc_1_psp_16_0_sva_16_11 <= 6'b000000;
    end
    else if ( BUTTERFLY_else_2_and_ssc & (mode_lpi_1_dfm | (~ inverse_lpi_1_dfm_1))
        ) begin
      BUTTERFLY_else_2_acc_1_psp_16_0_sva_16_11 <= z_out_58[16:11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0 <= 11'b00000000000;
    end
    else if ( rst ) begin
      BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0 <= 11'b00000000000;
    end
    else if ( BUTTERFLY_else_2_and_ssc & ((~(or_dcpl_338 | (fsm_output[10]) | (and_dcpl_219
        & (fsm_output[28])) | (and_dcpl_220 & (fsm_output[12])))) | or_954_rgt |
        or_955_rgt | or_956_cse | (fsm_output[9]) | or_959_rgt | or_960_rgt | (fsm_output[26])
        | BUTTERFLY_else_2_and_2_rgt) ) begin
      BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0 <= MUX1HOT_v_11_8_2((out_f_d_rsci_q_d[62:52]),
          (stage_PE_1_x_im_d_sva[62:52]), (stage_PE_1_tmp_im_d_1_sva_1_63_51[11:1]),
          return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w3,
          return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1,
          (in_f_d_rsci_q_d[62:52]), return_mult_generic_AC_RND_CONV_false_3_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w7,
          (z_out_58[10:0]), {or_954_rgt , or_955_rgt , or_956_cse , (fsm_output[9])
          , BUTTERFLY_else_2_and_8_nl , or_960_rgt , (fsm_output[26]) , BUTTERFLY_else_2_and_2_rgt});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~(BUTTERFLY_if_1_or_3_cse | return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_2_cse))
        ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0 <= MUX1HOT_v_51_11_2(return_add_generic_AC_RND_CONV_false_4_op1_mu_51_1_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_4_op2_mu_51_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_mx0w2,
          return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_mx0w4, return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_mx0w5,
          return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_mx0w6, return_add_generic_AC_RND_CONV_false_25_return_add_generic_AC_RND_CONV_false_25_and_4_nl,
          (z_out_34[51:1]), (~ (z_out_34[51:1])), (~ (return_add_generic_AC_RND_CONV_false_25_rshift_itm[51:1])),
          (return_add_generic_AC_RND_CONV_false_25_rshift_itm[51:1]), {or_tmp_388
          , or_tmp_389 , (fsm_output[8]) , (fsm_output[13]) , (fsm_output[24]) ,
          return_add_generic_AC_RND_CONV_false_18_and_15_nl , (fsm_output[30]) ,
          return_add_generic_AC_RND_CONV_false_11_op_smaller_and_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse
          , and_304_nl , return_add_generic_AC_RND_CONV_false_18_and_4_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_1_m_zero_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_1_m_zero_sva <= 1'b0;
    end
    else if ( run_wen & ((~(inverse_lpi_1_dfm_1 | or_tmp_543)) | (fsm_output[7])
        | (fsm_output[24])) ) begin
      return_extract_1_m_zero_sva <= MUX_s_1_2_2(return_extract_3_m_zero_sva_1, return_extract_54_m_zero_return_extract_54_m_zero_nor_nl,
          fsm_output[24]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & (~ (fsm_output[9])) ) begin
      return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm <= MUX1HOT_s_1_7_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_mx0w1, return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1,
          {(fsm_output[7]) , (fsm_output[8]) , (fsm_output[13]) , (fsm_output[23])
          , (fsm_output[25]) , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_13_cse
          , and_1808_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50 <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50 <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_511) ) begin
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50 <= MUX1HOT_s_1_4_2(return_extract_13_return_extract_13_or_1_cse_sva_1,
          stage_PE_tmp_im_d_1_lpi_3_dfm_51_mx0, return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50_mx2,
          return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_mx0w1, {return_add_generic_AC_RND_CONV_false_19_op2_mu_and_2_nl
          , return_add_generic_AC_RND_CONV_false_19_op2_mu_and_3_nl , (fsm_output[13])
          , (fsm_output[24])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm <= 1'b0;
    end
    else if ( rst ) begin
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_338 | (fsm_output[8]))) ) begin
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm <= MUX1HOT_s_1_12_2(return_extract_13_return_extract_13_or_1_cse_sva_1,
          return_extract_12_return_extract_12_or_1_tmp, BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx1,
          (BUTTERFLY_1_fry_9_0_sva[9]), reg_BUTTERFLY_1_i_9_0_ftd, drf_qr_lval_14_smx_0_lpi_3_dfm,
          (return_add_generic_AC_RND_CONV_false_20_ls_sva[0]), return_extract_45_return_extract_45_or_1_cse_sva_1,
          return_extract_44_return_extract_44_or_1_tmp, BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx3,
          return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1, (stage_PE_1_x_re_d_sva[52]),
          {(fsm_output[7]) , (fsm_output[9]) , (fsm_output[10]) , or_1195_nl , or_tmp_567
          , BUTTERFLY_1_fiy_and_1_nl , BUTTERFLY_1_fiy_and_2_nl , (fsm_output[23])
          , (fsm_output[25]) , (fsm_output[26]) , BUTTERFLY_1_fiy_and_4_cse , BUTTERFLY_1_fiy_and_5_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_12_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      drf_qr_lval_12_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_89 | (fsm_output[16]) | or_dcpl_551 | (fsm_output[8])))
        ) begin
      drf_qr_lval_12_smx_0_lpi_3_dfm <= MUX1HOT_s_1_10_2(return_add_generic_AC_RND_CONV_false_1_r_nan_or_1_nl,
          (return_add_generic_AC_RND_CONV_false_1_res_rounded_lpi_3_dfm_51_0_1[51]),
          return_add_generic_AC_RND_CONV_false_9_exp_mux1h_2_cse, return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm,
          (stage_PE_1_x_im_d_sva[52]), return_add_generic_AC_RND_CONV_false_14_r_nan_or_1_nl,
          return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1, (stage_PE_1_x_re_d_sva[52]),
          return_add_generic_AC_RND_CONV_false_23_r_nan_or_1_nl, (return_add_generic_AC_RND_CONV_false_23_res_rounded_lpi_3_dfm_51_0_1[51]),
          {return_add_generic_AC_RND_CONV_false_9_exp_and_1_nl , return_add_generic_AC_RND_CONV_false_9_exp_or_nl
          , (fsm_output[13]) , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_11_cse , return_add_generic_AC_RND_CONV_false_9_exp_and_5_nl
          , return_add_generic_AC_RND_CONV_false_9_exp_and_7_nl , and_1134_cse ,
          return_add_generic_AC_RND_CONV_false_9_exp_and_9_nl , return_add_generic_AC_RND_CONV_false_9_exp_and_10_nl});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_itm
          <= 10'b0000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_itm
          <= 10'b0000000000;
    end
    else if ( run_wen & (~((fsm_output[32]) | (fsm_output[24]) | (fsm_output[25])
        | or_dcpl_300)) ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_itm
          <= MUX_v_10_2_2(mux_25_nl, 10'b1111111111, or_1772_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm
          <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm
          <= 1'b0;
    end
    else if ( (((~(return_add_generic_AC_RND_CONV_false_10_ma1_lt_ma2_acc_1_itm_52
        & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_sva)) & (fsm_output[14])
        & (~ (return_add_generic_AC_RND_CONV_false_10_e_dif1_acc_1_tmp[11]))) | (fsm_output[13])
        | (fsm_output[10]) | (fsm_output[7]) | (fsm_output[23]) | (fsm_output[29])
        | (fsm_output[30])) & run_wen ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm
          <= MUX1HOT_s_1_7_2(return_add_generic_AC_RND_CONV_false_1_e_r_return_add_generic_AC_RND_CONV_false_1_e_r_or_1_nl,
          return_add_generic_AC_RND_CONV_false_6_exp_plus_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm_mx1,
          return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_nl,
          return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_25_e_r_qelse_return_add_generic_AC_RND_CONV_false_25_e_r_qelse_and_1_nl,
          {(fsm_output[7]) , (fsm_output[10]) , (fsm_output[13]) , (fsm_output[14])
          , (fsm_output[23]) , (fsm_output[29]) , (fsm_output[30])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_cse_sva
          <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_cse_sva
          <= 1'b0;
    end
    else if ( run_wen & (~((fsm_output[24]) | (fsm_output[9]) | (fsm_output[8])))
        ) begin
      return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_cse_sva
          <= MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_1_return_add_generic_AC_RND_CONV_false_6_op2_normal_return_extract_13_nor_tmp,
          return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_tmp,
          return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp,
          {(fsm_output[7]) , (fsm_output[23]) , (fsm_output[25])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_12_m_zero_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_12_m_zero_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_571 | or_dcpl_388 | (fsm_output[29]) | (fsm_output[8])))
        ) begin
      return_extract_12_m_zero_sva <= MUX1HOT_s_1_6_2(return_extract_13_m_zero_return_extract_13_m_zero_nor_nl,
          return_extract_12_m_zero_return_extract_12_m_zero_nor_nl, return_extract_20_m_zero_return_extract_20_m_zero_nor_nl,
          return_extract_25_m_zero_return_extract_25_m_zero_nor_nl, return_extract_15_m_zero_mux1h_3_cse,
          return_add_generic_AC_RND_CONV_false_17_e_r_qelse_or_svs_1, {(fsm_output[7])
          , (fsm_output[9]) , (fsm_output[10]) , (fsm_output[13]) , or_1266_cse ,
          (fsm_output[23])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~ or_tmp_606) ) begin
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0 <= MUX_v_51_2_2(stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0,
          stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx1, fsm_output[23]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_24_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_24_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_354 | or_dcpl_325 | (fsm_output[10]) | or_dcpl_551))
        ) begin
      operator_11_true_return_24_sva <= MUX1HOT_s_1_3_2(operator_11_true_return_3_sva_mx1w0,
          return_add_generic_AC_RND_CONV_false_7_op1_inf_sva_1, operator_11_true_return_26_sva_2,
          {(fsm_output[8]) , (fsm_output[14]) , (fsm_output[24])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_17_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_17_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_571 | or_dcpl_388 | (fsm_output[10]) | (fsm_output[15])))
        ) begin
      operator_11_true_return_17_sva <= MUX1HOT_s_1_4_2(operator_11_true_17_operator_11_true_17_and_nl,
          operator_11_true_22_operator_11_true_22_and_nl, return_add_generic_AC_RND_CONV_false_9_op1_nan_sva_1,
          operator_11_true_54_operator_11_true_54_and_nl, {(fsm_output[8]) , (fsm_output[9])
          , (fsm_output[14]) , (fsm_output[24])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_15_return_extract_15_nor_cse_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_extract_15_return_extract_15_nor_cse_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( return_extract_15_and_3_cse ) begin
      return_extract_15_return_extract_15_nor_cse_sva <= MUX_s_1_2_2(return_extract_15_return_extract_15_nor_nl,
          return_extract_47_return_extract_47_nor_nl, fsm_output[24]);
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0 <= MUX1HOT_v_50_3_2((stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0[50:1]),
          (stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0[49:0]), return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0_mx2,
          {return_add_generic_AC_RND_CONV_false_19_op2_mu_return_add_generic_AC_RND_CONV_false_19_op2_mu_nor_nl
          , return_add_generic_AC_RND_CONV_false_19_op2_mu_and_5_nl , (fsm_output[13])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_15_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_15_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_98 | (fsm_output[16]) | (fsm_output[13]) | (fsm_output[9])))
        ) begin
      operator_11_true_return_15_sva <= MUX1HOT_s_1_7_2(operator_11_true_15_operator_11_true_15_and_nl,
          return_add_generic_AC_RND_CONV_false_7_op1_nan_sva_1, operator_11_true_return_15_sva_mx1,
          return_add_generic_AC_RND_CONV_false_10_op1_nan_sva_1, operator_11_true_47_operator_11_true_47_and_nl,
          return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1, operator_11_true_return_15_sva_mx2,
          {(fsm_output[8]) , (fsm_output[10]) , (fsm_output[12]) , (fsm_output[15])
          , (fsm_output[24]) , (fsm_output[26]) , (fsm_output[28])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & (~ and_1747_cse) ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm <= MUX1HOT_s_1_6_2(return_extract_15_return_extract_15_or_1_nl,
          return_add_generic_AC_RND_CONV_false_11_op_smaller_mux_cse, return_add_generic_AC_RND_CONV_false_10_op1_mu_mux_1_cse,
          return_extract_47_return_extract_47_or_1_nl, return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0,
          (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[50]), {(fsm_output[8])
          , (fsm_output[13]) , (fsm_output[14]) , (fsm_output[24]) , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_13_cse
          , and_1808_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_89) ) begin
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm <= MUX1HOT_s_1_11_2(return_extract_17_return_extract_17_or_sva_1,
          return_mult_generic_AC_RND_CONV_false_1_or_nl, return_mult_generic_AC_RND_CONV_false_2_or_nl,
          return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx1, return_add_generic_AC_RND_CONV_false_18_res_mant_3_0_sva_1,
          (~ return_add_generic_AC_RND_CONV_false_18_res_mant_3_0_sva_1), return_extract_45_return_extract_45_or_1_cse_sva_1,
          stage_PE_1_tmp_im_d_1_lpi_3_dfm_51_mx1, return_mult_generic_AC_RND_CONV_false_5_or_nl,
          return_add_generic_AC_RND_CONV_false_24_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_24_res_mant_3_0_sva_1),
          {(fsm_output[8]) , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[13])
          , return_add_generic_AC_RND_CONV_false_17_and_7_cse , return_add_generic_AC_RND_CONV_false_17_and_8_cse
          , return_add_generic_AC_RND_CONV_false_10_op2_mu_and_3_nl , return_add_generic_AC_RND_CONV_false_10_op2_mu_and_4_nl
          , (fsm_output[27]) , return_add_generic_AC_RND_CONV_false_17_and_9_cse
          , return_add_generic_AC_RND_CONV_false_17_and_3_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_14_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      drf_qr_lval_14_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & (~((fsm_output[26]) | (fsm_output[31]) | or_dcpl_338 | (fsm_output[25])
        | (fsm_output[14]) | (fsm_output[15]))) ) begin
      drf_qr_lval_14_smx_0_lpi_3_dfm <= MUX1HOT_s_1_9_2(return_add_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_1,
          (return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1[50]), BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx1,
          return_add_generic_AC_RND_CONV_false_9_exp_mux1h_2_cse, return_add_generic_AC_RND_CONV_false_18_return_add_generic_AC_RND_CONV_false_18_and_5_nl,
          return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_2_nl,
          return_add_generic_AC_RND_CONV_false_10_op1_mu_mux1h_3_cse, return_add_generic_AC_RND_CONV_false_24_r_nan_or_1_nl,
          (return_add_generic_AC_RND_CONV_false_24_res_rounded_lpi_3_dfm_51_0_1[51]),
          {(fsm_output[8]) , return_add_generic_AC_RND_CONV_false_11_exp_and_1_cse
          , return_add_generic_AC_RND_CONV_false_11_exp_and_2_cse , (fsm_output[13])
          , (fsm_output[23]) , (fsm_output[24]) , (fsm_output[29]) , return_add_generic_AC_RND_CONV_false_11_exp_and_3_nl
          , return_add_generic_AC_RND_CONV_false_11_exp_and_4_nl});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_and_1_itm
          <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_and_1_itm
          <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_17_m_r_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm <= MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_4_m_r_51_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm_mx1, return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_and_8_nl,
          return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm_mx2, {(fsm_output[8])
          , (fsm_output[13]) , (fsm_output[23]) , (fsm_output[29])});
      return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_and_1_itm
          <= MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nor_nl,
          return_add_generic_AC_RND_CONV_false_23_e_r_return_add_generic_AC_RND_CONV_false_23_e_r_or_1_nl,
          return_add_generic_AC_RND_CONV_false_24_e_r_return_add_generic_AC_RND_CONV_false_24_e_r_or_1_nl,
          {(fsm_output[8]) , (fsm_output[23]) , (fsm_output[30]) , (fsm_output[31])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm
          <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm
          <= 1'b0;
    end
    else if ( run_wen & (~ (fsm_output[32])) ) begin
      return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm
          <= MUX1HOT_s_1_7_2(return_extract_17_return_extract_17_nor_tmp, z_out_20_11,
          return_add_generic_AC_RND_CONV_false_6_if_5_return_add_generic_AC_RND_CONV_false_6_if_5_and_nl,
          return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_nor_nl,
          return_add_generic_AC_RND_CONV_false_24_e_r_qelse_return_add_generic_AC_RND_CONV_false_24_e_r_qelse_and_1_nl,
          return_add_generic_AC_RND_CONV_false_25_e_r_return_add_generic_AC_RND_CONV_false_25_e_r_or_1_nl,
          {(fsm_output[8]) , return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_2_cse
          , (fsm_output[10]) , (fsm_output[13]) , (fsm_output[23]) , (fsm_output[30])
          , (fsm_output[31])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_22_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_22_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_571 | or_dcpl_388 | or_dcpl_106)) ) begin
      return_add_generic_AC_RND_CONV_false_22_unequal_tmp <= MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp,
          return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp,
          fsm_output[24]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_456 | or_dcpl_454 | or_dcpl_145)) ) begin
      return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm <= MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_1_op2_mu_51_1_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm_mx1, fsm_output[21]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_x_re_d_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      stage_PE_1_x_re_d_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~ or_tmp_543) ) begin
      stage_PE_1_x_re_d_sva <= MUX_v_64_2_2(out_f_d_rsci_q_d, in_f_d_rsci_q_d, fsm_output[24]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_21_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_21_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_437 | or_dcpl_443)) ) begin
      return_add_generic_AC_RND_CONV_false_21_unequal_tmp <= MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_nl,
          return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp,
          return_add_generic_AC_RND_CONV_false_24_exception_sva_1, {(fsm_output[9])
          , (fsm_output[24]) , (fsm_output[30])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_op2_nan_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_op2_nan_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_124 | (fsm_output[16]) | (fsm_output[10]))) )
        begin
      return_add_generic_AC_RND_CONV_false_10_op2_nan_sva <= MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_14_op2_nan_sva_1,
          return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1, return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1,
          {(fsm_output[9]) , (fsm_output[15]) , (fsm_output[24])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_op2_inf_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_op2_inf_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_125 | or_dcpl_147 | (fsm_output[10]))) ) begin
      return_add_generic_AC_RND_CONV_false_10_op2_inf_sva <= MUX1HOT_s_1_5_2(return_mult_generic_AC_RND_CONV_false_op1_zero_sva_1,
          return_add_generic_AC_RND_CONV_false_9_do_sub_return_add_generic_AC_RND_CONV_false_9_do_sub_xor_nl,
          return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1, return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1,
          return_add_generic_AC_RND_CONV_false_23_do_sub_return_add_generic_AC_RND_CONV_false_23_do_sub_xor_nl,
          {(fsm_output[9]) , (fsm_output[12]) , (fsm_output[15]) , (fsm_output[24])
          , (fsm_output[28])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_do_sub_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_do_sub_sva <= 1'b0;
    end
    else if ( run_wen & (~((fsm_output[29]) | (fsm_output[16]) | (fsm_output[13])
        | or_dcpl_133)) ) begin
      return_add_generic_AC_RND_CONV_false_12_do_sub_sva <= MUX1HOT_s_1_4_2(z_out_20_11,
          return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_xnor_nl,
          return_add_generic_AC_RND_CONV_false_4_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_xnor_nl,
          {return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_2_cse , (fsm_output[12])
          , (fsm_output[22]) , (fsm_output[28])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_else_2_tmp2_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      BUTTERFLY_1_else_2_tmp2_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & (~ mode_lpi_1_dfm) ) begin
      BUTTERFLY_1_else_2_tmp2_1_sva <= z_out_25;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm <= 1'b0;
    end
    else if ( run_wen & ((~(and_dcpl_228 | or_dcpl_353 | or_dcpl_523 | (fsm_output[15])))
        | (fsm_output[10]) | (fsm_output[13]) | (fsm_output[14]) | (fsm_output[24]))
        ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm <= MUX1HOT_s_1_7_2(return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_2_nl,
          return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm,
          return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm,
          return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0,
          {(fsm_output[10]) , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_11_cse , (fsm_output[24])
          , (fsm_output[29])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd
          <= 1'b0;
    end
    else if ( rst ) begin
      reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd
          <= 1'b0;
    end
    else if ( run_wen & (~ leading_sign_57_0_1_0_18_out_2) & mode_lpi_1_dfm ) begin
      reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd
          <= return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_1[50];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1
          <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1
          <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_338 | (fsm_output[15]))) ) begin
      reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1
          <= MUX1HOT_v_50_14_2((stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0[49:0]), (stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0[50:1]),
          (return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1[50:1]), (return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1[49:0]),
          return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[49:0]),
          return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0, (return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0[49:0]),
          (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1[49:0]), (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1[50:1]),
          (return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1[50:1]), (return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1[49:0]),
          return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_1[49:0]),
          {return_add_generic_AC_RND_CONV_false_14_op1_mu_and_6_cse , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_5_cse
          , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_8_cse , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_7_cse
          , and_1132_ssc , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse
          , and_1804_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_cse
          , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_2_cse , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_1_cse
          , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_12_cse , return_add_generic_AC_RND_CONV_false_14_op1_mu_and_11_cse
          , and_1145_ssc , (fsm_output[23])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      in_u_rsc_merge_sva_rsp_0 <= 6'b000000;
      in_u_rsc_merge_sva_rsp_1_rsp_0 <= 4'b0000;
      in_u_rsc_merge_sva_rsp_1_rsp_1 <= 6'b000000;
    end
    else if ( rst ) begin
      in_u_rsc_merge_sva_rsp_0 <= 6'b000000;
      in_u_rsc_merge_sva_rsp_1_rsp_0 <= 4'b0000;
      in_u_rsc_merge_sva_rsp_1_rsp_1 <= 6'b000000;
    end
    else if ( in_u_and_ssc ) begin
      in_u_rsc_merge_sva_rsp_0 <= MUX1HOT_v_6_4_2((out_u_rsci_q_d[15:10]), (in_u_mux1h_1_itm[15:10]),
          (in_u_rsci_q_d[15:10]), (z_out_64_31_16[15:10]), {(fsm_output[7]) , (fsm_output[10])
          , (fsm_output[21]) , (fsm_output[23])});
      in_u_rsc_merge_sva_rsp_1_rsp_0 <= MUX1HOT_v_4_5_2((out_u_rsci_q_d[9:6]), (in_u_mux1h_1_itm[9:6]),
          or_1486_nl, (in_u_rsci_q_d[9:6]), (z_out_64_31_16[9:6]), {(fsm_output[7])
          , (fsm_output[10]) , in_u_rsc_merge_sva_mx0c2 , (fsm_output[21]) , (fsm_output[23])});
      in_u_rsc_merge_sva_rsp_1_rsp_1 <= MUX1HOT_v_6_5_2((out_u_rsci_q_d[5:0]), (in_u_mux1h_1_itm[5:0]),
          or_1487_nl, (in_u_rsci_q_d[5:0]), (z_out_64_31_16[5:0]), {(fsm_output[7])
          , (fsm_output[10]) , in_u_rsc_merge_sva_mx0c2 , (fsm_output[21]) , (fsm_output[23])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_6_false_18_acc_psp_sva_10_0_rsp_0 <= 1'b0;
      operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0 <= 9'b000000000;
      operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1 <= 1'b0;
    end
    else if ( rst ) begin
      operator_6_false_18_acc_psp_sva_10_0_rsp_0 <= 1'b0;
      operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0 <= 9'b000000000;
      operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1 <= 1'b0;
    end
    else if ( operator_6_false_18_and_1_ssc ) begin
      operator_6_false_18_acc_psp_sva_10_0_rsp_0 <= MUX1HOT_s_1_4_2((operator_6_false_18_mux1h_itm_10_1[9]),
          (z_out_50[10]), (return_add_generic_AC_RND_CONV_false_9_e_dif1_acc_1_tmp[10]),
          (return_add_generic_AC_RND_CONV_false_10_e_dif1_acc_1_tmp[10]), {or_1285_itm
          , operator_6_false_18_or_cse , (fsm_output[13]) , (fsm_output[14])});
      operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0 <= MUX1HOT_v_9_5_2((operator_6_false_18_mux1h_itm_10_1[8:0]),
          (return_add_generic_AC_RND_CONV_false_6_exp_plus_1_12_1_lpi_3_dfm_1[9:1]),
          (z_out_50[9:1]), (return_add_generic_AC_RND_CONV_false_9_e_dif1_acc_1_tmp[9:1]),
          (return_add_generic_AC_RND_CONV_false_10_e_dif1_acc_1_tmp[9:1]), {or_1285_itm
          , (fsm_output[10]) , operator_6_false_18_or_cse , (fsm_output[13]) , (fsm_output[14])});
      operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1 <= MUX1HOT_s_1_5_2(and_2118_nl,
          (return_add_generic_AC_RND_CONV_false_6_exp_plus_1_12_1_lpi_3_dfm_1[0]),
          (z_out_50[0]), (return_add_generic_AC_RND_CONV_false_9_e_dif1_acc_1_tmp[0]),
          (return_add_generic_AC_RND_CONV_false_10_e_dif1_acc_1_tmp[0]), {or_1285_itm
          , (fsm_output[10]) , operator_6_false_18_or_cse , (fsm_output[13]) , (fsm_output[14])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_u_add_3_acc_itm_rsp_0 <= 4'b0000;
      stage_u_add_3_acc_itm_rsp_1 <= 13'b0000000000000;
    end
    else if ( rst ) begin
      stage_u_add_3_acc_itm_rsp_0 <= 4'b0000;
      stage_u_add_3_acc_itm_rsp_1 <= 13'b0000000000000;
    end
    else if ( stage_u_add_3_and_ssc ) begin
      stage_u_add_3_acc_itm_rsp_0 <= MUX1HOT_v_4_3_2((z_out_1[16:13]), (stage_u_add_3_mux1h_2_itm[16:13]),
          (z_out_22[16:13]), {(fsm_output[8]) , (fsm_output[11]) , stage_u_add_3_or_1_cse});
      stage_u_add_3_acc_itm_rsp_1 <= MUX1HOT_v_13_7_2((z_out_1[12:0]), return_mult_generic_AC_RND_CONV_false_1_exp_acc_tmp,
          operator_33_true_12_acc_tmp, z_out_16, (z_out_48[12:0]), (stage_u_add_3_mux1h_2_itm[12:0]),
          (z_out_22[12:0]), {stage_u_add_3_and_1_nl , stage_u_add_3_and_3_nl , (fsm_output[10])
          , operator_14_false_1_or_nl , (fsm_output[15]) , (fsm_output[11]) , stage_u_add_3_or_1_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0 <= 9'b000000000;
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1 <= 1'b0;
    end
    else if ( rst ) begin
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0 <= 9'b000000000;
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1 <= 1'b0;
    end
    else if ( and_2620_ssc ) begin
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0 <= MUX1HOT_v_9_8_2((out_u_rsci_q_d[9:1]),
          (z_out_15[9:1]), (and_2143_itm[9:1]), (in_u_rsci_q_d[9:1]), (BUTTERFLY_1_else_3_else_acc_4_sdt[9:1]),
          (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w0_10_1[8:0]), (stage_PE_1_tmp_im_d_1_sva_1_63_51[10:2]),
          (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w2_10_1[8:0]), {BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c0
          , BUTTERFLY_else_1_if_or_3_cse , or_965_itm , (fsm_output[22]) , (fsm_output[24])
          , BUTTERFLY_else_1_if_and_cse , BUTTERFLY_else_1_if_and_1_cse , BUTTERFLY_else_1_if_and_5_cse});
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1 <= MUX1HOT_s_1_8_2((out_u_rsci_q_d[0]),
          (z_out_15[0]), (and_2143_itm[0]), (in_u_rsci_q_d[0]), (BUTTERFLY_1_else_3_else_acc_4_sdt[0]),
          stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w0_0, (stage_PE_1_tmp_im_d_1_sva_1_63_51[1]),
          stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w2_0, {BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_mx0c0
          , BUTTERFLY_else_1_if_or_3_cse , or_965_itm , (fsm_output[22]) , (fsm_output[24])
          , BUTTERFLY_else_1_if_and_cse , BUTTERFLY_else_1_if_and_1_cse , BUTTERFLY_else_1_if_and_5_cse});
    end
  end
  assign nl_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_acc_nl = return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3
      + 11'b00000000001;
  assign return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_acc_nl = nl_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_acc_nl[10:0];
  assign return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl = (~ return_mult_generic_AC_RND_CONV_false_6_e_incr_lpi_2_dfm_2)
      & return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_6_else_2_else_mux_nl = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_acc_nl,
      return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3, return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl);
  assign return_mult_generic_AC_RND_CONV_false_6_else_2_else_return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl
      = MUX_v_11_2_2(11'b00000000000, return_mult_generic_AC_RND_CONV_false_6_else_2_else_mux_nl,
      return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_or_nl
      = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_6_else_2_else_return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_6_lor_lpi_2_dfm_1);
  assign BUTTERFLY_if_1_and_nl = (~ return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1)
      & out1_rsci_idat_63_0_mx0c1;
  assign BUTTERFLY_if_1_and_1_nl = return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1
      & out1_rsci_idat_63_0_mx0c1;
  assign return_mult_generic_AC_RND_CONV_false_6_oelse_3_not_1_nl = ~ return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1;
  assign return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_and_1_nl
      = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000, (z_out[50:0]),
      return_mult_generic_AC_RND_CONV_false_6_oelse_3_not_1_nl);
  assign stage_PE_index_const_mux_nl = MUX_s_1_2_2(stage_PE_index_const_15_lpi_2_dfm_mx0w0,
      stage_PE_1_index_const_15_lpi_2_dfm, fsm_output[18]);
  assign stage_PE_index_const_mux_3_nl = MUX_s_1_2_2(stage_PE_1_index_const_15_lpi_2_dfm,
      stage_PE_index_const_15_lpi_2_dfm_mx0w0, fsm_output[2]);
  assign stage_PE_index_const_mux_2_nl = MUX_s_1_2_2(stage_PE_index_const_10_lpi_2_dfm_mx0w0,
      stage_PE_1_index_const_10_lpi_2_dfm, fsm_output[18]);
  assign stage_PE_index_const_mux_7_nl = MUX_s_1_2_2(stage_PE_1_index_const_10_lpi_2_dfm,
      stage_PE_index_const_10_lpi_2_dfm_mx0w0, fsm_output[2]);
  assign stage_PE_mux1h_nl = MUX1HOT_s_1_3_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_8,
      t_in_10_0_lpi_1_dfm_1_10, stage_PE_1_index_const_9_1_lpi_2_dfm_8, {or_tmp_180
      , or_tmp_181 , (fsm_output[18])});
  assign stage_PE_mux1h_7_nl = MUX1HOT_s_1_3_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_8,
      t_in_10_0_lpi_1_dfm_1_10, stage_PE_1_index_const_9_1_lpi_2_dfm_8, {or_tmp_180
      , or_tmp_181 , (~ (fsm_output[2]))});
  assign stage_PE_mux1h_1_nl = MUX1HOT_s_1_3_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_7,
      t_in_10_0_lpi_1_dfm_1_9, stage_PE_1_index_const_9_1_lpi_2_dfm_7, {or_tmp_180
      , or_tmp_181 , (fsm_output[18])});
  assign stage_PE_mux1h_9_nl = MUX1HOT_s_1_3_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_7,
      t_in_10_0_lpi_1_dfm_1_9, stage_PE_1_index_const_9_1_lpi_2_dfm_7, {or_tmp_180
      , or_tmp_181 , (~ (fsm_output[2]))});
  assign stage_PE_mux1h_2_nl = MUX1HOT_s_1_3_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_6,
      t_in_10_0_lpi_1_dfm_1_8, stage_PE_1_index_const_9_1_lpi_2_dfm_6, {or_tmp_180
      , or_tmp_181 , (fsm_output[18])});
  assign stage_PE_mux1h_11_nl = MUX1HOT_s_1_3_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_6,
      t_in_10_0_lpi_1_dfm_1_8, stage_PE_1_index_const_9_1_lpi_2_dfm_6, {or_tmp_180
      , or_tmp_181 , (~ (fsm_output[2]))});
  assign BUTTERFLY_i_and_14_nl = (~ mode_lpi_1_dfm) & BUTTERFLY_i_or_4_ssc;
  assign BUTTERFLY_i_or_7_nl = (mode_lpi_1_dfm & BUTTERFLY_i_or_4_ssc) | BUTTERFLY_i_or_5_ssc;
  assign stage_PE_mux1h_3_nl = MUX1HOT_s_1_3_2(stage_PE_asn_13_mx0w0, t_in_10_0_lpi_1_dfm_1_1,
      stage_PE_1_index_const_0_lpi_2_dfm, {or_tmp_180 , or_tmp_181 , (fsm_output[18])});
  assign stage_PE_mux1h_13_nl = MUX1HOT_s_1_3_2(stage_PE_asn_13_mx0w0, t_in_10_0_lpi_1_dfm_1_1,
      stage_PE_1_index_const_0_lpi_2_dfm, {or_tmp_180 , or_tmp_181 , (~ (fsm_output[2]))});
  assign BUTTERFLY_i_mux_1_nl = MUX_v_9_2_2((z_out_49[8:0]), (BUTTERFLY_mux_5_itm_9_0[8:0]),
      or_tmp_46);
  assign t_in_not_nl = ~ nor_155_cse;
  assign stage_PE_stage_PE_stage_PE_mux_3_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_10,
      t_in_10_0_lpi_1_dfm_1_9, operator_11_true_return_26_sva);
  assign BUTTERFLY_if_mux_12_nl = MUX_s_1_2_2(stage_PE_stage_PE_stage_PE_mux_3_nl,
      stage_PE_1_qr_1_10_1_lpi_2_dfm_8, or_tmp_1041);
  assign BUTTERFLY_if_mux_13_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_8, stage_PE_1_qr_1_10_1_lpi_2_dfm_7,
      or_tmp_1041);
  assign BUTTERFLY_if_mux_14_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_7, stage_PE_1_qr_1_10_1_lpi_2_dfm_6,
      or_tmp_1041);
  assign BUTTERFLY_if_mux_15_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_6, stage_PE_1_qr_1_10_1_lpi_2_dfm_5,
      or_tmp_1041);
  assign BUTTERFLY_if_mux_16_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_5, stage_PE_1_qr_1_10_1_lpi_2_dfm_4,
      or_tmp_1041);
  assign BUTTERFLY_if_mux_17_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_4, stage_PE_1_qr_1_10_1_lpi_2_dfm_3,
      or_tmp_1041);
  assign BUTTERFLY_if_mux_18_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_3, stage_PE_1_qr_1_10_1_lpi_2_dfm_2,
      or_tmp_1041);
  assign BUTTERFLY_if_mux_19_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_2, stage_PE_1_qr_1_10_1_lpi_2_dfm_1,
      or_tmp_1041);
  assign BUTTERFLY_if_mux_20_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_1, stage_PE_1_qr_1_10_1_lpi_2_dfm_0,
      or_tmp_1041);
  assign BUTTERFLY_if_mux_21_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_0, stage_PE_1_qr_1_0_lpi_2_dfm,
      or_tmp_1041);
  assign nl_reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_addr_cse  = ({BUTTERFLY_if_mux_12_nl
      , BUTTERFLY_if_mux_13_nl , BUTTERFLY_if_mux_14_nl , BUTTERFLY_if_mux_15_nl
      , BUTTERFLY_if_mux_16_nl , BUTTERFLY_if_mux_17_nl , BUTTERFLY_if_mux_18_nl
      , BUTTERFLY_if_mux_19_nl , BUTTERFLY_if_mux_20_nl , BUTTERFLY_if_mux_21_nl})
      + conv_u2u_9_10(BUTTERFLY_i_div_cmp_z_oreg);
  assign return_add_generic_AC_RND_CONV_false_17_or_nl = (return_add_generic_AC_RND_CONV_false_4_do_sub_sva_1
      & (~ (fsm_output[29]))) | return_add_generic_AC_RND_CONV_false_17_and_3_cse;
  assign return_add_generic_AC_RND_CONV_false_18_return_add_generic_AC_RND_CONV_false_18_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_5_do_sub_sva_1 | (fsm_output[29]));
  assign return_add_generic_AC_RND_CONV_false_18_and_2_nl = return_add_generic_AC_RND_CONV_false_5_do_sub_sva_1
      & (~ (fsm_output[29]));
  assign return_add_generic_AC_RND_CONV_false_18_and_3_nl = (~ nor_99_ssc) & (fsm_output[29]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_3_return_mult_generic_AC_RND_CONV_false_1_if_3_or_1_nl
      = (~ return_mult_generic_AC_RND_CONV_false_1_zero_m_return_mult_generic_AC_RND_CONV_false_1_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_1_r_zero_return_mult_generic_AC_RND_CONV_false_1_r_zero_nor_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_1_lor_lpi_3_dfm_1;
  assign return_mult_generic_AC_RND_CONV_false_2_if_3_return_mult_generic_AC_RND_CONV_false_2_if_3_or_1_nl
      = (~ return_mult_generic_AC_RND_CONV_false_2_zero_m_return_mult_generic_AC_RND_CONV_false_2_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_2_r_zero_return_mult_generic_AC_RND_CONV_false_2_r_zero_nor_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_2_lor_lpi_3_dfm_1;
  assign return_mult_generic_AC_RND_CONV_false_5_if_3_return_mult_generic_AC_RND_CONV_false_5_if_3_or_1_nl
      = (~ return_mult_generic_AC_RND_CONV_false_5_zero_m_return_mult_generic_AC_RND_CONV_false_5_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_5_r_zero_return_mult_generic_AC_RND_CONV_false_5_r_zero_nor_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_5_lor_lpi_3_dfm_1;
  assign return_mult_generic_AC_RND_CONV_false_1_if_not_nl = ~ return_mult_generic_AC_RND_CONV_false_1_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_1_if_nand_1_nl = ~(MUX_v_4_2_2(4'b0000,
      (return_mult_generic_AC_RND_CONV_false_1_exp_acc_tmp[4:1]), return_mult_generic_AC_RND_CONV_false_1_if_not_nl));
  assign return_add_generic_AC_RND_CONV_false_11_mux_23_nl = MUX_s_1_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1,
      (return_add_generic_AC_RND_CONV_false_20_ls_sva[1]), return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1);
  assign not_681_nl = ~ (fsm_output[1]);
  assign stage_PE_qif_qelse_mux_18_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_5, t_in_10_0_lpi_1_dfm_1_4,
      mode_lpi_1_dfm);
  assign stage_PE_qif_qelse_mux_5_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_6, t_in_10_0_lpi_1_dfm_1_5,
      mode_lpi_1_dfm);
  assign stage_PE_qif_qelse_or_nl = (stage_PE_1_and_cse & (fsm_output[2])) | or_tmp_181;
  assign stage_PE_qif_qelse_mux_19_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_6, t_in_10_0_lpi_1_dfm_1_5,
      mode_lpi_1_dfm);
  assign BUTTERFLY_fry_BUTTERFLY_fry_mux_nl = MUX_v_10_2_2(z_out_27, (z_out_55[9:0]),
      fsm_output[37]);
  assign BUTTERFLY_n_BUTTERFLY_n_mux_nl = MUX_v_9_2_2((z_out_49[8:0]), (BUTTERFLY_mux_5_itm_9_0[8:0]),
      fsm_output[34]);
  assign nand_97_nl = ~(and_dcpl_164 & (~ (fsm_output[17])) & (~((fsm_output[4])
      | (fsm_output[18]))) & (~((fsm_output[34]) | (fsm_output[11]))) & (~((fsm_output[12])
      | (fsm_output[16]))) & (~((fsm_output[13]) | (fsm_output[6]) | (fsm_output[10])))
      & (~((fsm_output[7]) | (fsm_output[5]))) & nor_87_cse & nor_88_cse);
  assign BUTTERFLY_n_and_nl = MUX_v_9_2_2(9'b000000000, BUTTERFLY_n_BUTTERFLY_n_mux_nl,
      nand_97_nl);
  assign BUTTERFLY_i_or_2_nl = or_dcpl_325 | BUTTERFLY_1_i_9_0_sva_mx0c3;
  assign return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_3_nl
      = BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx3 | return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp;
  assign return_add_generic_AC_RND_CONV_false_25_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_23_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_23_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_14_op1_mu_and_3_nl = (~ and_255_tmp)
      & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_14_op1_mu_and_4_nl = and_255_tmp &
      (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_1_if_2_return_add_generic_AC_RND_CONV_false_1_if_2_and_2_nl
      = (out_f_d_rsci_q_d[63]) & (stage_PE_1_x_im_d_sva[63]);
  assign return_add_generic_AC_RND_CONV_false_9_if_2_return_add_generic_AC_RND_CONV_false_9_if_2_and_2_nl
      = return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 & (stage_PE_1_x_re_d_sva[63]);
  assign return_add_generic_AC_RND_CONV_false_16_if_2_return_add_generic_AC_RND_CONV_false_16_if_2_nor_1_nl
      = ~((in_f_d_rsci_q_d[63]) | (~ (stage_PE_1_x_im_d_sva[63])));
  assign return_add_generic_AC_RND_CONV_false_13_if_2_return_add_generic_AC_RND_CONV_false_13_if_2_and_2_nl
      = (stage_PE_1_tmp_im_d_1_sva_1_63_51[12]) & (in_f_d_rsci_q_d[63]);
  assign return_add_generic_AC_RND_CONV_false_10_and_2_nl = (~ and_258_tmp) & (fsm_output[6]);
  assign return_add_generic_AC_RND_CONV_false_10_or_5_nl = ((~ return_add_generic_AC_RND_CONV_false_1_op1_smaller_lor_lpi_3_dfm_2)
      & return_add_generic_AC_RND_CONV_false_10_and_3_m1c) | return_add_generic_AC_RND_CONV_false_10_and_18_cse
      | ((~ or_452_cse) & return_add_generic_AC_RND_CONV_false_10_and_9_m1c);
  assign return_add_generic_AC_RND_CONV_false_10_and_15_nl = return_add_generic_AC_RND_CONV_false_1_op1_smaller_lor_lpi_3_dfm_2
      & return_add_generic_AC_RND_CONV_false_10_and_3_m1c;
  assign return_add_generic_AC_RND_CONV_false_10_or_nl = return_add_generic_AC_RND_CONV_false_10_and_4_cse
      | return_add_generic_AC_RND_CONV_false_10_and_12_cse;
  assign return_add_generic_AC_RND_CONV_false_10_or_6_nl = return_add_generic_AC_RND_CONV_false_10_and_16_cse
      | return_add_generic_AC_RND_CONV_false_10_and_24_cse;
  assign return_add_generic_AC_RND_CONV_false_10_or_7_nl = return_add_generic_AC_RND_CONV_false_10_and_17_cse
      | return_add_generic_AC_RND_CONV_false_10_and_25_cse;
  assign return_add_generic_AC_RND_CONV_false_10_and_8_nl = (~ and_261_tmp) & (fsm_output[22]);
  assign return_add_generic_AC_RND_CONV_false_10_and_21_nl = or_452_cse & return_add_generic_AC_RND_CONV_false_10_and_9_m1c;
  assign return_add_generic_AC_RND_CONV_false_10_and_10_nl = (~ and_264_tmp) & (fsm_output[24]);
  assign return_add_generic_AC_RND_CONV_false_10_and_22_nl = (~ or_445_cse) & return_add_generic_AC_RND_CONV_false_10_and_11_m1c;
  assign return_add_generic_AC_RND_CONV_false_10_and_23_nl = or_445_cse & return_add_generic_AC_RND_CONV_false_10_and_11_m1c;
  assign return_extract_17_m_zero_return_extract_17_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_1
      | (return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_47_m_zero_return_extract_47_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm
      | (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_mx0w5!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_59_m_zero_return_extract_59_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm_mx2
      | (return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_mx0w6!=51'b000000000000000000000000000000000000000000000000000));
  assign or_916_nl = (fsm_output[28]) | (fsm_output[10]);
  assign return_extract_45_m_zero_return_extract_45_m_zero_nor_nl = ~(stage_PE_1_tmp_im_d_1_lpi_3_dfm_51_mx1
      | (stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_44_m_zero_return_extract_44_m_zero_nor_nl = ~(stage_PE_1_tmp_re_d_1_lpi_3_dfm_51_mx1
      | stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx2_50 | (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1[49:0]!=50'b00000000000000000000000000000000000000000000000000));
  assign return_extract_52_m_zero_return_extract_52_m_zero_nor_nl = ~(BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx3
      | (return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_57_m_zero_return_extract_57_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_17_m_zero_or_1_nl = (fsm_output[5]) | (fsm_output[8]);
  assign operator_11_true_12_operator_11_true_12_and_nl = (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_1==10'b1111111111)
      & stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0;
  assign operator_11_true_20_operator_11_true_20_and_nl = (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1==11'b11111111111);
  assign operator_11_true_25_operator_11_true_25_and_nl = (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1;
  assign operator_11_true_45_operator_11_true_45_and_nl = (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_1==10'b1111111111)
      & stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0;
  assign operator_11_true_44_operator_11_true_44_and_nl = (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx1_10_1==10'b1111111111)
      & stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx1_0;
  assign operator_11_true_52_operator_11_true_52_and_nl = (return_mult_generic_AC_RND_CONV_false_3_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w7==11'b11111111111);
  assign operator_11_true_57_operator_11_true_57_and_nl = (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1;
  assign or_934_nl = (fsm_output[24]) | (fsm_output[21]);
  assign BUTTERFLY_and_5_nl = (~ inverse_lpi_1_dfm_1) & (fsm_output[6]);
  assign BUTTERFLY_and_6_nl = inverse_lpi_1_dfm_1 & (fsm_output[6]);
  assign return_add_generic_AC_RND_CONV_false_24_if_7_return_add_generic_AC_RND_CONV_false_24_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_24_exception_sva_1 | leading_sign_57_0_1_0_24_out_2);
  assign return_add_generic_AC_RND_CONV_false_24_return_add_generic_AC_RND_CONV_false_24_and_4_nl
      = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000, (return_add_generic_AC_RND_CONV_false_24_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_24_if_7_return_add_generic_AC_RND_CONV_false_24_if_7_nor_nl);
  assign or_939_nl = (inverse_lpi_1_dfm_1 & return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp
      & (fsm_output[7])) | (return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp
      & (fsm_output[5]));
  assign or_940_nl = (inverse_lpi_1_dfm_1 & (~ return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp)
      & (fsm_output[7])) | ((~ return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp)
      & (fsm_output[5]));
  assign and_990_nl = return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp
      & or_dcpl_385;
  assign and_992_nl = (~ return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp)
      & or_dcpl_385;
  assign return_add_generic_AC_RND_CONV_false_17_or_4_nl = return_add_generic_AC_RND_CONV_false_17_and_7_cse
      | return_add_generic_AC_RND_CONV_false_17_and_9_cse;
  assign return_add_generic_AC_RND_CONV_false_17_or_5_nl = return_add_generic_AC_RND_CONV_false_17_and_8_cse
      | return_add_generic_AC_RND_CONV_false_17_and_3_cse;
  assign return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_3_nl
      = return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2 | return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_tmp;
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_nl = (~ return_add_generic_AC_RND_CONV_false_10_do_sub_sva)
      & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_nl = return_add_generic_AC_RND_CONV_false_10_do_sub_sva
      & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_nl = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse;
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_17_nl = MUX1HOT_v_56_4_2((~
      (z_out_30[56:1])), (z_out_30[56:1]), (z_out_29[56:1]), (~ (z_out_29[56:1])),
      {return_add_generic_AC_RND_CONV_false_3_or_4_cse , return_add_generic_AC_RND_CONV_false_3_or_5_cse
      , return_add_generic_AC_RND_CONV_false_3_and_8_cse , return_add_generic_AC_RND_CONV_false_3_and_9_cse});
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_18_nl = MUX1HOT_s_1_10_2((~
      return_add_generic_AC_RND_CONV_false_3_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_3_res_mant_3_0_sva_1,
      return_add_generic_AC_RND_CONV_false_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_res_mant_3_0_sva_1),
      (~ return_add_generic_AC_RND_CONV_false_16_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_16_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_15_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_15_res_mant_3_0_sva_1,
      return_add_generic_AC_RND_CONV_false_23_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_23_res_mant_3_0_sva_1),
      {return_add_generic_AC_RND_CONV_false_3_and_cse , return_add_generic_AC_RND_CONV_false_3_and_1_cse
      , return_add_generic_AC_RND_CONV_false_3_and_2_cse , return_add_generic_AC_RND_CONV_false_3_and_3_cse
      , return_add_generic_AC_RND_CONV_false_3_and_4_cse , return_add_generic_AC_RND_CONV_false_3_and_5_cse
      , return_add_generic_AC_RND_CONV_false_3_and_6_cse , return_add_generic_AC_RND_CONV_false_3_and_7_cse
      , return_add_generic_AC_RND_CONV_false_3_and_8_cse , return_add_generic_AC_RND_CONV_false_3_and_9_cse});
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_19_nl = MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_3_do_sub_sva_1,
      return_add_generic_AC_RND_CONV_false_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_16_do_sub_sva_1,
      return_add_generic_AC_RND_CONV_false_15_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_10_op2_inf_sva,
      {(fsm_output[6]) , (fsm_output[8]) , (fsm_output[22]) , (fsm_output[24]) ,
      (fsm_output[29])});
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_20_nl = MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_3_op_bigger_mux_1_cse,
      return_add_generic_AC_RND_CONV_false_op_bigger_mux_1_cse, return_add_generic_AC_RND_CONV_false_16_op_bigger_mux_1_cse,
      return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_1_cse, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0, {(fsm_output[6])
      , (fsm_output[8]) , (fsm_output[22]) , (fsm_output[24]) , return_add_generic_AC_RND_CONV_false_3_and_20_cse
      , and_1813_cse});
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_21_nl = MUX1HOT_s_1_6_2((return_add_generic_AC_RND_CONV_false_3_op_bigger_mux_2_cse[50]),
      (return_add_generic_AC_RND_CONV_false_op_bigger_mux_2_cse[50]), (return_add_generic_AC_RND_CONV_false_16_op_bigger_mux_2_cse[50]),
      (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_cse[50]), (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[50]),
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0, {(fsm_output[6])
      , (fsm_output[8]) , (fsm_output[22]) , (fsm_output[24]) , return_add_generic_AC_RND_CONV_false_3_and_20_cse
      , and_1813_cse});
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_22_nl = MUX1HOT_v_50_6_2((return_add_generic_AC_RND_CONV_false_3_op_bigger_mux_2_cse[49:0]),
      (return_add_generic_AC_RND_CONV_false_op_bigger_mux_2_cse[49:0]), (return_add_generic_AC_RND_CONV_false_16_op_bigger_mux_2_cse[49:0]),
      (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_cse[49:0]), (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[49:0]),
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0, {(fsm_output[6])
      , (fsm_output[8]) , (fsm_output[22]) , (fsm_output[24]) , return_add_generic_AC_RND_CONV_false_3_and_20_cse
      , and_1813_cse});
  assign return_add_generic_AC_RND_CONV_false_3_or_17_nl = return_add_generic_AC_RND_CONV_false_3_and_30_cse
      | return_add_generic_AC_RND_CONV_false_3_and_32_cse | return_add_generic_AC_RND_CONV_false_3_and_20_cse;
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_23_nl = MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1,
      {return_add_generic_AC_RND_CONV_false_3_or_17_nl , return_add_generic_AC_RND_CONV_false_3_or_14_cse
      , or_956_cse , return_add_generic_AC_RND_CONV_false_3_or_16_cse , and_1813_cse});
  assign nl_acc_4_nl = ({return_add_generic_AC_RND_CONV_false_3_mux1h_17_nl , return_add_generic_AC_RND_CONV_false_3_mux1h_18_nl
      , return_add_generic_AC_RND_CONV_false_3_mux1h_19_nl}) + conv_u2u_57_58({return_add_generic_AC_RND_CONV_false_3_mux1h_20_nl
      , return_add_generic_AC_RND_CONV_false_3_mux1h_21_nl , return_add_generic_AC_RND_CONV_false_3_mux1h_22_nl
      , return_add_generic_AC_RND_CONV_false_3_mux1h_23_nl , 4'b0001});
  assign acc_4_nl = nl_acc_4_nl[57:0];
  assign return_add_generic_AC_RND_CONV_false_15_res_mant_or_4_nl = return_add_generic_AC_RND_CONV_false_15_res_mant_or_cse
      | (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_15_res_mant_or_5_nl = (fsm_output[14])
      | return_add_generic_AC_RND_CONV_false_15_res_mant_or_1_cse;
  assign return_add_generic_AC_RND_CONV_false_10_do_sub_return_add_generic_AC_RND_CONV_false_10_do_sub_xor_nl
      = (stage_PE_1_x_im_d_sva[63]) ^ operator_11_true_return_15_sva_mx1;
  assign return_add_generic_AC_RND_CONV_false_19_do_sub_return_add_generic_AC_RND_CONV_false_19_do_sub_return_add_generic_AC_RND_CONV_false_19_do_sub_xnor_nl
      = ~(stage_PE_1_tmp_re_d_1_lpi_3_dfm_63_mx1 ^ stage_PE_1_tmp_im_d_1_lpi_3_dfm_63);
  assign return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_xnor_nl
      = ~((stage_PE_1_x_im_d_sva[63]) ^ operator_11_true_return_15_sva_mx2);
  assign return_add_generic_AC_RND_CONV_false_4_if_2_return_add_generic_AC_RND_CONV_false_4_if_2_nor_1_nl
      = ~(inverse_lpi_1_dfm_1 | (~ (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[63])));
  assign return_add_generic_AC_RND_CONV_false_4_r_sign_mux_1_nl = MUX_s_1_2_2((BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[63]),
      (~ inverse_lpi_1_dfm_1), return_add_generic_AC_RND_CONV_false_17_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_4_if_2_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_4_if_2_return_add_generic_AC_RND_CONV_false_4_if_2_nor_1_nl,
      return_add_generic_AC_RND_CONV_false_4_r_sign_mux_1_nl, or_dcpl_474);
  assign return_add_generic_AC_RND_CONV_false_25_r_sign_mux_1_nl = MUX_s_1_2_2((stage_PE_1_x_im_d_sva[63]),
      (~ operator_11_true_return_15_sva), return_add_generic_AC_RND_CONV_false_25_op1_smaller_return_add_generic_AC_RND_CONV_false_25_op1_smaller_or_cse);
  assign return_add_generic_AC_RND_CONV_false_12_if_2_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_12_if_2_return_add_generic_AC_RND_CONV_false_12_if_2_nor_mx3w0,
      return_add_generic_AC_RND_CONV_false_25_r_sign_mux_1_nl, or_dcpl_480);
  assign return_add_generic_AC_RND_CONV_false_5_if_2_return_add_generic_AC_RND_CONV_false_5_if_2_and_2_nl
      = inverse_lpi_1_dfm_1 & (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[63]);
  assign return_add_generic_AC_RND_CONV_false_5_r_sign_mux_1_nl = MUX_s_1_2_2((BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[63]),
      inverse_lpi_1_dfm_1, return_add_generic_AC_RND_CONV_false_17_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_3_if_2_return_add_generic_AC_RND_CONV_false_3_if_2_nor_1_nl
      = ~((out_f_d_rsci_q_d[63]) | (~ (stage_PE_1_x_im_d_sva[63])));
  assign return_add_generic_AC_RND_CONV_false_2_if_2_return_add_generic_AC_RND_CONV_false_2_if_2_nor_1_nl
      = ~((stage_PE_1_tmp_im_d_1_sva_1_63_51[12]) | (~ (out_f_d_rsci_q_d[63])));
  assign return_add_generic_AC_RND_CONV_false_14_if_2_return_add_generic_AC_RND_CONV_false_14_if_2_and_2_nl
      = (in_f_d_rsci_q_d[63]) & (stage_PE_1_x_im_d_sva[63]);
  assign return_add_generic_AC_RND_CONV_false_11_and_25_nl = (~ or_dcpl_356) & (fsm_output[6]);
  assign return_add_generic_AC_RND_CONV_false_11_or_4_nl = ((~ return_add_generic_AC_RND_CONV_false_1_op1_smaller_lor_lpi_3_dfm_2)
      & return_add_generic_AC_RND_CONV_false_11_and_26_m1c) | ((~ or_452_cse) & return_add_generic_AC_RND_CONV_false_11_and_32_m1c)
      | ((~ return_add_generic_AC_RND_CONV_false_25_op1_smaller_return_add_generic_AC_RND_CONV_false_25_op1_smaller_or_cse)
      & return_add_generic_AC_RND_CONV_false_11_and_34_m1c);
  assign return_add_generic_AC_RND_CONV_false_11_and_36_nl = return_add_generic_AC_RND_CONV_false_1_op1_smaller_lor_lpi_3_dfm_2
      & return_add_generic_AC_RND_CONV_false_11_and_26_m1c;
  assign return_add_generic_AC_RND_CONV_false_11_and_31_nl = (~ or_dcpl_359) & (fsm_output[22]);
  assign return_add_generic_AC_RND_CONV_false_11_and_42_nl = or_452_cse & return_add_generic_AC_RND_CONV_false_11_and_32_m1c;
  assign return_add_generic_AC_RND_CONV_false_11_and_33_nl = (~ or_dcpl_480) & (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_11_and_44_nl = return_add_generic_AC_RND_CONV_false_25_op1_smaller_return_add_generic_AC_RND_CONV_false_25_op1_smaller_or_cse
      & return_add_generic_AC_RND_CONV_false_11_and_34_m1c;
  assign return_add_generic_AC_RND_CONV_false_if_2_return_add_generic_AC_RND_CONV_false_if_2_and_2_nl
      = (stage_PE_1_tmp_im_d_1_sva_1_63_51[12]) & (out_f_d_rsci_q_d[63]);
  assign return_add_generic_AC_RND_CONV_false_7_do_sub_return_add_generic_AC_RND_CONV_false_7_do_sub_xor_nl
      = stage_d_mul_return_d_63_sva_1 ^ stage_d_mul_return_d_2_63_sva_1;
  assign return_add_generic_AC_RND_CONV_false_15_if_2_return_add_generic_AC_RND_CONV_false_15_if_2_nor_1_nl
      = ~((stage_PE_1_tmp_im_d_1_sva_1_63_51[12]) | (~ (in_f_d_rsci_q_d[63])));
  assign return_add_generic_AC_RND_CONV_false_20_do_sub_return_add_generic_AC_RND_CONV_false_20_do_sub_xor_nl
      = stage_d_mul_return_d_63_sva_1 ^ stage_d_mul_return_d_5_63_sva_1;
  assign return_add_generic_AC_RND_CONV_false_12_and_5_nl = (~ or_dcpl_360) & (fsm_output[24]);
  assign return_add_generic_AC_RND_CONV_false_12_and_13_nl = (~ or_445_cse) & return_add_generic_AC_RND_CONV_false_12_and_6_m1c;
  assign return_add_generic_AC_RND_CONV_false_12_and_14_nl = or_445_cse & return_add_generic_AC_RND_CONV_false_12_and_6_m1c;
  assign return_extract_50_and_nl = return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_if_1_return_add_generic_AC_RND_CONV_false_17_op2_normal_return_extract_41_nor_tmp
      & (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[51:0]==52'b0000000000000000000000000000000000000000000000000000);
  assign return_extract_15_m_zero_return_extract_15_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_4_m_r_51_lpi_3_dfm_1
      | (return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_mx0w2!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_27_m_zero_return_extract_27_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm_mx1
      | (return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_mx0w4!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_17_m_zero_or_2_nl = (fsm_output[21]) | (fsm_output[23]);
  assign operator_11_true_13_operator_11_true_13_and_nl = (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_1==10'b1111111111)
      & stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0;
  assign operator_11_true_53_operator_11_true_53_and_nl = (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1==11'b11111111111);
  assign operator_11_true_27_operator_11_true_27_and_nl = (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_mx0w2==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1;
  assign operator_11_true_59_operator_11_true_59_and_nl = (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_mx1w0==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_6_do_sub_return_add_generic_AC_RND_CONV_false_6_do_sub_return_add_generic_AC_RND_CONV_false_6_do_sub_xnor_nl
      = ~(return_add_generic_AC_RND_CONV_false_11_mux_19_cse ^ stage_PE_1_tmp_im_d_1_lpi_3_dfm_63);
  assign return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_xnor_nl
      = ~((stage_PE_1_x_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1);
  assign return_add_generic_AC_RND_CONV_false_21_do_sub_return_add_generic_AC_RND_CONV_false_21_do_sub_xor_nl
      = stage_d_mul_return_d_1_63_sva_1 ^ stage_d_mul_return_d_5_63_sva_1;
  assign return_add_generic_AC_RND_CONV_false_8_do_sub_return_add_generic_AC_RND_CONV_false_8_do_sub_xor_nl
      = stage_d_mul_return_d_1_63_sva_1 ^ stage_d_mul_return_d_2_63_sva_1;
  assign return_add_generic_AC_RND_CONV_false_22_do_sub_return_add_generic_AC_RND_CONV_false_22_do_sub_xor_nl
      = (stage_PE_1_x_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2;
  assign return_add_generic_AC_RND_CONV_false_14_mux1h_8_nl = MUX1HOT_v_51_6_2(return_add_generic_AC_RND_CONV_false_4_op2_mu_51_1_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_4_op1_mu_51_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_1_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1, return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1,
      (return_add_generic_AC_RND_CONV_false_23_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      {return_add_generic_AC_RND_CONV_false_11_op_bigger_and_4_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_5_cse
      , return_add_generic_AC_RND_CONV_false_14_or_cse , (fsm_output[10]) , (fsm_output[26])
      , (fsm_output[30])});
  assign nor_157_nl = ~(((return_add_generic_AC_RND_CONV_false_14_exception_sva_1
      | leading_sign_57_0_1_0_2_out_2) & (fsm_output[23])) | ((return_add_generic_AC_RND_CONV_false_1_exception_sva_1
      | leading_sign_57_0_1_0_2_out_2) & (fsm_output[7])) | ((leading_sign_57_0_1_0_15_out_2
      | return_add_generic_AC_RND_CONV_false_23_exception_sva_1) & (fsm_output[30])));
  assign stage_PE_1_tmp_im_d_and_5_nl = (~ inverse_lpi_1_dfm_1) & (fsm_output[23]);
  assign stage_PE_1_x_im_d_and_1_nl = (~ or_tmp_773) & return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_2_cse;
  assign mux1h_nl = MUX1HOT_v_4_11_2((r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[61:58]),
      (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[61:58]), (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1[9:6]),
      (stage_PE_1_x_re_d_sva[62:59]), in_u_rsc_merge_sva_rsp_1_rsp_0, (stage_PE_1_x_im_d_sva[62:59]),
      (z_out_12[9:6]), (operator_33_true_34_acc_psp_1_sva_1[10:7]), (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1[9:6]),
      (return_add_generic_AC_RND_CONV_false_24_exp_plus_1_12_1_lpi_3_dfm_1[9:6]),
      (operator_33_true_48_acc_tmp[10:7]), {and_2120_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_5_cse
      , and_1132_ssc , and_2123_cse , and_1804_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_11_cse
      , and_2126_cse , and_2127_cse , and_1145_ssc , and_2129_cse , and_2130_cse});
  assign not_730_nl = ~ or_dcpl_629;
  assign and_2119_nl = MUX_v_4_2_2(4'b0000, mux1h_nl, not_730_nl);
  assign mux1h_2_nl = MUX1HOT_v_6_11_2((r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[57:52]),
      (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[57:52]), (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1[5:0]),
      (stage_PE_1_x_re_d_sva[58:53]), in_u_rsc_merge_sva_rsp_1_rsp_1, (stage_PE_1_x_im_d_sva[58:53]),
      (z_out_12[5:0]), (operator_33_true_34_acc_psp_1_sva_1[6:1]), (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1[5:0]),
      (return_add_generic_AC_RND_CONV_false_24_exp_plus_1_12_1_lpi_3_dfm_1[5:0]),
      (operator_33_true_48_acc_tmp[6:1]), {and_2120_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_5_cse
      , and_1132_ssc , and_2123_cse , and_1804_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_11_cse
      , and_2126_cse , and_2127_cse , and_1145_ssc , and_2129_cse , and_2130_cse});
  assign not_732_nl = ~ or_dcpl_629;
  assign and_2131_nl = MUX_v_6_2_2(6'b000000, mux1h_2_nl, not_732_nl);
  assign and_2628_nl = (fsm_output[12]) & return_add_generic_AC_RND_CONV_false_7_op1_smaller_lor_lpi_3_dfm_2;
  assign mux_20_nl = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp[11]),
      return_add_generic_AC_RND_CONV_false_7_op1_smaller_lor_lpi_3_dfm_2, fsm_output[12]);
  assign or_1755_nl = (return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp[11])
      | return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp;
  assign mux_21_nl = MUX_s_1_2_2(mux_20_nl, or_1755_nl, return_add_generic_AC_RND_CONV_false_21_ma1_lt_ma2_acc_1_itm_52);
  assign mux_22_nl = MUX_s_1_2_2(and_2628_nl, mux_21_nl, fsm_output[28]);
  assign BUTTERFLY_else_2_and_8_nl = or_959_rgt & (~ BUTTERFLY_else_2_and_2_rgt);
  assign return_add_generic_AC_RND_CONV_false_25_if_7_return_add_generic_AC_RND_CONV_false_25_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_25_exception_sva_1 | leading_sign_57_0_1_0_25_out_2);
  assign return_add_generic_AC_RND_CONV_false_25_return_add_generic_AC_RND_CONV_false_25_and_4_nl
      = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000, (return_add_generic_AC_RND_CONV_false_25_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_25_if_7_return_add_generic_AC_RND_CONV_false_25_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_18_and_15_nl = (fsm_output[29]) & (or_dcpl_477
      | or_dcpl_387 | or_dcpl_300 | return_add_generic_AC_RND_CONV_false_18_and_8_cse);
  assign and_304_nl = (~ inverse_lpi_1_dfm_1) & return_add_generic_AC_RND_CONV_false_10_do_sub_sva
      & (fsm_output[29]);
  assign return_extract_54_m_zero_return_extract_54_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx6
      | (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_add_generic_AC_RND_CONV_false_19_op2_mu_and_2_nl = (~ return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_1_return_add_generic_AC_RND_CONV_false_6_op2_normal_return_extract_13_nor_tmp)
      & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_19_op2_mu_and_3_nl = return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_1_return_add_generic_AC_RND_CONV_false_6_op2_normal_return_extract_13_nor_tmp
      & (fsm_output[7]);
  assign or_1195_nl = (fsm_output[32]) | (fsm_output[16]) | (fsm_output[13]) | return_add_generic_AC_RND_CONV_false_18_and_8_cse;
  assign BUTTERFLY_1_fiy_and_1_nl = (~ return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1)
      & (fsm_output[15]);
  assign BUTTERFLY_1_fiy_and_2_nl = return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1
      & (fsm_output[15]);
  assign return_add_generic_AC_RND_CONV_false_1_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_14_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_14_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_13_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_14_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_14_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_14_op1_inf_sva_1
      & return_mult_generic_AC_RND_CONV_false_op1_zero_sva_1 & return_add_generic_AC_RND_CONV_false_13_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_23_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_23_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_23_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva);
  assign return_add_generic_AC_RND_CONV_false_9_exp_and_1_nl = (~ and_336_cse) &
      (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_9_exp_or_nl = (and_336_cse & (fsm_output[7]))
      | (and_336_cse & (fsm_output[23]));
  assign return_add_generic_AC_RND_CONV_false_9_exp_and_5_nl = (~ and_336_cse) &
      (fsm_output[23]);
  assign return_add_generic_AC_RND_CONV_false_9_exp_and_7_nl = (~ and_dcpl_241) &
      (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_9_exp_and_9_nl = (~ and_342_tmp) &
      (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_9_exp_and_10_nl = and_342_tmp & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_25_e_r_qelse_not_2_nl = ~ return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs;
  assign return_add_generic_AC_RND_CONV_false_25_e_r_qelse_return_add_generic_AC_RND_CONV_false_25_e_r_qelse_and_nl
      = MUX_v_10_2_2(10'b0000000000, ({reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0
      , reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1}), return_add_generic_AC_RND_CONV_false_25_e_r_qelse_not_2_nl);
  assign return_add_generic_AC_RND_CONV_false_14_e_r_mux1h_6_nl = MUX1HOT_v_10_5_2(return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_mx1w0, return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1,
      (stage_PE_1_x_re_d_sva[62:53]), return_add_generic_AC_RND_CONV_false_25_e_r_qelse_return_add_generic_AC_RND_CONV_false_25_e_r_qelse_and_nl,
      {(fsm_output[13]) , return_add_generic_AC_RND_CONV_false_18_and_8_cse , BUTTERFLY_1_fiy_and_4_cse
      , BUTTERFLY_1_fiy_and_5_cse , (fsm_output[31])});
  assign return_add_generic_AC_RND_CONV_false_14_e_r_nor_2_nl = ~((fsm_output[7])
      | (fsm_output[23]));
  assign return_add_generic_AC_RND_CONV_false_14_e_r_and_5_nl = MUX_v_10_2_2(10'b0000000000,
      return_add_generic_AC_RND_CONV_false_14_e_r_mux1h_6_nl, return_add_generic_AC_RND_CONV_false_14_e_r_nor_2_nl);
  assign or_1771_nl = ((~ return_add_generic_AC_RND_CONV_false_14_exception_sva_1)
      & (fsm_output[23])) | ((~ return_add_generic_AC_RND_CONV_false_1_exception_sva_1)
      & (fsm_output[7]));
  assign mux_25_nl = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_14_e_r_and_5_nl,
      return_add_generic_AC_RND_CONV_false_1_e_r_qelse_qr_10_1_lpi_3_dfm_1, or_1771_nl);
  assign or_1772_nl = (return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva & (fsm_output[31]))
      | (return_add_generic_AC_RND_CONV_false_14_exception_sva_1 & (fsm_output[23]))
      | (return_add_generic_AC_RND_CONV_false_1_exception_sva_1 & (fsm_output[7]));
  assign return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs, or_dcpl_159);
  assign return_add_generic_AC_RND_CONV_false_1_e_r_return_add_generic_AC_RND_CONV_false_1_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_32 & (~ return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_1_nl))
      | return_add_generic_AC_RND_CONV_false_1_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_5_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs, or_dcpl_159);
  assign return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_32 & (~ return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_5_nl))
      | return_add_generic_AC_RND_CONV_false_14_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_25_return_add_generic_AC_RND_CONV_false_25_and_5_nl
      = (operator_33_true_50_acc_tmp[0]) & return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11;
  assign return_add_generic_AC_RND_CONV_false_25_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_25_return_add_generic_AC_RND_CONV_false_25_and_5_nl,
      return_add_generic_AC_RND_CONV_false_25_exp_plus_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_25_res_rounded_acc_tmp[53]);
  assign or_312_nl = or_dcpl_250 | and_dcpl_141 | return_add_generic_AC_RND_CONV_false_25_r_inf_lpi_3_dfm_2;
  assign return_add_generic_AC_RND_CONV_false_25_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs, or_312_nl);
  assign return_add_generic_AC_RND_CONV_false_25_e_r_qelse_return_add_generic_AC_RND_CONV_false_25_e_r_qelse_and_1_nl
      = return_add_generic_AC_RND_CONV_false_25_mux_13_nl & (~ return_add_generic_AC_RND_CONV_false_25_e_r_qelse_mux_1_nl);
  assign return_extract_13_m_zero_return_extract_13_m_zero_nor_nl = ~(stage_PE_tmp_im_d_1_lpi_3_dfm_51_mx0
      | (stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_12_m_zero_return_extract_12_m_zero_nor_nl = ~(stage_PE_tmp_re_d_1_lpi_3_dfm_51_mx0
      | stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx1_50 | (stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0[49:0]!=50'b00000000000000000000000000000000000000000000000000));
  assign return_extract_20_m_zero_return_extract_20_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2
      | (return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_25_m_zero_return_extract_25_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign operator_11_true_17_operator_11_true_17_and_nl = (return_add_generic_AC_RND_CONV_false_5_e_r_qelse_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1;
  assign operator_11_true_22_operator_11_true_22_and_nl = (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w3==11'b11111111111);
  assign operator_11_true_54_operator_11_true_54_and_nl = (return_mult_generic_AC_RND_CONV_false_4_exp_1_11_0_lpi_3_dfm_3_10_0_1==11'b11111111111);
  assign return_extract_15_return_extract_15_nor_nl = ~((return_add_generic_AC_RND_CONV_false_4_e_r_qelse_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1);
  assign return_extract_47_return_extract_47_nor_nl = ~((return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_mx0w4_9_6!=4'b0000)
      | (return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_mx0w4_5_0!=6'b000000)
      | return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_and_1_itm);
  assign return_add_generic_AC_RND_CONV_false_19_op2_mu_return_add_generic_AC_RND_CONV_false_19_op2_mu_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_cse_sva
      | (fsm_output[13]));
  assign return_add_generic_AC_RND_CONV_false_19_op2_mu_and_5_nl = return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_cse_sva
      & (~ (fsm_output[13]));
  assign operator_11_true_15_operator_11_true_15_and_nl = (return_add_generic_AC_RND_CONV_false_4_e_r_qelse_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1;
  assign operator_11_true_47_operator_11_true_47_and_nl = (return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_mx0w4_9_6==4'b1111)
      & (return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_mx0w4_5_0==6'b111111)
      & return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_and_1_itm;
  assign return_extract_15_return_extract_15_or_1_nl = (return_add_generic_AC_RND_CONV_false_4_e_r_qelse_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1;
  assign return_extract_47_return_extract_47_or_1_nl = (return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_mx0w4_9_6!=4'b0000)
      | (return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_mx0w4_5_0!=6'b000000)
      | return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_and_1_itm;
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_or_nl = (z_out_54[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_or_2
      & (z_out_54[51]));
  assign return_mult_generic_AC_RND_CONV_false_1_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_1_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_1_else_1_sticky_bit_or_nl
      = ((z_out_26[105]) & (~ (z_out_38[52]))) | ((z_out_26[104]) & (~ (z_out_38[51])))
      | ((z_out_26[103]) & (~ (z_out_38[50]))) | ((z_out_26[102]) & (~ (z_out_38[49])))
      | ((z_out_26[101]) & (~ (z_out_38[48]))) | ((z_out_26[100]) & (~ (z_out_38[47])))
      | ((z_out_26[99]) & (~ (z_out_38[46]))) | ((z_out_26[98]) & (~ (z_out_38[45])))
      | ((z_out_26[97]) & (~ (z_out_38[44]))) | ((z_out_26[96]) & (~ (z_out_38[43])))
      | ((z_out_26[95]) & (~ (z_out_38[42]))) | ((z_out_26[94]) & (~ (z_out_38[41])))
      | ((z_out_26[93]) & (~ (z_out_38[40]))) | ((z_out_26[92]) & (~ (z_out_38[39])))
      | ((z_out_26[91]) & (~ (z_out_38[38]))) | ((z_out_26[90]) & (~ (z_out_38[37])))
      | ((z_out_26[89]) & (~ (z_out_38[36]))) | ((z_out_26[88]) & (~ (z_out_38[35])))
      | ((z_out_26[87]) & (~ (z_out_38[34]))) | ((z_out_26[86]) & (~ (z_out_38[33])))
      | ((z_out_26[85]) & (~ (z_out_38[32]))) | ((z_out_26[84]) & (~ (z_out_38[31])))
      | ((z_out_26[83]) & (~ (z_out_38[30]))) | ((z_out_26[82]) & (~ (z_out_38[29])))
      | ((z_out_26[81]) & (~ (z_out_38[28]))) | ((z_out_26[80]) & (~ (z_out_38[27])))
      | ((z_out_26[79]) & (~ (z_out_38[26]))) | ((z_out_26[78]) & (~ (z_out_38[25])))
      | ((z_out_26[77]) & (~ (z_out_38[24]))) | ((z_out_26[76]) & (~ (z_out_38[23])))
      | ((z_out_26[75]) & (~ (z_out_38[22]))) | ((z_out_26[74]) & (~ (z_out_38[21])))
      | ((z_out_26[73]) & (~ (z_out_38[20]))) | ((z_out_26[72]) & (~ (z_out_38[19])))
      | ((z_out_26[71]) & (~ (z_out_38[18]))) | ((z_out_26[70]) & (~ (z_out_38[17])))
      | ((z_out_26[69]) & (~ (z_out_38[16]))) | ((z_out_26[68]) & (~ (z_out_38[15])))
      | ((z_out_26[67]) & (~ (z_out_38[14]))) | ((z_out_26[66]) & (~ (z_out_38[13])))
      | ((z_out_26[65]) & (~ (z_out_38[12]))) | ((z_out_26[64]) & (~ (z_out_38[11])))
      | ((z_out_26[63]) & (~ (z_out_38[10]))) | ((z_out_26[62]) & (~ (z_out_38[9])))
      | ((z_out_26[61]) & (~ (z_out_38[8]))) | ((z_out_26[60]) & (~ (z_out_38[7])))
      | ((z_out_26[59]) & (~ (z_out_38[6]))) | ((z_out_26[58]) & (~ (z_out_38[5])))
      | ((z_out_26[57]) & (~ (z_out_38[4]))) | ((z_out_26[56]) & (~ (z_out_38[3])))
      | ((z_out_26[55]) & (~ (z_out_38[2]))) | ((z_out_26[54]) & (~ (z_out_38[1])))
      | ((z_out_26[53]) & (~ (z_out_38[0]))) | (z_out_26[52:0]!=53'b00000000000000000000000000000000000000000000000000000);
  assign return_mult_generic_AC_RND_CONV_false_1_mux_13_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_1_if_1_or_nl,
      return_mult_generic_AC_RND_CONV_false_1_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_1_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_1_else_1_sticky_bit_or_nl,
      stage_u_add_3_acc_itm_rsp_1[12]);
  assign return_mult_generic_AC_RND_CONV_false_1_or_nl = return_mult_generic_AC_RND_CONV_false_1_mux_13_nl
      | (z_out_53[1]);
  assign return_mult_generic_AC_RND_CONV_false_2_if_1_or_nl = (return_mult_generic_AC_RND_CONV_false_2_p_sva_1[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_or_2
      & (return_mult_generic_AC_RND_CONV_false_2_p_sva_1[51]));
  assign return_mult_generic_AC_RND_CONV_false_2_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_2_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_2_else_1_sticky_bit_or_nl
      = ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[105]) & (~ (z_out_38[52])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[104]) & (~ (z_out_38[51])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[103]) & (~ (z_out_38[50])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[102]) & (~ (z_out_38[49])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[101]) & (~ (z_out_38[48])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[100]) & (~ (z_out_38[47])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[99]) & (~ (z_out_38[46])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[98]) & (~ (z_out_38[45])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[97]) & (~ (z_out_38[44])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[96]) & (~ (z_out_38[43])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[95]) & (~ (z_out_38[42])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[94]) & (~ (z_out_38[41])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[93]) & (~ (z_out_38[40])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[92]) & (~ (z_out_38[39])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[91]) & (~ (z_out_38[38])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[90]) & (~ (z_out_38[37])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[89]) & (~ (z_out_38[36])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[88]) & (~ (z_out_38[35])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[87]) & (~ (z_out_38[34])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[86]) & (~ (z_out_38[33])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[85]) & (~ (z_out_38[32])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[84]) & (~ (z_out_38[31])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[83]) & (~ (z_out_38[30])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[82]) & (~ (z_out_38[29])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[81]) & (~ (z_out_38[28])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[80]) & (~ (z_out_38[27])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[79]) & (~ (z_out_38[26])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[78]) & (~ (z_out_38[25])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[77]) & (~ (z_out_38[24])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[76]) & (~ (z_out_38[23])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[75]) & (~ (z_out_38[22])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[74]) & (~ (z_out_38[21])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[73]) & (~ (z_out_38[20])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[72]) & (~ (z_out_38[19])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[71]) & (~ (z_out_38[18])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[70]) & (~ (z_out_38[17])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[69]) & (~ (z_out_38[16])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[68]) & (~ (z_out_38[15])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[67]) & (~ (z_out_38[14])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[66]) & (~ (z_out_38[13])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[65]) & (~ (z_out_38[12])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[64]) & (~ (z_out_38[11])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[63]) & (~ (z_out_38[10])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[62]) & (~ (z_out_38[9])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[61]) & (~ (z_out_38[8])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[60]) & (~ (z_out_38[7])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[59]) & (~ (z_out_38[6])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[58]) & (~ (z_out_38[5])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[57]) & (~ (z_out_38[4])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[56]) & (~ (z_out_38[3])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[55]) & (~ (z_out_38[2])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[54]) & (~ (z_out_38[1])))
      | ((return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[53]) & (~ (z_out_38[0])))
      | (return_mult_generic_AC_RND_CONV_false_2_p_1_sva_1[52:0]!=53'b00000000000000000000000000000000000000000000000000000);
  assign return_mult_generic_AC_RND_CONV_false_2_mux_13_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_2_if_1_or_nl,
      return_mult_generic_AC_RND_CONV_false_2_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_2_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_2_else_1_sticky_bit_or_nl,
      return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp[12]);
  assign return_mult_generic_AC_RND_CONV_false_2_or_nl = return_mult_generic_AC_RND_CONV_false_2_mux_13_nl
      | (z_out_53[1]);
  assign return_mult_generic_AC_RND_CONV_false_5_if_1_or_nl = (return_mult_generic_AC_RND_CONV_false_5_p_sva_1[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_or_2
      & (return_mult_generic_AC_RND_CONV_false_5_p_sva_1[51]));
  assign return_mult_generic_AC_RND_CONV_false_5_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_5_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_5_else_1_sticky_bit_or_nl
      = ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[105]) & (~ (z_out_38[52])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[104]) & (~ (z_out_38[51])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[103]) & (~ (z_out_38[50])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[102]) & (~ (z_out_38[49])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[101]) & (~ (z_out_38[48])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[100]) & (~ (z_out_38[47])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[99]) & (~ (z_out_38[46])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[98]) & (~ (z_out_38[45])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[97]) & (~ (z_out_38[44])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[96]) & (~ (z_out_38[43])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[95]) & (~ (z_out_38[42])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[94]) & (~ (z_out_38[41])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[93]) & (~ (z_out_38[40])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[92]) & (~ (z_out_38[39])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[91]) & (~ (z_out_38[38])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[90]) & (~ (z_out_38[37])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[89]) & (~ (z_out_38[36])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[88]) & (~ (z_out_38[35])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[87]) & (~ (z_out_38[34])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[86]) & (~ (z_out_38[33])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[85]) & (~ (z_out_38[32])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[84]) & (~ (z_out_38[31])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[83]) & (~ (z_out_38[30])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[82]) & (~ (z_out_38[29])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[81]) & (~ (z_out_38[28])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[80]) & (~ (z_out_38[27])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[79]) & (~ (z_out_38[26])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[78]) & (~ (z_out_38[25])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[77]) & (~ (z_out_38[24])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[76]) & (~ (z_out_38[23])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[75]) & (~ (z_out_38[22])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[74]) & (~ (z_out_38[21])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[73]) & (~ (z_out_38[20])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[72]) & (~ (z_out_38[19])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[71]) & (~ (z_out_38[18])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[70]) & (~ (z_out_38[17])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[69]) & (~ (z_out_38[16])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[68]) & (~ (z_out_38[15])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[67]) & (~ (z_out_38[14])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[66]) & (~ (z_out_38[13])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[65]) & (~ (z_out_38[12])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[64]) & (~ (z_out_38[11])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[63]) & (~ (z_out_38[10])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[62]) & (~ (z_out_38[9])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[61]) & (~ (z_out_38[8])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[60]) & (~ (z_out_38[7])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[59]) & (~ (z_out_38[6])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[58]) & (~ (z_out_38[5])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[57]) & (~ (z_out_38[4])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[56]) & (~ (z_out_38[3])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[55]) & (~ (z_out_38[2])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[54]) & (~ (z_out_38[1])))
      | ((return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[53]) & (~ (z_out_38[0])))
      | (return_mult_generic_AC_RND_CONV_false_5_p_1_sva_1[52:0]!=53'b00000000000000000000000000000000000000000000000000000);
  assign return_mult_generic_AC_RND_CONV_false_5_mux_13_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_5_if_1_or_nl,
      return_mult_generic_AC_RND_CONV_false_5_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_5_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_5_else_1_sticky_bit_or_nl,
      return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp[12]);
  assign return_mult_generic_AC_RND_CONV_false_5_or_nl = return_mult_generic_AC_RND_CONV_false_5_mux_13_nl
      | (z_out_53[1]);
  assign return_add_generic_AC_RND_CONV_false_10_op2_mu_and_3_nl = (~ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_tmp)
      & (fsm_output[23]);
  assign return_add_generic_AC_RND_CONV_false_10_op2_mu_and_4_nl = return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_tmp
      & (fsm_output[23]);
  assign return_add_generic_AC_RND_CONV_false_18_return_add_generic_AC_RND_CONV_false_18_and_5_nl
      = (return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_1[51])
      & (~ leading_sign_57_0_1_0_18_out_2);
  assign return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_2_nl
      = return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx6 | return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp;
  assign return_add_generic_AC_RND_CONV_false_24_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_22_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_22_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1 & return_add_generic_AC_RND_CONV_false_12_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_11_exp_and_3_nl = (~ and_352_tmp) &
      (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_11_exp_and_4_nl = and_352_tmp & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_and_8_nl
      = (return_add_generic_AC_RND_CONV_false_17_res_rounded_lpi_3_dfm_51_0_1[51])
      & (~ leading_sign_57_0_1_0_17_out_2);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nand_nl = ~((operator_33_true_34_acc_psp_1_sva_1[0])
      & return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nor_nl = ~((z_out_14[0])
      | (~ return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10));
  assign return_add_generic_AC_RND_CONV_false_17_mux_19_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nand_nl,
      return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nor_nl, return_add_generic_AC_RND_CONV_false_17_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_17_mux_19_nl | return_add_generic_AC_RND_CONV_false_17_e_r_qelse_or_svs_1);
  assign return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_and_4_nl
      = (operator_33_true_46_acc_tmp[0]) & return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_23_mux_20_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_and_4_nl,
      return_add_generic_AC_RND_CONV_false_23_exp_plus_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_23_res_rounded_acc_tmp[53]);
  assign or_319_nl = return_add_generic_AC_RND_CONV_false_23_r_inf_lpi_3_dfm_2 |
      operator_11_true_return_13_sva | and_dcpl_143 | operator_11_true_return_26_sva;
  assign return_add_generic_AC_RND_CONV_false_23_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs, or_319_nl);
  assign return_add_generic_AC_RND_CONV_false_23_e_r_return_add_generic_AC_RND_CONV_false_23_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_23_mux_20_nl & (~ return_add_generic_AC_RND_CONV_false_23_e_r_qelse_mux_1_nl))
      | return_add_generic_AC_RND_CONV_false_23_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_24_e_r_return_add_generic_AC_RND_CONV_false_24_e_r_or_1_nl
      = return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm
      | return_add_generic_AC_RND_CONV_false_21_unequal_tmp;
  assign return_add_generic_AC_RND_CONV_false_6_if_5_return_add_generic_AC_RND_CONV_false_6_if_5_and_nl
      = (return_add_generic_AC_RND_CONV_false_6_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_6_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_6_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_18_e_r_qelse_nand_nl = ~((operator_33_true_36_acc_psp_1_sva_1[0])
      & return_add_generic_AC_RND_CONV_false_18_acc_2_itm_10);
  assign return_add_generic_AC_RND_CONV_false_18_e_r_qelse_nor_nl = ~((operator_6_false_40_acc_psp_1_sva_1[0])
      | (~ return_add_generic_AC_RND_CONV_false_18_acc_2_itm_10));
  assign return_add_generic_AC_RND_CONV_false_18_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_18_e_r_qelse_nand_nl,
      return_add_generic_AC_RND_CONV_false_18_e_r_qelse_nor_nl, return_add_generic_AC_RND_CONV_false_18_res_rounded_acc_tmp[53]);
  assign return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_18_mux_13_nl | return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_svs_1);
  assign return_add_generic_AC_RND_CONV_false_24_return_add_generic_AC_RND_CONV_false_24_and_2_nl
      = (operator_33_true_48_acc_tmp[0]) & return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11;
  assign return_add_generic_AC_RND_CONV_false_24_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_24_return_add_generic_AC_RND_CONV_false_24_and_2_nl,
      return_add_generic_AC_RND_CONV_false_24_exp_plus_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_24_res_rounded_acc_tmp[53]);
  assign or_306_nl = or_dcpl_172 | and_dcpl_139 | return_add_generic_AC_RND_CONV_false_24_r_inf_lpi_3_dfm_2;
  assign return_add_generic_AC_RND_CONV_false_24_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs, or_306_nl);
  assign return_add_generic_AC_RND_CONV_false_24_e_r_qelse_return_add_generic_AC_RND_CONV_false_24_e_r_qelse_and_1_nl
      = return_add_generic_AC_RND_CONV_false_24_mux_13_nl & (~ return_add_generic_AC_RND_CONV_false_24_e_r_qelse_mux_1_nl);
  assign return_add_generic_AC_RND_CONV_false_25_e_r_return_add_generic_AC_RND_CONV_false_25_e_r_or_1_nl
      = return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm
      | return_add_generic_AC_RND_CONV_false_21_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_nl
      = (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w3!=11'b00000000000);
  assign return_add_generic_AC_RND_CONV_false_9_do_sub_return_add_generic_AC_RND_CONV_false_9_do_sub_xor_nl
      = (stage_PE_1_x_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1;
  assign return_add_generic_AC_RND_CONV_false_23_do_sub_return_add_generic_AC_RND_CONV_false_23_do_sub_xor_nl
      = (stage_PE_1_x_im_d_sva[63]) ^ operator_11_true_return_15_sva_mx2;
  assign return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_xnor_nl
      = ~((stage_PE_1_x_im_d_sva[63]) ^ operator_11_true_return_15_sva_mx1);
  assign return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_xnor_nl
      = ~((stage_PE_1_x_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2);
  assign return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_2_nl
      = BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx1 | return_add_generic_AC_RND_CONV_false_21_unequal_tmp;
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_mux1h_nl = MUX1HOT_v_4_9_2((return_add_generic_AC_RND_CONV_false_4_e_r_qelse_qr_10_1_lpi_3_dfm_1[9:6]),
      in_u_rsc_merge_sva_rsp_1_rsp_0, (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_mx0w2[9:6]),
      (stage_PE_1_x_im_d_sva[62:59]), return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_mx0w4_9_6,
      (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_mx1w0[9:6]),
      (operator_33_true_46_acc_tmp[10:7]), (return_add_generic_AC_RND_CONV_false_23_exp_plus_1_12_1_lpi_3_dfm_1[9:6]),
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1, {(fsm_output[8]) , or_1342_ssc , (fsm_output[13])
      , or_1344_ssc , (fsm_output[24]) , and_1813_cse , return_add_generic_AC_RND_CONV_false_4_e_r_qelse_and_cse
      , return_add_generic_AC_RND_CONV_false_4_e_r_qelse_and_1_cse , (fsm_output[31])});
  assign not_724_nl = ~ or_tmp;
  assign and_2115_nl = MUX_v_4_2_2(4'b0000, return_add_generic_AC_RND_CONV_false_4_e_r_qelse_mux1h_nl,
      not_724_nl);
  assign or_1486_nl = MUX_v_4_2_2(and_2115_nl, 4'b1111, or_tmp_829);
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_mux1h_1_nl = MUX1HOT_v_6_9_2((return_add_generic_AC_RND_CONV_false_4_e_r_qelse_qr_10_1_lpi_3_dfm_1[5:0]),
      in_u_rsc_merge_sva_rsp_1_rsp_1, (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_mx0w2[5:0]),
      (stage_PE_1_x_im_d_sva[58:53]), return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_mx0w4_5_0,
      (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_mx1w0[5:0]),
      (operator_33_true_46_acc_tmp[6:1]), (return_add_generic_AC_RND_CONV_false_23_exp_plus_1_12_1_lpi_3_dfm_1[5:0]),
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2, {(fsm_output[8]) , or_1342_ssc , (fsm_output[13])
      , or_1344_ssc , (fsm_output[24]) , and_1813_cse , return_add_generic_AC_RND_CONV_false_4_e_r_qelse_and_cse
      , return_add_generic_AC_RND_CONV_false_4_e_r_qelse_and_1_cse , (fsm_output[31])});
  assign not_725_nl = ~ or_tmp;
  assign and_2116_nl = MUX_v_6_2_2(6'b000000, return_add_generic_AC_RND_CONV_false_4_e_r_qelse_mux1h_1_nl,
      not_725_nl);
  assign or_1487_nl = MUX_v_6_2_2(and_2116_nl, 6'b111111, or_tmp_829);
  assign stage_PE_tmp_im_d_mux1h_1_nl = MUX1HOT_s_1_6_2(stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_0,
      (stage_PE_1_tmp_im_d_1_sva_1_63_51[1]), (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_1[0]),
      (z_out_24[0]), stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w4_0, (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_1[0]),
      {and_1585_rgt , and_1587_rgt , stage_PE_tmp_im_d_and_cse , stage_PE_tmp_im_d_or_cse
      , stage_PE_1_tmp_im_d_and_6_cse , stage_PE_tmp_im_d_and_2_cse});
  assign and_2118_nl = stage_PE_tmp_im_d_mux1h_1_nl & (~ or_tmp_830);
  assign stage_u_add_3_and_1_nl = (~ mode_lpi_1_dfm) & (fsm_output[8]);
  assign stage_u_add_3_and_3_nl = (fsm_output[8]) & (mode_lpi_1_dfm | return_add_generic_AC_RND_CONV_false_15_res_mant_or_1_cse
      | (fsm_output[12]) | (fsm_output[16]) | or_dcpl_505);
  assign operator_14_false_1_or_nl = (fsm_output[12]) | (fsm_output[14]) | (fsm_output[16])
      | (fsm_output[26]) | (fsm_output[28]);
  assign return_mult_generic_AC_RND_CONV_false_mux1h_2_nl = MUX1HOT_v_52_3_2((return_mult_generic_AC_RND_CONV_false_res_bef_rnd_3_53_1_lpi_3_dfm_1[52:1]),
      (return_mult_generic_AC_RND_CONV_false_3_res_bef_rnd_3_53_1_lpi_3_dfm_1[52:1]),
      (return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1[52:1]),
      {(fsm_output[10]) , (fsm_output[26]) , (fsm_output[36])});
  assign return_mult_generic_AC_RND_CONV_false_and_3_nl = (return_mult_generic_AC_RND_CONV_false_res_bef_rnd_3_53_1_lpi_3_dfm_1[0])
      & (return_mult_generic_AC_RND_CONV_false_mux_15 | (return_mult_generic_AC_RND_CONV_false_res_bef_rnd_3_53_1_lpi_3_dfm_1[1]));
  assign return_mult_generic_AC_RND_CONV_false_3_and_3_nl = (return_mult_generic_AC_RND_CONV_false_3_res_bef_rnd_3_53_1_lpi_3_dfm_1[0])
      & (return_mult_generic_AC_RND_CONV_false_mux_15 | (return_mult_generic_AC_RND_CONV_false_3_res_bef_rnd_3_53_1_lpi_3_dfm_1[1]));
  assign return_mult_generic_AC_RND_CONV_false_6_if_1_or_1_nl = (z_out_54[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_or_2
      & (z_out_54[51]));
  assign return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[51]))) | ((out_f_d_rsci_q_d[51])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[50]))) | ((out_f_d_rsci_q_d[50])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[49]))) | ((out_f_d_rsci_q_d[49])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[48]))) | ((out_f_d_rsci_q_d[48])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[47]))) | ((out_f_d_rsci_q_d[47])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[46]))) | ((out_f_d_rsci_q_d[46])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[45]))) | ((out_f_d_rsci_q_d[45])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[44]))) | ((out_f_d_rsci_q_d[44])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[43]))) | ((out_f_d_rsci_q_d[43])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[42]))) | ((out_f_d_rsci_q_d[42])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[41]))) | ((out_f_d_rsci_q_d[41])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[40]))) | ((out_f_d_rsci_q_d[40])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[39]))) | ((out_f_d_rsci_q_d[39])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[38]))) | ((out_f_d_rsci_q_d[38])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[37]))) | ((out_f_d_rsci_q_d[37])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[36]))) | ((out_f_d_rsci_q_d[36])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[35]))) | ((out_f_d_rsci_q_d[35])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[34]))) | ((out_f_d_rsci_q_d[34])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[33]))) | ((out_f_d_rsci_q_d[33])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[32]))) | ((out_f_d_rsci_q_d[32])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[31]))) | ((out_f_d_rsci_q_d[31])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[30]))) | ((out_f_d_rsci_q_d[30])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[29]))) | ((out_f_d_rsci_q_d[29])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[28]))) | ((out_f_d_rsci_q_d[28])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[27]))) | ((out_f_d_rsci_q_d[27])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[26]))) | ((out_f_d_rsci_q_d[26])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[25]))) | ((out_f_d_rsci_q_d[25])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[24]))) | ((out_f_d_rsci_q_d[24])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[23]))) | ((out_f_d_rsci_q_d[23])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[22]))) | ((out_f_d_rsci_q_d[22])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[21]))) | ((out_f_d_rsci_q_d[21])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[20]))) | ((out_f_d_rsci_q_d[20])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[19]))) | ((out_f_d_rsci_q_d[19])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[18]))) | ((out_f_d_rsci_q_d[18])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[17]))) | ((out_f_d_rsci_q_d[17])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[16]))) | ((out_f_d_rsci_q_d[16])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[15]))) | ((out_f_d_rsci_q_d[15])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[14]))) | ((out_f_d_rsci_q_d[14])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[13]))) | ((out_f_d_rsci_q_d[13])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[12]))) | ((out_f_d_rsci_q_d[12])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[11]))) | ((out_f_d_rsci_q_d[11])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[10]))) | ((out_f_d_rsci_q_d[10])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[9]))) | ((out_f_d_rsci_q_d[9])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[8]))) | ((out_f_d_rsci_q_d[8])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[7]))) | ((out_f_d_rsci_q_d[7])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[6]))) | ((out_f_d_rsci_q_d[6])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[5]))) | ((out_f_d_rsci_q_d[5])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[4]))) | ((out_f_d_rsci_q_d[4])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[3]))) | ((out_f_d_rsci_q_d[3])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[2]))) | ((out_f_d_rsci_q_d[2])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[1]))) | ((out_f_d_rsci_q_d[1])
      & (~ (return_mult_generic_AC_RND_CONV_false_6_else_1_lshift_itm[0]))) | (out_f_d_rsci_q_d[0]);
  assign return_mult_generic_AC_RND_CONV_false_6_mux_12_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_6_if_1_or_1_nl,
      return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_or_1_nl,
      z_out_51[11]);
  assign return_mult_generic_AC_RND_CONV_false_6_and_3_nl = (return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1[0])
      & (return_mult_generic_AC_RND_CONV_false_6_mux_12_nl | (return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1[1]));
  assign return_mult_generic_AC_RND_CONV_false_mux1h_3_nl = MUX1HOT_s_1_3_2(return_mult_generic_AC_RND_CONV_false_and_3_nl,
      return_mult_generic_AC_RND_CONV_false_3_and_3_nl, return_mult_generic_AC_RND_CONV_false_6_and_3_nl,
      {(fsm_output[10]) , (fsm_output[26]) , (fsm_output[36])});
  assign nl_z_out = return_mult_generic_AC_RND_CONV_false_mux1h_2_nl + conv_u2u_1_52(return_mult_generic_AC_RND_CONV_false_mux1h_3_nl);
  assign z_out = nl_z_out[51:0];
  assign operator_32_false_operator_32_false_or_3_nl = MUX_v_4_2_2((in_u_rsc_merge_sva_rsp_0[5:2]),
      4'b1111, or_1495_cse_1);
  assign operator_32_false_mux_7_nl = MUX_v_6_2_2((~ in_u_rsc_merge_sva_rsp_0), in_u_rsc_merge_sva_rsp_0,
      or_1495_cse_1);
  assign operator_32_false_mux_8_nl = MUX_v_4_2_2((~ in_u_rsc_merge_sva_rsp_1_rsp_0),
      in_u_rsc_merge_sva_rsp_1_rsp_0, or_1495_cse_1);
  assign operator_32_false_mux_9_nl = MUX_v_6_2_2((~ in_u_rsc_merge_sva_rsp_1_rsp_1),
      in_u_rsc_merge_sva_rsp_1_rsp_1, or_1495_cse_1);
  assign nl_z_out_1 = ({1'b1 , ({{1{or_1495_cse_1}}, or_1495_cse_1}) , 2'b00 , ({{7{or_1495_cse_1}},
      or_1495_cse_1}) , operator_32_false_operator_32_false_or_3_nl}) + conv_u2u_16_17({operator_32_false_mux_7_nl
      , operator_32_false_mux_8_nl , operator_32_false_mux_9_nl});
  assign z_out_1 = nl_z_out_1[16:0];
  assign return_add_generic_AC_RND_CONV_false_9_ma1_lt_ma2_mux_4_nl = MUX_s_1_2_2((~
      return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0), (~ return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0),
      fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_9_ma1_lt_ma2_mux_5_nl = MUX_v_51_2_2((~
      return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1), (~ return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1),
      fsm_output[29]);
  assign nl_acc_2_nl = ({1'b1 , (stage_PE_1_x_re_d_sva[51:0]) , 1'b1}) + conv_u2u_53_54({return_add_generic_AC_RND_CONV_false_9_ma1_lt_ma2_mux_4_nl
      , return_add_generic_AC_RND_CONV_false_9_ma1_lt_ma2_mux_5_nl , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[53:0];
  assign z_out_2_52 = readslicef_54_1_53(acc_2_nl);
  assign return_add_generic_AC_RND_CONV_false_3_ma1_lt_ma2_mux_3_nl = MUX_v_52_2_2((~
      (out_f_d_rsci_q_d[51:0])), (~ (in_f_d_rsci_q_d[51:0])), fsm_output[22]);
  assign nl_acc_3_nl = ({1'b1 , (stage_PE_1_x_im_d_sva[51:0]) , 1'b1}) + conv_u2u_53_54({return_add_generic_AC_RND_CONV_false_3_ma1_lt_ma2_mux_3_nl
      , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[53:0];
  assign z_out_3_52 = readslicef_54_1_53(acc_3_nl);
  assign return_add_generic_AC_RND_CONV_false_17_mux_32_nl = MUX_v_5_2_2(return_add_generic_AC_RND_CONV_false_17_mux_7_itm_55_51,
      return_add_generic_AC_RND_CONV_false_18_mux_1_itm_55_51, fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_17_mux_33_nl = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0,
      return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0, fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_17_mux_34_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm, fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_17_mux_35_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_12_do_sub_sva,
      return_add_generic_AC_RND_CONV_false_10_do_sub_sva, fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_17_mux_36_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm, fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_17_mux_37_nl = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[50]),
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm, fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_17_mux_38_nl = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[49:0]),
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm, fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_17_mux_39_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm, fsm_output[30]);
  assign nl_acc_5_nl = ({return_add_generic_AC_RND_CONV_false_17_mux_32_nl , return_add_generic_AC_RND_CONV_false_17_mux_33_nl
      , return_add_generic_AC_RND_CONV_false_17_mux_34_nl , return_add_generic_AC_RND_CONV_false_17_mux_35_nl})
      + conv_u2u_57_58({return_add_generic_AC_RND_CONV_false_17_mux_36_nl , return_add_generic_AC_RND_CONV_false_17_mux_37_nl
      , return_add_generic_AC_RND_CONV_false_17_mux_38_nl , return_add_generic_AC_RND_CONV_false_17_mux_39_nl
      , 4'b0001});
  assign acc_5_nl = nl_acc_5_nl[57:0];
  assign z_out_5 = readslicef_58_57_1(acc_5_nl);
  assign return_add_generic_AC_RND_CONV_false_18_mux_23_nl = MUX_v_5_2_2(return_add_generic_AC_RND_CONV_false_18_mux_1_itm_55_51,
      return_add_generic_AC_RND_CONV_false_17_mux_7_itm_55_51, fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_18_mux_24_nl = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0,
      return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0, fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_18_mux_25_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm, fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_18_mux_26_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_do_sub_sva,
      return_add_generic_AC_RND_CONV_false_12_do_sub_sva, fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_18_mux_27_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm, fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_18_mux_28_nl = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[50]),
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm, fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_18_mux_29_nl = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[49:0]),
      reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1,
      fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_18_mux_30_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm, fsm_output[30]);
  assign nl_acc_6_nl = ({return_add_generic_AC_RND_CONV_false_18_mux_23_nl , return_add_generic_AC_RND_CONV_false_18_mux_24_nl
      , return_add_generic_AC_RND_CONV_false_18_mux_25_nl , return_add_generic_AC_RND_CONV_false_18_mux_26_nl})
      + conv_u2u_57_58({return_add_generic_AC_RND_CONV_false_18_mux_27_nl , return_add_generic_AC_RND_CONV_false_18_mux_28_nl
      , return_add_generic_AC_RND_CONV_false_18_mux_29_nl , return_add_generic_AC_RND_CONV_false_18_mux_30_nl
      , 4'b0001});
  assign acc_6_nl = nl_acc_6_nl[57:0];
  assign z_out_6 = readslicef_58_57_1(acc_6_nl);
  assign return_add_generic_AC_RND_CONV_false_1_or_13_nl = return_add_generic_AC_RND_CONV_false_1_and_8_cse
      | return_add_generic_AC_RND_CONV_false_1_and_14_cse;
  assign return_add_generic_AC_RND_CONV_false_1_or_14_nl = return_add_generic_AC_RND_CONV_false_1_and_9_cse
      | return_add_generic_AC_RND_CONV_false_1_and_15_cse;
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_20_nl = MUX1HOT_v_56_4_2((z_out_29[56:1]),
      (~ (z_out_29[56:1])), (z_out_30[56:1]), (~ (z_out_30[56:1])), {return_add_generic_AC_RND_CONV_false_3_or_4_cse
      , return_add_generic_AC_RND_CONV_false_3_or_5_cse , return_add_generic_AC_RND_CONV_false_1_or_13_nl
      , return_add_generic_AC_RND_CONV_false_1_or_14_nl});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_21_nl = MUX1HOT_s_1_12_2(return_add_generic_AC_RND_CONV_false_1_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_1_res_mant_3_0_sva_1), (~ return_add_generic_AC_RND_CONV_false_2_res_mant_3_0_sva_1),
      return_add_generic_AC_RND_CONV_false_2_res_mant_3_0_sva_1, return_add_generic_AC_RND_CONV_false_9_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_9_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_14_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_14_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_13_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_13_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_22_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_22_res_mant_3_0_sva_1), {return_add_generic_AC_RND_CONV_false_3_and_cse
      , return_add_generic_AC_RND_CONV_false_3_and_1_cse , return_add_generic_AC_RND_CONV_false_3_and_2_cse
      , return_add_generic_AC_RND_CONV_false_3_and_3_cse , return_add_generic_AC_RND_CONV_false_1_and_8_cse
      , return_add_generic_AC_RND_CONV_false_1_and_9_cse , return_add_generic_AC_RND_CONV_false_3_and_4_cse
      , return_add_generic_AC_RND_CONV_false_3_and_5_cse , return_add_generic_AC_RND_CONV_false_3_and_6_cse
      , return_add_generic_AC_RND_CONV_false_3_and_7_cse , return_add_generic_AC_RND_CONV_false_1_and_14_cse
      , return_add_generic_AC_RND_CONV_false_1_and_15_cse});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_22_nl = MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1,
      return_add_generic_AC_RND_CONV_false_2_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_10_op2_inf_sva,
      return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_13_do_sub_sva_1,
      return_add_generic_AC_RND_CONV_false_15_do_sub_sva, {(fsm_output[6]) , (fsm_output[8])
      , (fsm_output[13]) , (fsm_output[22]) , (fsm_output[24]) , (fsm_output[29])});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_23_nl = MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_3_op_bigger_mux_1_cse,
      return_add_generic_AC_RND_CONV_false_op_bigger_mux_1_cse, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_16_op_bigger_mux_1_cse,
      return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_1_cse, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm,
      return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0, {(fsm_output[6])
      , (fsm_output[8]) , return_add_generic_AC_RND_CONV_false_1_and_28_cse , and_1132_ssc
      , (fsm_output[22]) , (fsm_output[24]) , return_add_generic_AC_RND_CONV_false_1_and_30_cse
      , and_1145_ssc});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_24_nl = MUX1HOT_s_1_8_2((return_add_generic_AC_RND_CONV_false_3_op_bigger_mux_2_cse[50]),
      (return_add_generic_AC_RND_CONV_false_op_bigger_mux_2_cse[50]), (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[50]),
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_16_op_bigger_mux_2_cse[50]),
      (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_cse[50]), (return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0[50]),
      return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0, {(fsm_output[6])
      , (fsm_output[8]) , return_add_generic_AC_RND_CONV_false_1_and_28_cse , and_1132_ssc
      , (fsm_output[22]) , (fsm_output[24]) , return_add_generic_AC_RND_CONV_false_1_and_30_cse
      , and_1145_ssc});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_25_nl = MUX1HOT_v_50_8_2((return_add_generic_AC_RND_CONV_false_3_op_bigger_mux_2_cse[49:0]),
      (return_add_generic_AC_RND_CONV_false_op_bigger_mux_2_cse[49:0]), (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[49:0]),
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_16_op_bigger_mux_2_cse[49:0]),
      (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_cse[49:0]), (return_add_generic_AC_RND_CONV_false_17_mux_7_itm_50_0[49:0]),
      return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0, {(fsm_output[6])
      , (fsm_output[8]) , return_add_generic_AC_RND_CONV_false_1_and_28_cse , and_1132_ssc
      , (fsm_output[22]) , (fsm_output[24]) , return_add_generic_AC_RND_CONV_false_1_and_30_cse
      , and_1145_ssc});
  assign return_add_generic_AC_RND_CONV_false_1_or_15_nl = return_add_generic_AC_RND_CONV_false_3_and_30_cse
      | return_add_generic_AC_RND_CONV_false_3_and_32_cse;
  assign return_add_generic_AC_RND_CONV_false_1_or_16_nl = return_add_generic_AC_RND_CONV_false_1_and_28_cse
      | return_add_generic_AC_RND_CONV_false_1_and_30_cse;
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_26_nl = MUX1HOT_s_1_7_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1,
      {return_add_generic_AC_RND_CONV_false_1_or_15_nl , return_add_generic_AC_RND_CONV_false_3_or_14_cse
      , or_956_cse , return_add_generic_AC_RND_CONV_false_1_or_16_nl , and_1132_ssc
      , return_add_generic_AC_RND_CONV_false_3_or_16_cse , and_1145_ssc});
  assign nl_acc_7_nl = ({return_add_generic_AC_RND_CONV_false_1_mux1h_20_nl , return_add_generic_AC_RND_CONV_false_1_mux1h_21_nl
      , return_add_generic_AC_RND_CONV_false_1_mux1h_22_nl}) + conv_u2u_57_58({return_add_generic_AC_RND_CONV_false_1_mux1h_23_nl
      , return_add_generic_AC_RND_CONV_false_1_mux1h_24_nl , return_add_generic_AC_RND_CONV_false_1_mux1h_25_nl
      , return_add_generic_AC_RND_CONV_false_1_mux1h_26_nl , 4'b0001});
  assign acc_7_nl = nl_acc_7_nl[57:0];
  assign z_out_7 = readslicef_58_57_1(acc_7_nl);
  assign return_add_generic_AC_RND_CONV_false_20_op_bigger_mux_7_tmp = MUX_s_1_2_2(or_450_cse,
      return_add_generic_AC_RND_CONV_false_7_op1_smaller_lor_lpi_3_dfm_2, fsm_output[12]);
  assign return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_nor_1_nl
      = ~(return_add_generic_AC_RND_CONV_false_12_mux_itm | (fsm_output[16]));
  assign return_add_generic_AC_RND_CONV_false_7_and_4_nl = return_add_generic_AC_RND_CONV_false_12_mux_itm
      & (~ (fsm_output[16]));
  assign return_add_generic_AC_RND_CONV_false_7_and_5_nl = (~ return_add_generic_AC_RND_CONV_false_12_do_sub_sva)
      & (fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_7_and_6_nl = return_add_generic_AC_RND_CONV_false_12_do_sub_sva
      & (fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_mux1h_1_nl
      = MUX1HOT_v_56_4_2((return_add_generic_AC_RND_CONV_false_7_rshift_itm[56:1]),
      (~ (return_add_generic_AC_RND_CONV_false_7_rshift_itm[56:1])), (z_out_32[56:1]),
      (~ (z_out_32[56:1])), {return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_nor_1_nl
      , return_add_generic_AC_RND_CONV_false_7_and_4_nl , return_add_generic_AC_RND_CONV_false_7_and_5_nl
      , return_add_generic_AC_RND_CONV_false_7_and_6_nl});
  assign return_add_generic_AC_RND_CONV_false_7_mux_41_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_7_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_12_mux_itm);
  assign return_add_generic_AC_RND_CONV_false_12_mux_23_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_sticky_bit_return_add_generic_AC_RND_CONV_false_11_sticky_bit_return_add_generic_AC_RND_CONV_false_11_sticky_bit_or_cse,
      (~ return_add_generic_AC_RND_CONV_false_11_sticky_bit_return_add_generic_AC_RND_CONV_false_11_sticky_bit_return_add_generic_AC_RND_CONV_false_11_sticky_bit_or_cse),
      return_add_generic_AC_RND_CONV_false_12_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_7_mux_40_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_mux_41_nl,
      return_add_generic_AC_RND_CONV_false_12_mux_23_nl, fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_7_mux_42_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_12_mux_itm,
      return_add_generic_AC_RND_CONV_false_12_do_sub_sva, fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_7_op_bigger_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_7_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_7_mux_43_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_op_bigger_mux_13_nl,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm, fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_7_op_bigger_mux_14_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_7_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_7_mux_44_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_op_bigger_mux_14_nl,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm, fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_7_and_nl = return_add_generic_AC_RND_CONV_false_20_op_bigger_mux_7_tmp
      & (~ (fsm_output[16]));
  assign return_add_generic_AC_RND_CONV_false_7_mux_45_nl = MUX_v_50_2_2(reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_7_and_nl);
  assign return_add_generic_AC_RND_CONV_false_7_op_bigger_mux_15_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_7_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_7_mux_46_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_op_bigger_mux_15_nl,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm, fsm_output[16]);
  assign nl_acc_8_nl = ({return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_mux1h_1_nl
      , return_add_generic_AC_RND_CONV_false_7_mux_40_nl , return_add_generic_AC_RND_CONV_false_7_mux_42_nl})
      + conv_u2u_57_58({return_add_generic_AC_RND_CONV_false_7_mux_43_nl , return_add_generic_AC_RND_CONV_false_7_mux_44_nl
      , return_add_generic_AC_RND_CONV_false_7_mux_45_nl , return_add_generic_AC_RND_CONV_false_7_mux_46_nl
      , 4'b0001});
  assign acc_8_nl = nl_acc_8_nl[57:0];
  assign z_out_8 = readslicef_58_57_1(acc_8_nl);
  assign return_add_generic_AC_RND_CONV_false_11_or_7_nl = return_add_generic_AC_RND_CONV_false_11_and_45_cse
      | return_add_generic_AC_RND_CONV_false_11_and_1_cse;
  assign return_add_generic_AC_RND_CONV_false_11_or_8_nl = return_add_generic_AC_RND_CONV_false_11_and_46_cse
      | return_add_generic_AC_RND_CONV_false_11_and_2_cse;
  assign return_add_generic_AC_RND_CONV_false_11_mux1h_17_nl = MUX1HOT_v_56_4_2((z_out_32[56:1]),
      (~ (z_out_32[56:1])), (return_add_generic_AC_RND_CONV_false_20_rshift_itm[56:1]),
      (~ (return_add_generic_AC_RND_CONV_false_20_rshift_itm[56:1])), {return_add_generic_AC_RND_CONV_false_11_or_7_nl
      , return_add_generic_AC_RND_CONV_false_11_or_8_nl , return_add_generic_AC_RND_CONV_false_11_and_3_cse
      , return_add_generic_AC_RND_CONV_false_11_and_4_cse});
  assign return_add_generic_AC_RND_CONV_false_11_mux1h_18_nl = MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_11_sticky_bit_return_add_generic_AC_RND_CONV_false_11_sticky_bit_return_add_generic_AC_RND_CONV_false_11_sticky_bit_or_cse,
      (~ return_add_generic_AC_RND_CONV_false_11_sticky_bit_return_add_generic_AC_RND_CONV_false_11_sticky_bit_return_add_generic_AC_RND_CONV_false_11_sticky_bit_or_cse),
      return_add_generic_AC_RND_CONV_false_19_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_19_res_mant_3_0_sva_1),
      return_add_generic_AC_RND_CONV_false_20_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_20_res_mant_3_0_sva_1),
      {return_add_generic_AC_RND_CONV_false_11_and_45_cse , return_add_generic_AC_RND_CONV_false_11_and_46_cse
      , return_add_generic_AC_RND_CONV_false_11_and_1_cse , return_add_generic_AC_RND_CONV_false_11_and_2_cse
      , return_add_generic_AC_RND_CONV_false_11_and_3_cse , return_add_generic_AC_RND_CONV_false_11_and_4_cse});
  assign return_add_generic_AC_RND_CONV_false_11_mux1h_19_nl = MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_13_do_sub_sva,
      return_add_generic_AC_RND_CONV_false_10_do_sub_sva, return_add_generic_AC_RND_CONV_false_12_mux_itm,
      {(fsm_output[14]) , (fsm_output[26]) , (fsm_output[28])});
  assign return_add_generic_AC_RND_CONV_false_11_mux1h_20_nl = MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm,
      return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1, {(fsm_output[14])
      , return_add_generic_AC_RND_CONV_false_11_or_cse , return_add_generic_AC_RND_CONV_false_11_and_12_cse
      , and_1029_cse});
  assign return_add_generic_AC_RND_CONV_false_11_mux1h_21_nl = MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm,
      return_add_generic_AC_RND_CONV_false_14_op1_mu_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0, {(fsm_output[14])
      , return_add_generic_AC_RND_CONV_false_11_or_cse , return_add_generic_AC_RND_CONV_false_11_and_12_cse
      , and_1029_cse});
  assign return_add_generic_AC_RND_CONV_false_11_or_9_nl = (fsm_output[14]) | return_add_generic_AC_RND_CONV_false_11_and_11_cse
      | ((~ return_add_generic_AC_RND_CONV_false_20_op_bigger_mux_7_tmp) & (fsm_output[28]));
  assign return_add_generic_AC_RND_CONV_false_11_and_48_nl = return_add_generic_AC_RND_CONV_false_20_op_bigger_mux_7_tmp
      & (fsm_output[28]);
  assign return_add_generic_AC_RND_CONV_false_11_mux1h_22_nl = MUX1HOT_v_50_3_2(reg_return_add_generic_AC_RND_CONV_false_18_res_rounded_lpi_3_dfm_51_0_ftd_1,
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0,
      {return_add_generic_AC_RND_CONV_false_11_or_9_nl , return_add_generic_AC_RND_CONV_false_11_and_12_cse
      , return_add_generic_AC_RND_CONV_false_11_and_48_nl});
  assign return_add_generic_AC_RND_CONV_false_11_mux1h_23_nl = MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm,
      return_add_generic_AC_RND_CONV_false_19_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1,
      {(fsm_output[14]) , return_add_generic_AC_RND_CONV_false_11_and_11_cse , return_add_generic_AC_RND_CONV_false_11_and_12_cse
      , return_add_generic_AC_RND_CONV_false_11_and_13_cse , and_1029_cse});
  assign nl_acc_9_nl = ({return_add_generic_AC_RND_CONV_false_11_mux1h_17_nl , return_add_generic_AC_RND_CONV_false_11_mux1h_18_nl
      , return_add_generic_AC_RND_CONV_false_11_mux1h_19_nl}) + conv_u2u_57_58({return_add_generic_AC_RND_CONV_false_11_mux1h_20_nl
      , return_add_generic_AC_RND_CONV_false_11_mux1h_21_nl , return_add_generic_AC_RND_CONV_false_11_mux1h_22_nl
      , return_add_generic_AC_RND_CONV_false_11_mux1h_23_nl , 4'b0001});
  assign acc_9_nl = nl_acc_9_nl[57:0];
  assign z_out_9 = readslicef_58_57_1(acc_9_nl);
  assign nl_z_out_12 = (z_out_14[10:1]) + 10'b0000000001;
  assign z_out_12 = nl_z_out_12[9:0];
  assign for_mux1h_11_nl = MUX1HOT_s_1_4_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[10]),
      (in_u_rsc_merge_sva_rsp_1_rsp_0[3]), (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0[8]),
      (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1[3]), {or_1531_cse , (fsm_output[15])
      , for_or_5_cse , (fsm_output[17])});
  assign for_and_4_nl = for_mux1h_11_nl & (~ (fsm_output[8])) & (~ mode_or_cse);
  assign for_mux1h_12_nl = MUX1HOT_v_3_5_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[9:7]),
      (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0[8:6]), (in_u_rsc_merge_sva_rsp_1_rsp_0[2:0]),
      (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0[7:5]), (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1[2:0]),
      {or_1531_cse , (fsm_output[8]) , (fsm_output[15]) , for_or_5_cse , (fsm_output[17])});
  assign not_889_nl = ~ mode_or_cse;
  assign for_and_5_nl = MUX_v_3_2_2(3'b000, for_mux1h_12_nl, not_889_nl);
  assign for_mux1h_13_nl = MUX1HOT_v_5_5_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[6:2]),
      (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0[5:1]), (in_u_rsc_merge_sva_rsp_1_rsp_1[5:1]),
      (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0[4:0]), (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[5:1]),
      {or_1531_cse , (fsm_output[8]) , (fsm_output[15]) , for_or_5_cse , (fsm_output[17])});
  assign not_890_nl = ~ mode_or_cse;
  assign for_and_6_nl = MUX_v_5_2_2(5'b00000, for_mux1h_13_nl, not_890_nl);
  assign for_mux1h_14_nl = MUX1HOT_s_1_5_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[1]),
      (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0[0]), (in_u_rsc_merge_sva_rsp_1_rsp_1[0]),
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1, (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[0]),
      {or_1531_cse , (fsm_output[8]) , (fsm_output[15]) , for_or_5_cse , (fsm_output[17])});
  assign for_and_7_nl = for_mux1h_14_nl & (~ mode_or_cse);
  assign for_mux1h_15_nl = MUX1HOT_s_1_5_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[0]),
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1, return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm,
      drf_qr_lval_14_smx_0_lpi_3_dfm, drf_qr_lval_12_smx_0_lpi_3_dfm, {or_1531_cse
      , (fsm_output[8]) , (fsm_output[15]) , for_or_5_cse , (fsm_output[17])});
  assign for_or_14_nl = for_mux1h_15_nl | mode_or_cse;
  assign for_or_15_nl = (~(mode_or_cse | or_1531_cse)) | (fsm_output[8]) | (fsm_output[15])
      | (fsm_output[16]) | (fsm_output[17]) | (fsm_output[30]);
  assign for_mux_1_nl = MUX_s_1_2_2((for_i_3_0_sva[3]), (operator_6_false_6_operator_6_false_6_conc_2_6_1[5]),
      or_1531_cse);
  assign for_for_or_1_nl = for_mux_1_nl | (fsm_output[8]) | (fsm_output[15]) | (fsm_output[16])
      | (fsm_output[17]) | (fsm_output[30]);
  assign for_mux1h_16_nl = MUX1HOT_s_1_5_2((for_i_3_0_sva[3]), (operator_6_false_6_operator_6_false_6_conc_2_6_1[4]),
      (~ (return_add_generic_AC_RND_CONV_false_20_ls_sva[5])), (~ return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_0),
      (~ (leading_sign_57_0_1_0_15_out_3[5])), {mode_or_cse , or_1531_cse , for_or_4_cse
      , for_or_10_cse_1 , (fsm_output[30])});
  assign for_mux1h_17_nl = MUX1HOT_s_1_5_2((for_i_3_0_sva[3]), (operator_6_false_6_operator_6_false_6_conc_2_6_1[3]),
      (~ (return_add_generic_AC_RND_CONV_false_20_ls_sva[4])), (~ return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_1),
      (~ (leading_sign_57_0_1_0_15_out_3[4])), {mode_or_cse , or_1531_cse , for_or_4_cse
      , for_or_10_cse_1 , (fsm_output[30])});
  assign for_mux1h_18_nl = MUX1HOT_s_1_5_2((for_i_3_0_sva[3]), (operator_6_false_6_operator_6_false_6_conc_2_6_1[2]),
      (~ (return_add_generic_AC_RND_CONV_false_20_ls_sva[3])), (~ (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2[3])),
      (~ (leading_sign_57_0_1_0_15_out_3[3])), {mode_or_cse , or_1531_cse , for_or_4_cse
      , for_or_10_cse_1 , (fsm_output[30])});
  assign for_mux1h_19_nl = MUX1HOT_v_2_5_2((for_i_3_0_sva[2:1]), (operator_6_false_6_operator_6_false_6_conc_2_6_1[1:0]),
      (~ (return_add_generic_AC_RND_CONV_false_20_ls_sva[2:1])), (~ (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2[2:1])),
      (~ (leading_sign_57_0_1_0_15_out_3[2:1])), {mode_or_cse , or_1531_cse , for_or_4_cse
      , for_or_10_cse_1 , (fsm_output[30])});
  assign for_mux1h_20_nl = MUX1HOT_s_1_5_2((for_i_3_0_sva[0]), (~ (leading_sign_57_0_1_0_15_out_3[0])),
      (~ (return_add_generic_AC_RND_CONV_false_20_ls_sva[0])), (~ (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2[0])),
      (~ (leading_sign_57_0_1_0_15_out_3[0])), {mode_or_cse , or_1531_cse , for_or_4_cse
      , for_or_10_cse_1 , (fsm_output[30])});
  assign nl_acc_11_nl = conv_u2u_12_14({for_and_4_nl , for_and_5_nl , for_and_6_nl
      , for_and_7_nl , for_or_14_nl , for_or_15_nl}) + conv_s2u_8_14({for_for_or_1_nl
      , for_mux1h_16_nl , for_mux1h_17_nl , for_mux1h_18_nl , for_mux1h_19_nl , for_mux1h_20_nl
      , 1'b1});
  assign acc_11_nl = nl_acc_11_nl[13:0];
  assign z_out_13 = readslicef_14_13_1(acc_11_nl);
  assign operator_6_false_9_mux_6_nl = MUX_s_1_2_2((~ return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_0),
      (~ (leading_sign_57_0_1_0_17_out_3[5])), fsm_output[23]);
  assign operator_6_false_9_mux_7_nl = MUX_s_1_2_2((~ return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_1),
      (~ (leading_sign_57_0_1_0_17_out_3[4])), fsm_output[23]);
  assign operator_6_false_9_mux_8_nl = MUX_v_4_2_2((~ return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2),
      (~ (leading_sign_57_0_1_0_17_out_3[3:0])), fsm_output[23]);
  assign nl_acc_12_nl = conv_u2u_11_12({reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1 ,
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2 , 1'b1}) + conv_s2u_8_12({1'b1 , operator_6_false_9_mux_6_nl
      , operator_6_false_9_mux_7_nl , operator_6_false_9_mux_8_nl , 1'b1});
  assign acc_12_nl = nl_acc_12_nl[11:0];
  assign z_out_14 = readslicef_12_11_1(acc_12_nl);
  assign operator_6_false_19_mux_5_nl = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_7_op_bigger_mux_6_itm[10]),
      drf_qr_lval_10_smx_lpi_3_dfm_mx2_10, fsm_output[28]);
  assign operator_6_false_19_mux_6_nl = MUX_v_4_2_2((return_add_generic_AC_RND_CONV_false_7_op_bigger_mux_6_itm[9:6]),
      drf_qr_lval_10_smx_lpi_3_dfm_mx2_9_6, fsm_output[28]);
  assign operator_6_false_19_mux_7_nl = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_7_op_bigger_mux_6_itm[5:0]),
      drf_qr_lval_10_smx_lpi_3_dfm_mx2_5_0, fsm_output[28]);
  assign nl_operator_6_false_19_acc_1_nl = ({1'b1 , (~ (leading_sign_57_0_1_0_8_out_3[5:1]))})
      + 6'b000001;
  assign operator_6_false_19_acc_1_nl = nl_operator_6_false_19_acc_1_nl[5:0];
  assign nl_operator_6_false_48_acc_1_nl = ({1'b1 , (~ (leading_sign_57_0_1_0_21_out_3[5:1]))})
      + 6'b000001;
  assign operator_6_false_48_acc_1_nl = nl_operator_6_false_48_acc_1_nl[5:0];
  assign operator_6_false_19_mux_8_nl = MUX_v_6_2_2(operator_6_false_19_acc_1_nl,
      operator_6_false_48_acc_1_nl, fsm_output[28]);
  assign operator_6_false_19_mux_9_nl = MUX_s_1_2_2((~ (leading_sign_57_0_1_0_8_out_3[0])),
      (~ (leading_sign_57_0_1_0_21_out_3[0])), fsm_output[28]);
  assign nl_z_out_15 = conv_u2u_11_13({operator_6_false_19_mux_5_nl , operator_6_false_19_mux_6_nl
      , operator_6_false_19_mux_7_nl}) + conv_s2u_7_13({operator_6_false_19_mux_8_nl
      , operator_6_false_19_mux_9_nl});
  assign z_out_15 = nl_z_out_15[12:0];
  assign operator_6_false_17_mux1h_7_nl = MUX1HOT_s_1_5_2(drf_qr_lval_10_smx_lpi_3_dfm_mx1_10,
      (return_add_generic_AC_RND_CONV_false_10_exp_conc_5_itm_10_7[3]), (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1[3]),
      (drf_qr_lval_26_smx_lpi_3_dfm_mx0[10]), drf_qr_lval_6_smx_lpi_3_dfm_mx0_10,
      {(fsm_output[12]) , (fsm_output[14]) , (fsm_output[16]) , (fsm_output[28])
      , (fsm_output[26])});
  assign operator_6_false_17_mux1h_8_nl = MUX1HOT_v_3_5_2((drf_qr_lval_10_smx_lpi_3_dfm_mx1_9_6[3:1]),
      (return_add_generic_AC_RND_CONV_false_10_exp_conc_5_itm_10_7[2:0]), (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1[2:0]),
      (drf_qr_lval_26_smx_lpi_3_dfm_mx0[9:7]), (drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_0[9:7]),
      {(fsm_output[12]) , (fsm_output[14]) , (fsm_output[16]) , (fsm_output[28])
      , (fsm_output[26])});
  assign operator_6_false_17_mux1h_9_nl = MUX1HOT_s_1_5_2((drf_qr_lval_10_smx_lpi_3_dfm_mx1_9_6[0]),
      (return_add_generic_AC_RND_CONV_false_10_exp_conc_5_itm_6_1[5]), (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[5]),
      (drf_qr_lval_26_smx_lpi_3_dfm_mx0[6]), (drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_0[6]),
      {(fsm_output[12]) , (fsm_output[14]) , (fsm_output[16]) , (fsm_output[28])
      , (fsm_output[26])});
  assign operator_6_false_17_mux1h_10_nl = MUX1HOT_v_5_5_2((drf_qr_lval_10_smx_lpi_3_dfm_mx1_5_0[5:1]),
      (return_add_generic_AC_RND_CONV_false_10_exp_conc_5_itm_6_1[4:0]), (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2[4:0]),
      (drf_qr_lval_26_smx_lpi_3_dfm_mx0[5:1]), (drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_0[5:1]),
      {(fsm_output[12]) , (fsm_output[14]) , (fsm_output[16]) , (fsm_output[28])
      , (fsm_output[26])});
  assign operator_6_false_17_mux1h_11_nl = MUX1HOT_s_1_5_2((drf_qr_lval_10_smx_lpi_3_dfm_mx1_5_0[0]),
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm_mx1,
      drf_qr_lval_12_smx_0_lpi_3_dfm, (drf_qr_lval_26_smx_lpi_3_dfm_mx0[0]), (drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_0[0]),
      {(fsm_output[12]) , (fsm_output[14]) , (fsm_output[16]) , (fsm_output[28])
      , (fsm_output[26])});
  assign nl_operator_6_false_17_acc_1_nl = ({1'b1 , (~ (rtn_out_1[5:1]))}) + 6'b000001;
  assign operator_6_false_17_acc_1_nl = nl_operator_6_false_17_acc_1_nl[5:0];
  assign nl_operator_6_false_23_acc_1_nl = ({1'b1 , (~ (leading_sign_57_0_1_0_10_out_3[5:1]))})
      + 6'b000001;
  assign operator_6_false_23_acc_1_nl = nl_operator_6_false_23_acc_1_nl[5:0];
  assign nl_operator_6_false_27_acc_1_nl = ({1'b1 , (~ (rtn_out_1[5:1]))}) + 6'b000001;
  assign operator_6_false_27_acc_1_nl = nl_operator_6_false_27_acc_1_nl[5:0];
  assign nl_operator_6_false_46_acc_1_nl = ({1'b1 , (~ (leading_sign_57_0_1_0_20_out_3[5:1]))})
      + 6'b000001;
  assign operator_6_false_46_acc_1_nl = nl_operator_6_false_46_acc_1_nl[5:0];
  assign nl_operator_6_false_41_acc_1_nl = ({1'b1 , (~ (leading_sign_57_0_1_0_19_out_3[5:1]))})
      + 6'b000001;
  assign operator_6_false_41_acc_1_nl = nl_operator_6_false_41_acc_1_nl[5:0];
  assign operator_6_false_17_mux1h_12_nl = MUX1HOT_v_6_5_2(operator_6_false_17_acc_1_nl,
      operator_6_false_23_acc_1_nl, operator_6_false_27_acc_1_nl, operator_6_false_46_acc_1_nl,
      operator_6_false_41_acc_1_nl, {(fsm_output[12]) , (fsm_output[14]) , (fsm_output[16])
      , (fsm_output[28]) , (fsm_output[26])});
  assign operator_6_false_17_mux1h_13_nl = MUX1HOT_s_1_4_2((~ (rtn_out_1[0])), (~
      (leading_sign_57_0_1_0_10_out_3[0])), (~ (leading_sign_57_0_1_0_20_out_3[0])),
      (~ (leading_sign_57_0_1_0_19_out_3[0])), {return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse
      , (fsm_output[14]) , (fsm_output[28]) , (fsm_output[26])});
  assign nl_z_out_16 = conv_u2u_11_13({operator_6_false_17_mux1h_7_nl , operator_6_false_17_mux1h_8_nl
      , operator_6_false_17_mux1h_9_nl , operator_6_false_17_mux1h_10_nl , operator_6_false_17_mux1h_11_nl})
      + conv_s2u_7_13({operator_6_false_17_mux1h_12_nl , operator_6_false_17_mux1h_13_nl});
  assign z_out_16 = nl_z_out_16[12:0];
  assign return_add_generic_AC_RND_CONV_false_1_e_dif_qif_return_add_generic_AC_RND_CONV_false_1_e_dif_qif_mux_2_nl
      = MUX_v_11_2_2((out_f_d_rsci_q_d[62:52]), (in_f_d_rsci_q_d[62:52]), or_1266_cse);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif_qif_return_add_generic_AC_RND_CONV_false_1_e_dif_qif_mux_3_nl
      = MUX_v_11_2_2((~ (stage_PE_1_x_im_d_sva[62:52])), (~ (stage_PE_1_tmp_im_d_1_sva_1_63_51[11:1])),
      or_1495_cse_1);
  assign nl_acc_15_nl = ({1'b1 , return_add_generic_AC_RND_CONV_false_1_e_dif_qif_return_add_generic_AC_RND_CONV_false_1_e_dif_qif_mux_2_nl
      , 1'b1}) + conv_u2u_12_13({return_add_generic_AC_RND_CONV_false_1_e_dif_qif_return_add_generic_AC_RND_CONV_false_1_e_dif_qif_mux_3_nl
      , 1'b1});
  assign acc_15_nl = nl_acc_15_nl[12:0];
  assign z_out_17 = readslicef_13_12_1(acc_15_nl);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_return_add_generic_AC_RND_CONV_false_1_e_dif1_mux_2_nl
      = MUX_v_11_2_2((stage_PE_1_x_im_d_sva[62:52]), (stage_PE_1_tmp_im_d_1_sva_1_63_51[11:1]),
      or_1495_cse_1);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_return_add_generic_AC_RND_CONV_false_1_e_dif1_mux_3_nl
      = MUX_v_11_2_2((~ (out_f_d_rsci_q_d[62:52])), (~ (in_f_d_rsci_q_d[62:52])),
      or_1266_cse);
  assign nl_acc_16_nl = ({1'b1 , return_add_generic_AC_RND_CONV_false_1_e_dif1_return_add_generic_AC_RND_CONV_false_1_e_dif1_mux_2_nl
      , 1'b1}) + conv_u2u_12_13({return_add_generic_AC_RND_CONV_false_1_e_dif1_return_add_generic_AC_RND_CONV_false_1_e_dif1_mux_3_nl
      , 1'b1});
  assign acc_16_nl = nl_acc_16_nl[12:0];
  assign z_out_18 = readslicef_13_12_1(acc_16_nl);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_8_nl = MUX_s_1_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0,
      operator_6_false_18_acc_psp_sva_10_0_rsp_0, or_tmp_900);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_9_nl = MUX_v_9_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0,
      operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0, or_tmp_900);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_10_nl = MUX_s_1_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1,
      operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1, or_tmp_900);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_11_nl = MUX_s_1_2_2((~
      operator_6_false_18_acc_psp_sva_10_0_rsp_0), (~ reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0),
      or_tmp_900);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_12_nl = MUX_v_9_2_2((~
      operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0), (~ reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0),
      or_tmp_900);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_13_nl = MUX_s_1_2_2((~
      operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1), (~ reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1),
      or_tmp_900);
  assign nl_acc_17_nl = ({1'b1 , return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_8_nl
      , return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_9_nl , return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_10_nl
      , 1'b1}) + conv_u2u_12_13({return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_11_nl
      , return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_12_nl , return_add_generic_AC_RND_CONV_false_6_e_dif_qelse_mux_13_nl
      , 1'b1});
  assign acc_17_nl = nl_acc_17_nl[12:0];
  assign z_out_19 = readslicef_13_12_1(acc_17_nl);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_4_nl = MUX_v_10_2_2(stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_1,
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx1_10_1, fsm_output[25]);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_5_nl = MUX_s_1_2_2(stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0,
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx1_0, fsm_output[25]);
  assign nl_acc_18_nl = ({1'b1 , return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_4_nl
      , return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_5_nl , 1'b1}) + conv_u2u_12_13({(~
      operator_6_false_18_acc_psp_sva_10_0_rsp_0) , (~ operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0)
      , (~ operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1) , 1'b1});
  assign acc_18_nl = nl_acc_18_nl[12:0];
  assign z_out_20_11 = readslicef_13_1_12(acc_18_nl);
  assign nl_z_out_21 = conv_s2u_11_12(z_out_51[11:1]) + 12'b000000000001;
  assign z_out_21 = nl_z_out_21[11:0];
  assign operator_32_false_nor_2_nl = ~((fsm_output[11]) | (fsm_output[13]) | or_1367_cse);
  assign operator_32_false_operator_32_false_and_2_nl = MUX_v_6_2_2(6'b000000, (operator_32_false_2_mul_atp_sva_1[9:4]),
      operator_32_false_nor_2_nl);
  assign operator_32_false_mux_10_nl = MUX_v_2_2_2((in_u_rsc_merge_sva_rsp_0[5:4]),
      (operator_32_false_2_mul_atp_sva_1[3:2]), fsm_output[36]);
  assign operator_32_false_nor_3_nl = ~((fsm_output[13]) | or_1367_cse);
  assign operator_32_false_operator_32_false_and_3_nl = MUX_v_2_2_2(2'b00, operator_32_false_mux_10_nl,
      operator_32_false_nor_3_nl);
  assign operator_32_false_mux1h_11_nl = MUX1HOT_v_2_4_2((in_u_rsc_merge_sva_rsp_0[3:2]),
      (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd[2:1]), (in_u_rsci_q_d[15:14]),
      (operator_32_false_2_mul_atp_sva_1[1:0]), {(fsm_output[11]) , (fsm_output[13])
      , or_1367_cse , (fsm_output[36])});
  assign operator_32_false_mux1h_12_nl = MUX1HOT_s_1_3_2((in_u_rsc_merge_sva_rsp_0[1]),
      (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd[0]), (in_u_rsci_q_d[13]),
      {(fsm_output[11]) , (fsm_output[13]) , or_1367_cse});
  assign operator_32_false_and_5_nl = operator_32_false_mux1h_12_nl & (~ (fsm_output[36]));
  assign operator_32_false_mux1h_13_nl = MUX1HOT_s_1_3_2((in_u_rsc_merge_sva_rsp_0[0]),
      (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_2_1[1]), (in_u_rsci_q_d[12]),
      {(fsm_output[11]) , (fsm_output[13]) , or_1367_cse});
  assign operator_32_false_and_6_nl = operator_32_false_mux1h_13_nl & (~ (fsm_output[36]));
  assign operator_32_false_mux1h_14_nl = MUX1HOT_s_1_3_2((in_u_rsc_merge_sva_rsp_1_rsp_0[3]),
      (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_2_1[0]), (in_u_rsci_q_d[11]),
      {(fsm_output[11]) , (fsm_output[13]) , or_1367_cse});
  assign operator_32_false_and_7_nl = operator_32_false_mux1h_14_nl & (~ (fsm_output[36]));
  assign operator_32_false_mux1h_15_nl = MUX1HOT_s_1_3_2((in_u_rsc_merge_sva_rsp_1_rsp_0[2]),
      reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0, (in_u_rsci_q_d[10]),
      {(fsm_output[11]) , (fsm_output[13]) , or_1367_cse});
  assign operator_32_false_and_8_nl = operator_32_false_mux1h_15_nl & (~ (fsm_output[36]));
  assign operator_32_false_mux1h_16_nl = MUX1HOT_v_2_4_2((in_u_rsc_merge_sva_rsp_1_rsp_0[1:0]),
      (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0[8:7]), (in_u_rsci_q_d[9:8]),
      (operator_32_false_2_mul_atp_sva_1[9:8]), {(fsm_output[11]) , (fsm_output[13])
      , or_1367_cse , (fsm_output[36])});
  assign operator_32_false_mux1h_17_nl = MUX1HOT_v_6_4_2(in_u_rsc_merge_sva_rsp_1_rsp_1,
      (reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0[6:1]), (in_u_rsci_q_d[7:2]),
      (operator_32_false_2_mul_atp_sva_1[7:2]), {(fsm_output[11]) , (fsm_output[13])
      , or_1367_cse , (fsm_output[36])});
  assign operator_32_false_mux1h_18_nl = MUX1HOT_s_1_3_2((reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0[0]),
      (in_u_rsci_q_d[1]), (operator_32_false_2_mul_atp_sva_1[1]), {(fsm_output[13])
      , or_1367_cse , (fsm_output[36])});
  assign operator_32_false_and_9_nl = operator_32_false_mux1h_18_nl & (~ (fsm_output[11]));
  assign operator_32_false_mux1h_19_nl = MUX1HOT_s_1_3_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1,
      (in_u_rsci_q_d[0]), (operator_32_false_2_mul_atp_sva_1[0]), {(fsm_output[13])
      , or_1367_cse , (fsm_output[36])});
  assign operator_32_false_or_3_nl = operator_32_false_mux1h_19_nl | (fsm_output[11]);
  assign operator_32_false_or_4_nl = (fsm_output[11]) | stage_u_add_3_or_1_cse;
  assign operator_32_false_operator_32_false_or_4_nl = MUX_v_7_2_2((z_out_57[10:4]),
      7'b1111111, operator_32_false_or_4_nl);
  assign operator_32_false_mux1h_20_nl = MUX1HOT_v_4_3_2((z_out_1[15:12]), 4'b1100,
      (z_out_57[3:0]), {(fsm_output[11]) , stage_u_add_3_or_1_cse , (fsm_output[36])});
  assign operator_32_false_mux_11_nl = MUX_v_12_2_2((z_out_1[11:0]), (in_u_rsci_q_d[11:0]),
      fsm_output[36]);
  assign operator_32_false_operator_32_false_or_5_nl = MUX_v_12_2_2(operator_32_false_mux_11_nl,
      12'b111111111111, stage_u_add_3_or_1_cse);
  assign nl_z_out_22 = ({operator_32_false_operator_32_false_and_2_nl , operator_32_false_operator_32_false_and_3_nl
      , operator_32_false_mux1h_11_nl , operator_32_false_and_5_nl , operator_32_false_and_6_nl
      , operator_32_false_and_7_nl , operator_32_false_and_8_nl , operator_32_false_mux1h_16_nl
      , operator_32_false_mux1h_17_nl , operator_32_false_and_9_nl , operator_32_false_or_3_nl})
      + conv_s2u_23_24({operator_32_false_operator_32_false_or_4_nl , operator_32_false_mux1h_20_nl
      , operator_32_false_operator_32_false_or_5_nl});
  assign z_out_22 = nl_z_out_22[23:0];
  assign nl_z_out_23 = conv_s2u_17_18(z_out_28) + conv_u2u_14_18(signext_14_13({(z_out_28[16])
      , 11'b00000000000 , (z_out_28[16])}));
  assign z_out_23 = nl_z_out_23[17:0];
  assign return_mult_generic_AC_RND_CONV_false_2_exp_plus_1_mux_1_nl = MUX_v_12_2_2(return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_1,
      return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_1, fsm_output[27]);
  assign nl_z_out_24 = return_mult_generic_AC_RND_CONV_false_2_exp_plus_1_mux_1_nl
      + 12'b000000000001;
  assign z_out_24 = nl_z_out_24[11:0];
  assign BUTTERFLY_1_else_2_mux_5_nl = MUX_v_4_2_2((BUTTERFLY_1_if_mux_itm[13:10]),
      BUTTERFLY_mux_5_itm_13_10, fsm_output[10]);
  assign BUTTERFLY_1_else_2_mux_6_nl = MUX_v_10_2_2((BUTTERFLY_1_if_mux_itm[9:0]),
      BUTTERFLY_mux_5_itm_9_0, fsm_output[10]);
  assign BUTTERFLY_1_else_1_BUTTERFLY_1_else_1_and_1_nl = MUX_v_2_2_2(2'b00, (z_out_23[17:16]),
      inverse_lpi_1_dfm_1);
  assign BUTTERFLY_1_else_1_mux_9_nl = MUX_v_6_2_2(in_u_rsc_merge_sva_rsp_0, (z_out_23[15:10]),
      inverse_lpi_1_dfm_1);
  assign BUTTERFLY_1_else_1_mux_10_nl = MUX_v_4_2_2(in_u_rsc_merge_sva_rsp_1_rsp_0,
      (z_out_23[9:6]), inverse_lpi_1_dfm_1);
  assign BUTTERFLY_1_else_1_mux_11_nl = MUX_v_6_2_2(in_u_rsc_merge_sva_rsp_1_rsp_1,
      (z_out_23[5:0]), inverse_lpi_1_dfm_1);
  assign nl_z_out_25 = $signed(conv_u2s_14_15({BUTTERFLY_1_else_2_mux_5_nl , BUTTERFLY_1_else_2_mux_6_nl}))
      * $signed(({BUTTERFLY_1_else_1_BUTTERFLY_1_else_1_and_1_nl , BUTTERFLY_1_else_1_mux_9_nl
      , BUTTERFLY_1_else_1_mux_10_nl , BUTTERFLY_1_else_1_mux_11_nl}));
  assign z_out_25 = nl_z_out_25[31:0];
  assign BUTTERFLY_i_and_16_nl = BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm
      & (~ or_dcpl_83);
  assign BUTTERFLY_i_BUTTERFLY_i_mux_3_nl = MUX_s_1_2_2(stage_PE_1_tmp_im_d_1_lpi_3_dfm_51,
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_51, or_1556_cse);
  assign BUTTERFLY_i_and_17_nl = BUTTERFLY_i_BUTTERFLY_i_mux_3_nl & (~ or_dcpl_83);
  assign BUTTERFLY_i_mux_12_nl = MUX_v_42_2_2((stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0[50:9]),
      (stage_PE_1_tmp_im_d_1_sva_1_50_0[50:9]), or_1556_cse);
  assign not_898_nl = ~ or_dcpl_83;
  assign BUTTERFLY_i_BUTTERFLY_i_and_1_nl = MUX_v_42_2_2(42'b000000000000000000000000000000000000000000,
      BUTTERFLY_i_mux_12_nl, not_898_nl);
  assign BUTTERFLY_i_or_8_nl = (fsm_output[9]) | (fsm_output[24]);
  assign BUTTERFLY_i_mux1h_22_nl = MUX1HOT_v_9_3_2(BUTTERFLY_i_div_cmp_z_oreg, (stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0[8:0]),
      (stage_PE_1_tmp_im_d_1_sva_1_50_0[8:0]), {or_dcpl_83 , BUTTERFLY_i_or_8_nl
      , or_1556_cse});
  assign BUTTERFLY_i_mux1h_23_nl = MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm, return_extract_49_return_extract_49_or_sva_1,
      {(fsm_output[9]) , or_1556_cse , (fsm_output[24])});
  assign BUTTERFLY_i_and_18_nl = BUTTERFLY_i_mux1h_23_nl & (~ or_dcpl_83);
  assign BUTTERFLY_i_BUTTERFLY_i_mux_4_nl = MUX_s_1_2_2(drf_qr_lval_14_smx_0_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_17_m_r_51_lpi_3_dfm, or_1556_cse);
  assign BUTTERFLY_i_and_19_nl = BUTTERFLY_i_BUTTERFLY_i_mux_4_nl & (~ or_dcpl_83);
  assign BUTTERFLY_i_mux1h_24_nl = MUX1HOT_s_1_3_2((return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm[50]),
      (return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[50]), return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_50,
      {(fsm_output[9]) , or_1556_cse , (fsm_output[24])});
  assign BUTTERFLY_i_and_20_nl = BUTTERFLY_i_mux1h_24_nl & (~ or_dcpl_83);
  assign BUTTERFLY_i_mux1h_25_nl = MUX1HOT_v_40_3_2((return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm[49:10]),
      (return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[49:10]), (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0[49:10]),
      {(fsm_output[9]) , or_1556_cse , (fsm_output[24])});
  assign not_902_nl = ~ or_dcpl_83;
  assign BUTTERFLY_i_and_21_nl = MUX_v_40_2_2(40'b0000000000000000000000000000000000000000,
      BUTTERFLY_i_mux1h_25_nl, not_902_nl);
  assign BUTTERFLY_i_mux1h_26_nl = MUX1HOT_s_1_4_2(stage_PE_1_index_const_9_1_lpi_2_dfm_8,
      (return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm[9]), (return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[9]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0[9]), {or_dcpl_83
      , (fsm_output[9]) , or_1556_cse , (fsm_output[24])});
  assign BUTTERFLY_i_mux1h_27_nl = MUX1HOT_s_1_4_2(stage_PE_1_index_const_9_1_lpi_2_dfm_7,
      (return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm[8]), (return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[8]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0[8]), {or_dcpl_83
      , (fsm_output[9]) , or_1556_cse , (fsm_output[24])});
  assign BUTTERFLY_i_mux1h_28_nl = MUX1HOT_s_1_4_2(stage_PE_1_index_const_9_1_lpi_2_dfm_6,
      (return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm[7]), (return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[7]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0[7]), {or_dcpl_83
      , (fsm_output[9]) , or_1556_cse , (fsm_output[24])});
  assign BUTTERFLY_i_mux1h_29_nl = MUX1HOT_s_1_4_2(stage_PE_1_index_const_9_1_lpi_2_dfm_5,
      (return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm[6]), (return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[6]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0[6]), {or_dcpl_83
      , (fsm_output[9]) , or_1556_cse , (fsm_output[24])});
  assign BUTTERFLY_i_mux1h_30_nl = MUX1HOT_s_1_4_2(stage_PE_1_index_const_9_1_lpi_2_dfm_4,
      (return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm[5]), (return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[5]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0[5]), {or_dcpl_83
      , (fsm_output[9]) , or_1556_cse , (fsm_output[24])});
  assign BUTTERFLY_i_mux1h_31_nl = MUX1HOT_s_1_4_2(stage_PE_1_index_const_9_1_lpi_2_dfm_3,
      (return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm[4]), (return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[4]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0[4]), {or_dcpl_83
      , (fsm_output[9]) , or_1556_cse , (fsm_output[24])});
  assign BUTTERFLY_i_mux1h_32_nl = MUX1HOT_s_1_4_2(stage_PE_1_index_const_9_1_lpi_2_dfm_2,
      (return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm[3]), (return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[3]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0[3]), {or_dcpl_83
      , (fsm_output[9]) , or_1556_cse , (fsm_output[24])});
  assign BUTTERFLY_i_mux1h_33_nl = MUX1HOT_s_1_4_2(stage_PE_1_index_const_9_1_lpi_2_dfm_1,
      (return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm[2]), (return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[2]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0[2]), {or_dcpl_83
      , (fsm_output[9]) , or_1556_cse , (fsm_output[24])});
  assign BUTTERFLY_i_mux1h_34_nl = MUX1HOT_s_1_4_2(stage_PE_1_index_const_9_1_lpi_2_dfm_0,
      (return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm[1]), (return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[1]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0[1]), {or_dcpl_83
      , (fsm_output[9]) , or_1556_cse , (fsm_output[24])});
  assign BUTTERFLY_i_mux1h_35_nl = MUX1HOT_s_1_4_2(stage_PE_1_index_const_0_lpi_2_dfm,
      (return_mult_generic_AC_RND_CONV_false_3_if_mux_2_itm[0]), (return_add_generic_AC_RND_CONV_false_18_mux_1_itm_50_0[0]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm_1_49_0[0]), {or_dcpl_83
      , (fsm_output[9]) , or_1556_cse , (fsm_output[24])});
  assign z_out_26 = ({BUTTERFLY_i_and_16_nl , BUTTERFLY_i_and_17_nl , BUTTERFLY_i_BUTTERFLY_i_and_1_nl
      , BUTTERFLY_i_mux1h_22_nl}) * ({BUTTERFLY_i_and_18_nl , BUTTERFLY_i_and_19_nl
      , BUTTERFLY_i_and_20_nl , BUTTERFLY_i_and_21_nl , BUTTERFLY_i_mux1h_26_nl ,
      BUTTERFLY_i_mux1h_27_nl , BUTTERFLY_i_mux1h_28_nl , BUTTERFLY_i_mux1h_29_nl
      , BUTTERFLY_i_mux1h_30_nl , BUTTERFLY_i_mux1h_31_nl , BUTTERFLY_i_mux1h_32_nl
      , BUTTERFLY_i_mux1h_33_nl , BUTTERFLY_i_mux1h_34_nl , BUTTERFLY_i_mux1h_35_nl});
  assign BUTTERFLY_fry_mux_10_nl = MUX_s_1_2_2(stage_PE_1_qr_0_lpi_2_dfm, stage_PE_1_qr_10_1_lpi_2_dfm_8,
      or_tmp_920);
  assign BUTTERFLY_fry_mux_11_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_8, stage_PE_1_qr_10_1_lpi_2_dfm_7,
      or_tmp_920);
  assign BUTTERFLY_fry_mux_12_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_7, stage_PE_1_qr_10_1_lpi_2_dfm_6,
      or_tmp_920);
  assign BUTTERFLY_fry_mux_13_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_6, stage_PE_1_qr_10_1_lpi_2_dfm_5,
      or_tmp_920);
  assign BUTTERFLY_fry_mux_14_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_5, stage_PE_1_qr_10_1_lpi_2_dfm_4,
      or_tmp_920);
  assign BUTTERFLY_fry_mux_15_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_4, stage_PE_1_qr_10_1_lpi_2_dfm_3,
      or_tmp_920);
  assign BUTTERFLY_fry_mux_16_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_3, stage_PE_1_qr_10_1_lpi_2_dfm_2,
      or_tmp_920);
  assign BUTTERFLY_fry_mux_17_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_2, stage_PE_1_qr_10_1_lpi_2_dfm_1,
      or_tmp_920);
  assign BUTTERFLY_fry_mux_18_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_1, stage_PE_1_qr_10_1_lpi_2_dfm_0,
      or_tmp_920);
  assign BUTTERFLY_fry_mux_19_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_0, stage_PE_1_qr_0_lpi_2_dfm,
      or_tmp_920);
  assign nl_z_out_27 = BUTTERFLY_i_9_0_sva_1 + ({BUTTERFLY_fry_mux_10_nl , BUTTERFLY_fry_mux_11_nl
      , BUTTERFLY_fry_mux_12_nl , BUTTERFLY_fry_mux_13_nl , BUTTERFLY_fry_mux_14_nl
      , BUTTERFLY_fry_mux_15_nl , BUTTERFLY_fry_mux_16_nl , BUTTERFLY_fry_mux_17_nl
      , BUTTERFLY_fry_mux_18_nl , BUTTERFLY_fry_mux_19_nl});
  assign z_out_27 = nl_z_out_27[9:0];
  assign nl_acc_24_nl = ({1'b1 , BUTTERFLY_else_1_if_mux_4_cse , BUTTERFLY_else_1_if_mux_5_cse
      , BUTTERFLY_else_1_if_mux_6_cse , BUTTERFLY_else_1_if_mux_7_cse_9_1 , BUTTERFLY_else_1_if_mux_7_cse_0
      , 1'b1}) + conv_u2u_17_18({(~ in_u_rsc_merge_sva_rsp_0) , (~ in_u_rsc_merge_sva_rsp_1_rsp_0)
      , (~ in_u_rsc_merge_sva_rsp_1_rsp_1) , 1'b1});
  assign acc_24_nl = nl_acc_24_nl[17:0];
  assign z_out_28 = readslicef_18_17_1(acc_24_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_exp_acc_4_nl = conv_u2s_11_12({in_u_rsc_merge_sva_rsp_1_rsp_0
      , in_u_rsc_merge_sva_rsp_1_rsp_1 , return_add_generic_AC_RND_CONV_false_17_e_r_qelse_return_add_generic_AC_RND_CONV_false_17_e_r_qelse_and_1_itm})
      + conv_s2s_11_12({10'b1000000000 , (~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm)})
      + 12'b000000000001;
  assign return_mult_generic_AC_RND_CONV_false_exp_acc_4_nl = nl_return_mult_generic_AC_RND_CONV_false_exp_acc_4_nl[11:0];
  assign nl_return_mult_generic_AC_RND_CONV_false_4_exp_acc_2_nl = conv_u2s_11_12({return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1_9_1
      , return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1_0 , return_add_generic_AC_RND_CONV_false_18_e_r_qelse_return_add_generic_AC_RND_CONV_false_18_e_r_qelse_and_1_itm})
      + conv_s2s_11_12({10'b1000000000 , (~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm)})
      + 12'b000000000001;
  assign return_mult_generic_AC_RND_CONV_false_4_exp_acc_2_nl = nl_return_mult_generic_AC_RND_CONV_false_4_exp_acc_2_nl[11:0];
  assign return_mult_generic_AC_RND_CONV_false_3_exp_mux_5_nl = MUX_v_12_2_2(return_mult_generic_AC_RND_CONV_false_exp_acc_4_nl,
      return_mult_generic_AC_RND_CONV_false_4_exp_acc_2_nl, fsm_output[24]);
  assign return_mult_generic_AC_RND_CONV_false_3_exp_mux_6_nl = MUX_s_1_2_2(return_extract_15_return_extract_15_nor_cse_sva,
      return_extract_49_return_extract_49_nor_tmp, fsm_output[24]);
  assign return_mult_generic_AC_RND_CONV_false_3_exp_mux_7_nl = MUX_s_1_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_1_0,
      operator_6_false_18_acc_psp_sva_10_0_rsp_0, fsm_output[24]);
  assign return_mult_generic_AC_RND_CONV_false_3_exp_mux_8_nl = MUX_v_9_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0,
      operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_0, fsm_output[24]);
  assign return_mult_generic_AC_RND_CONV_false_3_exp_mux_9_nl = MUX_s_1_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1,
      operator_6_false_18_acc_psp_sva_10_0_rsp_1_rsp_1, fsm_output[24]);
  assign nl_acc_25_nl = conv_s2u_13_14({return_mult_generic_AC_RND_CONV_false_3_exp_mux_5_nl
      , return_mult_generic_AC_RND_CONV_false_3_exp_mux_6_nl}) + conv_u2u_12_14({return_mult_generic_AC_RND_CONV_false_3_exp_mux_7_nl
      , return_mult_generic_AC_RND_CONV_false_3_exp_mux_8_nl , return_mult_generic_AC_RND_CONV_false_3_exp_mux_9_nl
      , 1'b1});
  assign acc_25_nl = nl_acc_25_nl[13:0];
  assign z_out_45 = readslicef_14_13_1(acc_25_nl);
  assign return_add_generic_AC_RND_CONV_false_5_res_rounded_return_add_generic_AC_RND_CONV_false_5_res_rounded_mux_2_nl
      = MUX_v_53_2_2((z_out_37[56:4]), (z_out_39[56:4]), return_add_generic_AC_RND_CONV_false_5_res_rounded_or_1_cse);
  assign return_add_generic_AC_RND_CONV_false_5_res_rounded_and_1_nl = (z_out_37[3])
      & ((z_out_37[0]) | (z_out_37[1]) | (z_out_37[2]) | (z_out_37[4]));
  assign return_add_generic_AC_RND_CONV_false_5_res_rounded_return_add_generic_AC_RND_CONV_false_5_res_rounded_mux_3_nl
      = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_5_res_rounded_and_1_nl,
      return_add_generic_AC_RND_CONV_false_21_res_rounded_and_cse, return_add_generic_AC_RND_CONV_false_5_res_rounded_or_1_cse);
  assign nl_z_out_46 = conv_u2u_53_54(return_add_generic_AC_RND_CONV_false_5_res_rounded_return_add_generic_AC_RND_CONV_false_5_res_rounded_mux_2_nl)
      + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_5_res_rounded_return_add_generic_AC_RND_CONV_false_5_res_rounded_mux_3_nl);
  assign z_out_46 = nl_z_out_46[53:0];
  assign nl_z_out_47 = conv_u2u_53_54(z_out_36[56:4]) + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_1_res_rounded_and_1_cse);
  assign z_out_47 = nl_z_out_47[53:0];
  assign operator_6_false_25_mux_5_nl = MUX_v_14_2_2(({{8{operator_6_false_10_operator_6_false_10_conc_2_6_1[5]}},
      operator_6_false_10_operator_6_false_10_conc_2_6_1}), 14'b10011111111111, fsm_output[36]);
  assign operator_6_false_25_operator_6_false_25_or_1_nl = (~ (return_add_generic_AC_RND_CONV_false_20_ls_sva[0]))
      | (fsm_output[36]);
  assign operator_6_false_25_operator_6_false_25_and_1_nl = MUX_v_3_2_2(3'b000, (z_out_22[23:21]),
      (fsm_output[36]));
  assign operator_6_false_25_mux_6_nl = MUX_v_9_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_0,
      (z_out_22[20:12]), fsm_output[36]);
  assign operator_6_false_25_mux_7_nl = MUX_s_1_2_2(reg_BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_ftd_2_rsp_1,
      (z_out_22[11]), fsm_output[36]);
  assign operator_6_false_25_mux_8_nl = MUX_s_1_2_2(drf_qr_lval_14_smx_0_lpi_3_dfm,
      (z_out_22[10]), fsm_output[36]);
  assign nl_z_out_48 = ({operator_6_false_25_mux_5_nl , operator_6_false_25_operator_6_false_25_or_1_nl})
      + conv_u2u_14_15({operator_6_false_25_operator_6_false_25_and_1_nl , operator_6_false_25_mux_6_nl
      , operator_6_false_25_mux_7_nl , operator_6_false_25_mux_8_nl});
  assign z_out_48 = nl_z_out_48[14:0];
  assign BUTTERFLY_1_BUTTERFLY_1_and_3_nl = (BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[10])
      & BUTTERFLY_1_nor_1_cse;
  assign BUTTERFLY_1_mux_1548_nl = MUX_s_1_2_2((reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1[3]),
      (BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[9]), fsm_output[13]);
  assign BUTTERFLY_1_BUTTERFLY_1_and_4_nl = BUTTERFLY_1_mux_1548_nl & (~ or_tmp_1003);
  assign BUTTERFLY_1_mux1h_7_nl = MUX1HOT_v_3_3_2((operator_6_false_49_acc_psp_sva_8_0[8:6]),
      (reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1[2:0]), (BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[8:6]),
      {or_tmp_1003 , (fsm_output[8]) , (fsm_output[13])});
  assign BUTTERFLY_1_mux1h_8_nl = MUX1HOT_v_6_3_2((operator_6_false_49_acc_psp_sva_8_0[5:0]),
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2, (BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[5:0]),
      {or_tmp_1003 , (fsm_output[8]) , (fsm_output[13])});
  assign BUTTERFLY_1_or_1_nl = BUTTERFLY_1_nor_1_cse | (fsm_output[13]);
  assign BUTTERFLY_1_BUTTERFLY_1_or_2_nl = ((operator_6_false_8_operator_6_false_8_conc_itm_6_1[5])
      & (~ or_tmp_1003)) | (fsm_output[13]);
  assign BUTTERFLY_1_mux_1549_nl = MUX_v_5_2_2((operator_6_false_8_operator_6_false_8_conc_itm_6_1[4:0]),
      (~ (return_add_generic_AC_RND_CONV_false_20_ls_sva[5:1])), fsm_output[13]);
  assign not_905_nl = ~ or_tmp_1003;
  assign BUTTERFLY_1_BUTTERFLY_1_and_5_nl = MUX_v_5_2_2(5'b00000, BUTTERFLY_1_mux_1549_nl,
      not_905_nl);
  assign BUTTERFLY_1_mux_1550_nl = MUX_s_1_2_2((~ (return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_rsp_2[0])),
      (~ (return_add_generic_AC_RND_CONV_false_20_ls_sva[0])), fsm_output[13]);
  assign BUTTERFLY_1_BUTTERFLY_1_or_3_nl = BUTTERFLY_1_mux_1550_nl | or_tmp_1003;
  assign nl_acc_29_nl = conv_u2u_12_13({BUTTERFLY_1_BUTTERFLY_1_and_3_nl , BUTTERFLY_1_BUTTERFLY_1_and_4_nl
      , BUTTERFLY_1_mux1h_7_nl , BUTTERFLY_1_mux1h_8_nl , BUTTERFLY_1_or_1_nl}) +
      conv_s2u_8_13({BUTTERFLY_1_BUTTERFLY_1_or_2_nl , BUTTERFLY_1_BUTTERFLY_1_and_5_nl
      , BUTTERFLY_1_BUTTERFLY_1_or_3_nl , 1'b1});
  assign acc_29_nl = nl_acc_29_nl[12:0];
  assign z_out_49 = readslicef_13_12_1(acc_29_nl);
  assign operator_6_false_18_mux1h_22_nl = MUX1HOT_s_1_3_2(drf_qr_lval_10_smx_lpi_3_dfm_mx1_10,
      drf_qr_lval_6_smx_lpi_3_dfm_mx0_10, (drf_qr_lval_26_smx_lpi_3_dfm_mx0[10]),
      {(fsm_output[12]) , (fsm_output[26]) , (fsm_output[28])});
  assign operator_6_false_18_mux1h_23_nl = MUX1HOT_v_4_3_2(drf_qr_lval_10_smx_lpi_3_dfm_mx1_9_6,
      (drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_0[9:6]), (drf_qr_lval_26_smx_lpi_3_dfm_mx0[9:6]),
      {(fsm_output[12]) , (fsm_output[26]) , (fsm_output[28])});
  assign operator_6_false_18_mux1h_24_nl = MUX1HOT_v_6_3_2(drf_qr_lval_10_smx_lpi_3_dfm_mx1_5_0,
      (drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_0[5:0]), (drf_qr_lval_26_smx_lpi_3_dfm_mx0[5:0]),
      {(fsm_output[12]) , (fsm_output[26]) , (fsm_output[28])});
  assign operator_6_false_18_mux1h_25_nl = MUX1HOT_v_6_3_2((~ rtn_out_1), (~ leading_sign_57_0_1_0_19_out_3),
      (~ leading_sign_57_0_1_0_20_out_3), {(fsm_output[12]) , (fsm_output[26]) ,
      (fsm_output[28])});
  assign nl_acc_30_nl = conv_u2u_12_13({operator_6_false_18_mux1h_22_nl , operator_6_false_18_mux1h_23_nl
      , operator_6_false_18_mux1h_24_nl , 1'b1}) + conv_s2u_8_13({1'b1 , operator_6_false_18_mux1h_25_nl
      , 1'b1});
  assign acc_30_nl = nl_acc_30_nl[12:0];
  assign z_out_50 = readslicef_13_12_1(acc_30_nl);
  assign operator_6_false_3_mux1h_6_nl = MUX1HOT_v_4_3_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[10:7]),
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_1, (out_f_d_rsci_q_d[62:59]), {or_1531_cse
      , or_tmp_567 , (fsm_output[36])});
  assign operator_6_false_3_mux1h_7_nl = MUX1HOT_v_6_3_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[6:1]),
      reg_drf_qr_lval_10_smx_lpi_3_dfm_ftd_2, (out_f_d_rsci_q_d[58:53]), {or_1531_cse
      , or_tmp_567 , (fsm_output[36])});
  assign operator_6_false_3_mux1h_8_nl = MUX1HOT_s_1_3_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[0]),
      drf_qr_lval_12_smx_0_lpi_3_dfm, (out_f_d_rsci_q_d[52]), {or_1531_cse , or_tmp_567
      , (fsm_output[36])});
  assign operator_6_false_3_mux1h_9_nl = MUX1HOT_v_5_3_2((~ (leading_sign_57_0_1_0_2_out_3[5:1])),
      (~ (leading_sign_57_0_1_0_2_out_3[5:1])), 5'b11011, {or_1531_cse , or_tmp_567
      , (fsm_output[36])});
  assign operator_6_false_3_mux1h_10_nl = MUX1HOT_s_1_3_2((~ (leading_sign_57_0_1_0_2_out_3[0])),
      (~ (leading_sign_57_0_1_0_2_out_3[0])), (~ return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp),
      {or_1531_cse , or_tmp_567 , (fsm_output[36])});
  assign nl_acc_31_nl = conv_u2u_12_13({operator_6_false_3_mux1h_6_nl , operator_6_false_3_mux1h_7_nl
      , operator_6_false_3_mux1h_8_nl , 1'b1}) + conv_s2u_8_13({1'b1 , operator_6_false_3_mux1h_9_nl
      , operator_6_false_3_mux1h_10_nl , 1'b1});
  assign acc_31_nl = nl_acc_31_nl[12:0];
  assign z_out_51 = readslicef_13_12_1(acc_31_nl);
  assign operator_6_false_7_mux_5_nl = MUX_v_4_2_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[10:7]),
      in_u_rsc_merge_sva_rsp_1_rsp_0, fsm_output[30]);
  assign operator_6_false_7_mux_6_nl = MUX_v_6_2_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[6:1]),
      in_u_rsc_merge_sva_rsp_1_rsp_1, fsm_output[30]);
  assign operator_6_false_7_mux_7_nl = MUX_s_1_2_2((BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0[0]),
      return_add_generic_AC_RND_CONV_false_10_op1_mu_52_lpi_3_dfm, fsm_output[30]);
  assign operator_6_false_7_mux_8_nl = MUX_v_6_2_2((~ leading_sign_57_0_1_0_15_out_3),
      (~ leading_sign_57_0_1_0_25_out_3), fsm_output[30]);
  assign nl_acc_32_nl = conv_u2u_12_13({operator_6_false_7_mux_5_nl , operator_6_false_7_mux_6_nl
      , operator_6_false_7_mux_7_nl , 1'b1}) + conv_s2u_8_13({1'b1 , operator_6_false_7_mux_8_nl
      , 1'b1});
  assign acc_32_nl = nl_acc_32_nl[12:0];
  assign z_out_52 = readslicef_13_12_1(acc_32_nl);
  assign return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_mux_1_nl = MUX_v_2_2_2((return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_1[11:10]),
      (return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_1_cse[11:10]),
      return_mult_generic_AC_RND_CONV_false_1_else_1_or_cse);
  assign not_906_nl = ~ (fsm_output[37]);
  assign return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_and_1_nl
      = MUX_v_2_2_2(2'b00, return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_mux_1_nl,
      not_906_nl);
  assign return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_mux1h_2_nl = MUX1HOT_v_10_3_2((return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_1[9:0]),
      (return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_1_cse[9:0]),
      BUTTERFLY_1_fry_9_0_sva, {(fsm_output[9]) , return_mult_generic_AC_RND_CONV_false_1_else_1_or_cse
      , (fsm_output[37])});
  assign nl_z_out_55 = ({return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_and_1_nl
      , return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_mux1h_2_nl}) + 12'b000000000001;
  assign z_out_55 = nl_z_out_55[11:0];
  assign nl_z_out_56 = conv_s2u_11_12(z_out_13[11:1]) + 12'b000000000001;
  assign z_out_56 = nl_z_out_56[11:0];
  assign operator_6_false_15_not_1_nl = ~ (fsm_output[36]);
  assign operator_6_false_15_operator_6_false_15_and_1_nl = MUX_v_2_2_2(2'b00, (stage_u_add_3_acc_itm_rsp_1[12:11]),
      operator_6_false_15_not_1_nl);
  assign nl_operator_32_false_2_acc_7_nl = conv_u2u_10_11(~ operator_32_false_2_mul_atp_sva_1)
      + conv_u2u_4_11(in_u_rsci_q_d[15:12]);
  assign operator_32_false_2_acc_7_nl = nl_operator_32_false_2_acc_7_nl[10:0];
  assign operator_6_false_15_mux_3_nl = MUX_v_11_2_2((stage_u_add_3_acc_itm_rsp_1[10:0]),
      operator_32_false_2_acc_7_nl, fsm_output[36]);
  assign operator_6_false_15_or_1_nl = (~ (fsm_output[36])) | (fsm_output[9]);
  assign operator_6_false_15_mux_4_nl = MUX_v_6_2_2((~ return_add_generic_AC_RND_CONV_false_20_ls_sva),
      6'b000001, fsm_output[36]);
  assign nl_acc_35_nl = ({operator_6_false_15_operator_6_false_15_and_1_nl , operator_6_false_15_mux_3_nl
      , operator_6_false_15_or_1_nl}) + conv_s2u_12_14({1'b1 , (~ (fsm_output[36]))
      , (~ (fsm_output[36])) , (~ (fsm_output[36])) , (~ (fsm_output[36])) , operator_6_false_15_mux_4_nl
      , 1'b1});
  assign acc_35_nl = nl_acc_35_nl[13:0];
  assign z_out_57 = readslicef_14_13_1(acc_35_nl);
  assign BUTTERFLY_else_2_mux_5_nl = MUX_v_4_2_2(stage_u_add_3_acc_itm_rsp_0, (z_out_1[16:13]),
      fsm_output[24]);
  assign BUTTERFLY_else_2_mux_6_nl = MUX_v_13_2_2(stage_u_add_3_acc_itm_rsp_1, (z_out_1[12:0]),
      fsm_output[24]);
  assign nl_z_out_58 = ({BUTTERFLY_else_2_mux_5_nl , BUTTERFLY_else_2_mux_6_nl})
      + conv_u2u_14_17(signext_14_13({BUTTERFLY_else_2_mux_1_cse , 11'b00000000000
      , BUTTERFLY_else_2_mux_1_cse}));
  assign z_out_58 = nl_z_out_58[16:0];
  assign BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_3_nl = MUX_v_16_2_2((z_out_60[15:0]),
      (z_out_61[15:0]), or_dcpl_551);
  assign nl_z_out_59 = BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_3_nl +
      conv_u2u_14_16(signext_14_13({BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_1_cse
      , 11'b00000000000 , BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_1_cse}));
  assign z_out_59 = nl_z_out_59[15:0];
  assign stage_u_add_3_mux_2_nl = MUX_v_6_2_2(BUTTERFLY_else_2_acc_1_psp_16_0_sva_16_11,
      (z_out_58[16:11]), fsm_output[24]);
  assign stage_u_add_3_mux_3_nl = MUX_v_11_2_2(BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0,
      (z_out_58[10:0]), fsm_output[24]);
  assign nl_z_out_60 = conv_s2u_17_18({stage_u_add_3_acc_itm_rsp_0 , stage_u_add_3_acc_itm_rsp_1})
      + conv_s2u_17_18({stage_u_add_3_mux_2_nl , stage_u_add_3_mux_3_nl});
  assign z_out_60 = nl_z_out_60[17:0];
  assign stage_u_add_mux_5_nl = MUX_v_4_2_2(stage_u_add_3_acc_itm_rsp_0, (~ (BUTTERFLY_else_2_acc_1_psp_16_0_sva_16_11[5:2])),
      fsm_output[15]);
  assign stage_u_add_mux_6_nl = MUX_v_2_2_2((stage_u_add_3_acc_itm_rsp_1[12:11]),
      (~ (BUTTERFLY_else_2_acc_1_psp_16_0_sva_16_11[1:0])), fsm_output[15]);
  assign stage_u_add_mux_7_nl = MUX_v_11_2_2((stage_u_add_3_acc_itm_rsp_1[10:0]),
      (~ BUTTERFLY_else_2_acc_1_psp_16_0_sva_10_0), fsm_output[15]);
  assign stage_u_add_or_5_nl = (~((fsm_output[9]) | (fsm_output[22]))) | (fsm_output[15]);
  assign nl_acc_39_nl = conv_s2u_18_19({stage_u_add_mux_5_nl , stage_u_add_mux_6_nl
      , stage_u_add_mux_7_nl , stage_u_add_or_5_nl}) + conv_u2u_17_19({BUTTERFLY_else_1_if_mux_4_cse
      , BUTTERFLY_else_1_if_mux_5_cse , BUTTERFLY_else_1_if_mux_6_cse , BUTTERFLY_else_1_if_mux_7_cse_9_1
      , BUTTERFLY_else_1_if_mux_7_cse_0 , 1'b1});
  assign acc_39_nl = nl_acc_39_nl[18:0];
  assign z_out_61 = readslicef_19_18_1(acc_39_nl);
  assign operator_6_false_43_mux_3_nl = MUX_v_6_2_2((~ leading_sign_53_0_out_1),
      (~ leading_sign_53_0_4_out_1), fsm_output[24]);
  assign nl_acc_41_nl = ({z_out_45 , 1'b1}) + conv_s2u_8_14({1'b1 , operator_6_false_43_mux_3_nl
      , 1'b1});
  assign acc_41_nl = nl_acc_41_nl[13:0];
  assign z_out_63 = readslicef_14_13_1(acc_41_nl);
  assign nl_operator_32_false_1_acc_8_nl = conv_u2s_4_16(operator_32_false_1_mul_atp_sva_1[15:12])
      + (~ operator_32_false_1_mul_atp_sva_1);
  assign operator_32_false_1_acc_8_nl = nl_operator_32_false_1_acc_8_nl[15:0];
  assign nl_operator_32_false_1_acc_7_nl = ({operator_32_false_1_mul_atp_sva_1 ,
      2'b01}) + conv_s2u_17_18({1'b1 , operator_32_false_1_acc_8_nl});
  assign operator_32_false_1_acc_7_nl = nl_operator_32_false_1_acc_7_nl[17:0];
  assign operator_32_false_1_mux_4_nl = MUX_v_18_2_2(operator_32_false_1_acc_7_nl,
      (z_out_22[17:0]), fsm_output[11]);
  assign operator_32_false_1_mux_5_nl = MUX_v_2_2_2((operator_32_false_1_mul_atp_sva_1[11:10]),
      (in_u_rsc_merge_sva_rsp_0[1:0]), fsm_output[11]);
  assign operator_32_false_1_mux_6_nl = MUX_v_4_2_2((operator_32_false_1_mul_atp_sva_1[9:6]),
      in_u_rsc_merge_sva_rsp_1_rsp_0, fsm_output[11]);
  assign operator_32_false_1_mux_7_nl = MUX_v_6_2_2((operator_32_false_1_mul_atp_sva_1[5:0]),
      in_u_rsc_merge_sva_rsp_1_rsp_1, fsm_output[11]);
  assign nl_operator_32_false_1_acc_nl_1 = BUTTERFLY_1_else_2_tmp2_1_sva + conv_u2u_30_32({operator_32_false_1_mux_4_nl
      , operator_32_false_1_mux_5_nl , operator_32_false_1_mux_6_nl , operator_32_false_1_mux_7_nl});
  assign operator_32_false_1_acc_nl_1 = nl_operator_32_false_1_acc_nl_1[31:0];
  assign z_out_64_31_16 = readslicef_32_16_16(operator_32_false_1_acc_nl_1);
  assign return_add_generic_AC_RND_CONV_false_8_op_bigger_mux_6_nl = MUX_s_1_2_2(or_451_cse,
      return_add_generic_AC_RND_CONV_false_21_op1_smaller_lor_lpi_3_dfm_2, fsm_output[28]);
  assign z_out_10 = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_50_1_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_8_op_bigger_mux_6_nl);
  assign return_add_generic_AC_RND_CONV_false_7_mux_47_nl = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_7_res_rounded_acc_tmp[53]),
      (return_add_generic_AC_RND_CONV_false_20_res_rounded_acc_tmp[53]), fsm_output[29]);
  assign z_out_44 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_and_9,
      (return_add_generic_AC_RND_CONV_false_7_exp_plus_1_12_1_lpi_3_dfm_1[9:0]),
      return_add_generic_AC_RND_CONV_false_7_mux_47_nl);
  assign return_mult_generic_AC_RND_CONV_false_1_return_mult_generic_AC_RND_CONV_false_1_nor_1_nl
      = ~(return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_tmp_1 | (stage_u_add_3_acc_itm_rsp_1[12]));
  assign return_mult_generic_AC_RND_CONV_false_2_return_mult_generic_AC_RND_CONV_false_2_nor_1_nl
      = ~(return_mult_generic_AC_RND_CONV_false_2_if_1_and_1_tmp_1 | (return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp[12]));
  assign return_mult_generic_AC_RND_CONV_false_5_return_mult_generic_AC_RND_CONV_false_5_nor_1_nl
      = ~(return_mult_generic_AC_RND_CONV_false_5_if_1_and_1_tmp_1 | (return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp[12]));
  assign return_mult_generic_AC_RND_CONV_false_1_mux1h_8_m1c = MUX1HOT_s_1_3_2(return_mult_generic_AC_RND_CONV_false_1_return_mult_generic_AC_RND_CONV_false_1_nor_1_nl,
      return_mult_generic_AC_RND_CONV_false_2_return_mult_generic_AC_RND_CONV_false_2_nor_1_nl,
      return_mult_generic_AC_RND_CONV_false_5_return_mult_generic_AC_RND_CONV_false_5_nor_1_nl,
      {(fsm_output[9]) , (fsm_output[11]) , (fsm_output[27])});
  assign return_mult_generic_AC_RND_CONV_false_1_and_5_nl = return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_tmp_1
      & (~ (stage_u_add_3_acc_itm_rsp_1[12]));
  assign return_mult_generic_AC_RND_CONV_false_2_and_3_nl = return_mult_generic_AC_RND_CONV_false_2_if_1_and_1_tmp_1
      & (~ (return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp[12]));
  assign return_mult_generic_AC_RND_CONV_false_5_and_3_nl = return_mult_generic_AC_RND_CONV_false_5_if_1_and_1_tmp_1
      & (~ (return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp[12]));
  assign return_mult_generic_AC_RND_CONV_false_1_mux1h_9_m1c = MUX1HOT_s_1_3_2(return_mult_generic_AC_RND_CONV_false_1_and_5_nl,
      return_mult_generic_AC_RND_CONV_false_2_and_3_nl, return_mult_generic_AC_RND_CONV_false_5_and_3_nl,
      {(fsm_output[9]) , (fsm_output[11]) , (fsm_output[27])});
  assign return_mult_generic_AC_RND_CONV_false_1_mux1h_10_m1c = MUX1HOT_s_1_3_2((stage_u_add_3_acc_itm_rsp_1[12]),
      (return_mult_generic_AC_RND_CONV_false_2_exp_acc_tmp[12]), (return_mult_generic_AC_RND_CONV_false_5_exp_acc_tmp[12]),
      {(fsm_output[9]) , (fsm_output[11]) , (fsm_output[27])});
  assign return_mult_generic_AC_RND_CONV_false_1_and_nl = (fsm_output[9]) & return_mult_generic_AC_RND_CONV_false_1_mux1h_8_m1c;
  assign return_mult_generic_AC_RND_CONV_false_1_and_6_nl = (fsm_output[11]) & return_mult_generic_AC_RND_CONV_false_1_mux1h_8_m1c;
  assign return_mult_generic_AC_RND_CONV_false_1_and_7_nl = (fsm_output[27]) & return_mult_generic_AC_RND_CONV_false_1_mux1h_8_m1c;
  assign return_mult_generic_AC_RND_CONV_false_1_and_8_nl = (fsm_output[9]) & return_mult_generic_AC_RND_CONV_false_1_mux1h_9_m1c;
  assign return_mult_generic_AC_RND_CONV_false_1_and_9_nl = (fsm_output[11]) & return_mult_generic_AC_RND_CONV_false_1_mux1h_9_m1c;
  assign return_mult_generic_AC_RND_CONV_false_1_and_10_nl = (fsm_output[27]) & return_mult_generic_AC_RND_CONV_false_1_mux1h_9_m1c;
  assign return_mult_generic_AC_RND_CONV_false_1_and_11_nl = (~ or_dcpl_338) & return_mult_generic_AC_RND_CONV_false_1_mux1h_10_m1c;
  assign return_mult_generic_AC_RND_CONV_false_1_and_12_nl = or_dcpl_338 & return_mult_generic_AC_RND_CONV_false_1_mux1h_10_m1c;
  assign z_out_53 = MUX1HOT_v_53_8_2((z_out_54[104:52]), (return_mult_generic_AC_RND_CONV_false_2_p_sva_1[104:52]),
      (return_mult_generic_AC_RND_CONV_false_5_p_sva_1[104:52]), (z_out_54[103:51]),
      (return_mult_generic_AC_RND_CONV_false_2_p_sva_1[103:51]), (return_mult_generic_AC_RND_CONV_false_5_p_sva_1[103:51]),
      (z_out_35[53:1]), (z_out_34[53:1]), {return_mult_generic_AC_RND_CONV_false_1_and_nl
      , return_mult_generic_AC_RND_CONV_false_1_and_6_nl , return_mult_generic_AC_RND_CONV_false_1_and_7_nl
      , return_mult_generic_AC_RND_CONV_false_1_and_8_nl , return_mult_generic_AC_RND_CONV_false_1_and_9_nl
      , return_mult_generic_AC_RND_CONV_false_1_and_10_nl , return_mult_generic_AC_RND_CONV_false_1_and_11_nl
      , return_mult_generic_AC_RND_CONV_false_1_and_12_nl});

  function automatic  MUX1HOT_s_1_10_2;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [9:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    MUX1HOT_s_1_10_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_11_2;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [10:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    MUX1HOT_s_1_11_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_12_2;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [11:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    MUX1HOT_s_1_12_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_13_2;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [12:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    MUX1HOT_s_1_13_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_15_2;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [14:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    MUX1HOT_s_1_15_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_16_2;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [15:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    MUX1HOT_s_1_16_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_5_2;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [4:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_6_2;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [5:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_7_2;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [6:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_8_2;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [7:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    MUX1HOT_s_1_8_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_9_2;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [8:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    MUX1HOT_s_1_9_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_10_2;
    input [9:0] input_9;
    input [9:0] input_8;
    input [9:0] input_7;
    input [9:0] input_6;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [9:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    result = result | (input_3 & {10{sel[3]}});
    result = result | (input_4 & {10{sel[4]}});
    result = result | (input_5 & {10{sel[5]}});
    result = result | (input_6 & {10{sel[6]}});
    result = result | (input_7 & {10{sel[7]}});
    result = result | (input_8 & {10{sel[8]}});
    result = result | (input_9 & {10{sel[9]}});
    MUX1HOT_v_10_10_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_3_2;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [2:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    MUX1HOT_v_10_3_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_4_2;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [3:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    result = result | (input_3 & {10{sel[3]}});
    MUX1HOT_v_10_4_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_5_2;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [4:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    result = result | (input_3 & {10{sel[3]}});
    result = result | (input_4 & {10{sel[4]}});
    MUX1HOT_v_10_5_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_6_2;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [5:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    result = result | (input_3 & {10{sel[3]}});
    result = result | (input_4 & {10{sel[4]}});
    result = result | (input_5 & {10{sel[5]}});
    MUX1HOT_v_10_6_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_9_2;
    input [9:0] input_8;
    input [9:0] input_7;
    input [9:0] input_6;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [8:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    result = result | (input_3 & {10{sel[3]}});
    result = result | (input_4 & {10{sel[4]}});
    result = result | (input_5 & {10{sel[5]}});
    result = result | (input_6 & {10{sel[6]}});
    result = result | (input_7 & {10{sel[7]}});
    result = result | (input_8 & {10{sel[8]}});
    MUX1HOT_v_10_9_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_3_2;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [2:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    MUX1HOT_v_11_3_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_8_2;
    input [10:0] input_7;
    input [10:0] input_6;
    input [10:0] input_5;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [7:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    result = result | (input_3 & {11{sel[3]}});
    result = result | (input_4 & {11{sel[4]}});
    result = result | (input_5 & {11{sel[5]}});
    result = result | (input_6 & {11{sel[6]}});
    result = result | (input_7 & {11{sel[7]}});
    MUX1HOT_v_11_8_2 = result;
  end
  endfunction


  function automatic [12:0] MUX1HOT_v_13_7_2;
    input [12:0] input_6;
    input [12:0] input_5;
    input [12:0] input_4;
    input [12:0] input_3;
    input [12:0] input_2;
    input [12:0] input_1;
    input [12:0] input_0;
    input [6:0] sel;
    reg [12:0] result;
  begin
    result = input_0 & {13{sel[0]}};
    result = result | (input_1 & {13{sel[1]}});
    result = result | (input_2 & {13{sel[2]}});
    result = result | (input_3 & {13{sel[3]}});
    result = result | (input_4 & {13{sel[4]}});
    result = result | (input_5 & {13{sel[5]}});
    result = result | (input_6 & {13{sel[6]}});
    MUX1HOT_v_13_7_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_5_2;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [4:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    MUX1HOT_v_2_5_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_6_2;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [5:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    MUX1HOT_v_2_6_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_5_2;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [4:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    MUX1HOT_v_3_5_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_6_2;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [5:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    result = result | (input_5 & {3{sel[5]}});
    MUX1HOT_v_3_6_2 = result;
  end
  endfunction


  function automatic [39:0] MUX1HOT_v_40_3_2;
    input [39:0] input_2;
    input [39:0] input_1;
    input [39:0] input_0;
    input [2:0] sel;
    reg [39:0] result;
  begin
    result = input_0 & {40{sel[0]}};
    result = result | (input_1 & {40{sel[1]}});
    result = result | (input_2 & {40{sel[2]}});
    MUX1HOT_v_40_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_10_2;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [9:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    MUX1HOT_v_4_10_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_11_2;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [10:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    MUX1HOT_v_4_11_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_5_2;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [4:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    MUX1HOT_v_4_5_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_8_2;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [7:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    MUX1HOT_v_4_8_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_9_2;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [8:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    MUX1HOT_v_4_9_2 = result;
  end
  endfunction


  function automatic [49:0] MUX1HOT_v_50_14_2;
    input [49:0] input_13;
    input [49:0] input_12;
    input [49:0] input_11;
    input [49:0] input_10;
    input [49:0] input_9;
    input [49:0] input_8;
    input [49:0] input_7;
    input [49:0] input_6;
    input [49:0] input_5;
    input [49:0] input_4;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [13:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    result = result | (input_3 & {50{sel[3]}});
    result = result | (input_4 & {50{sel[4]}});
    result = result | (input_5 & {50{sel[5]}});
    result = result | (input_6 & {50{sel[6]}});
    result = result | (input_7 & {50{sel[7]}});
    result = result | (input_8 & {50{sel[8]}});
    result = result | (input_9 & {50{sel[9]}});
    result = result | (input_10 & {50{sel[10]}});
    result = result | (input_11 & {50{sel[11]}});
    result = result | (input_12 & {50{sel[12]}});
    result = result | (input_13 & {50{sel[13]}});
    MUX1HOT_v_50_14_2 = result;
  end
  endfunction


  function automatic [49:0] MUX1HOT_v_50_3_2;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [2:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    MUX1HOT_v_50_3_2 = result;
  end
  endfunction


  function automatic [49:0] MUX1HOT_v_50_4_2;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [3:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    result = result | (input_3 & {50{sel[3]}});
    MUX1HOT_v_50_4_2 = result;
  end
  endfunction


  function automatic [49:0] MUX1HOT_v_50_5_2;
    input [49:0] input_4;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [4:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    result = result | (input_3 & {50{sel[3]}});
    result = result | (input_4 & {50{sel[4]}});
    MUX1HOT_v_50_5_2 = result;
  end
  endfunction


  function automatic [49:0] MUX1HOT_v_50_6_2;
    input [49:0] input_5;
    input [49:0] input_4;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [5:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    result = result | (input_3 & {50{sel[3]}});
    result = result | (input_4 & {50{sel[4]}});
    result = result | (input_5 & {50{sel[5]}});
    MUX1HOT_v_50_6_2 = result;
  end
  endfunction


  function automatic [49:0] MUX1HOT_v_50_8_2;
    input [49:0] input_7;
    input [49:0] input_6;
    input [49:0] input_5;
    input [49:0] input_4;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [7:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    result = result | (input_3 & {50{sel[3]}});
    result = result | (input_4 & {50{sel[4]}});
    result = result | (input_5 & {50{sel[5]}});
    result = result | (input_6 & {50{sel[6]}});
    result = result | (input_7 & {50{sel[7]}});
    MUX1HOT_v_50_8_2 = result;
  end
  endfunction


  function automatic [50:0] MUX1HOT_v_51_11_2;
    input [50:0] input_10;
    input [50:0] input_9;
    input [50:0] input_8;
    input [50:0] input_7;
    input [50:0] input_6;
    input [50:0] input_5;
    input [50:0] input_4;
    input [50:0] input_3;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [10:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | (input_1 & {51{sel[1]}});
    result = result | (input_2 & {51{sel[2]}});
    result = result | (input_3 & {51{sel[3]}});
    result = result | (input_4 & {51{sel[4]}});
    result = result | (input_5 & {51{sel[5]}});
    result = result | (input_6 & {51{sel[6]}});
    result = result | (input_7 & {51{sel[7]}});
    result = result | (input_8 & {51{sel[8]}});
    result = result | (input_9 & {51{sel[9]}});
    result = result | (input_10 & {51{sel[10]}});
    MUX1HOT_v_51_11_2 = result;
  end
  endfunction


  function automatic [50:0] MUX1HOT_v_51_3_2;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [2:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | (input_1 & {51{sel[1]}});
    result = result | (input_2 & {51{sel[2]}});
    MUX1HOT_v_51_3_2 = result;
  end
  endfunction


  function automatic [50:0] MUX1HOT_v_51_4_2;
    input [50:0] input_3;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [3:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | (input_1 & {51{sel[1]}});
    result = result | (input_2 & {51{sel[2]}});
    result = result | (input_3 & {51{sel[3]}});
    MUX1HOT_v_51_4_2 = result;
  end
  endfunction


  function automatic [50:0] MUX1HOT_v_51_6_2;
    input [50:0] input_5;
    input [50:0] input_4;
    input [50:0] input_3;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [5:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | (input_1 & {51{sel[1]}});
    result = result | (input_2 & {51{sel[2]}});
    result = result | (input_3 & {51{sel[3]}});
    result = result | (input_4 & {51{sel[4]}});
    result = result | (input_5 & {51{sel[5]}});
    MUX1HOT_v_51_6_2 = result;
  end
  endfunction


  function automatic [50:0] MUX1HOT_v_51_7_2;
    input [50:0] input_6;
    input [50:0] input_5;
    input [50:0] input_4;
    input [50:0] input_3;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [6:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | (input_1 & {51{sel[1]}});
    result = result | (input_2 & {51{sel[2]}});
    result = result | (input_3 & {51{sel[3]}});
    result = result | (input_4 & {51{sel[4]}});
    result = result | (input_5 & {51{sel[5]}});
    result = result | (input_6 & {51{sel[6]}});
    MUX1HOT_v_51_7_2 = result;
  end
  endfunction


  function automatic [51:0] MUX1HOT_v_52_3_2;
    input [51:0] input_2;
    input [51:0] input_1;
    input [51:0] input_0;
    input [2:0] sel;
    reg [51:0] result;
  begin
    result = input_0 & {52{sel[0]}};
    result = result | (input_1 & {52{sel[1]}});
    result = result | (input_2 & {52{sel[2]}});
    MUX1HOT_v_52_3_2 = result;
  end
  endfunction


  function automatic [52:0] MUX1HOT_v_53_3_2;
    input [52:0] input_2;
    input [52:0] input_1;
    input [52:0] input_0;
    input [2:0] sel;
    reg [52:0] result;
  begin
    result = input_0 & {53{sel[0]}};
    result = result | (input_1 & {53{sel[1]}});
    result = result | (input_2 & {53{sel[2]}});
    MUX1HOT_v_53_3_2 = result;
  end
  endfunction


  function automatic [52:0] MUX1HOT_v_53_8_2;
    input [52:0] input_7;
    input [52:0] input_6;
    input [52:0] input_5;
    input [52:0] input_4;
    input [52:0] input_3;
    input [52:0] input_2;
    input [52:0] input_1;
    input [52:0] input_0;
    input [7:0] sel;
    reg [52:0] result;
  begin
    result = input_0 & {53{sel[0]}};
    result = result | (input_1 & {53{sel[1]}});
    result = result | (input_2 & {53{sel[2]}});
    result = result | (input_3 & {53{sel[3]}});
    result = result | (input_4 & {53{sel[4]}});
    result = result | (input_5 & {53{sel[5]}});
    result = result | (input_6 & {53{sel[6]}});
    result = result | (input_7 & {53{sel[7]}});
    MUX1HOT_v_53_8_2 = result;
  end
  endfunction


  function automatic [55:0] MUX1HOT_v_56_4_2;
    input [55:0] input_3;
    input [55:0] input_2;
    input [55:0] input_1;
    input [55:0] input_0;
    input [3:0] sel;
    reg [55:0] result;
  begin
    result = input_0 & {56{sel[0]}};
    result = result | (input_1 & {56{sel[1]}});
    result = result | (input_2 & {56{sel[2]}});
    result = result | (input_3 & {56{sel[3]}});
    MUX1HOT_v_56_4_2 = result;
  end
  endfunction


  function automatic [56:0] MUX1HOT_v_57_3_2;
    input [56:0] input_2;
    input [56:0] input_1;
    input [56:0] input_0;
    input [2:0] sel;
    reg [56:0] result;
  begin
    result = input_0 & {57{sel[0]}};
    result = result | (input_1 & {57{sel[1]}});
    result = result | (input_2 & {57{sel[2]}});
    MUX1HOT_v_57_3_2 = result;
  end
  endfunction


  function automatic [56:0] MUX1HOT_v_57_5_2;
    input [56:0] input_4;
    input [56:0] input_3;
    input [56:0] input_2;
    input [56:0] input_1;
    input [56:0] input_0;
    input [4:0] sel;
    reg [56:0] result;
  begin
    result = input_0 & {57{sel[0]}};
    result = result | (input_1 & {57{sel[1]}});
    result = result | (input_2 & {57{sel[2]}});
    result = result | (input_3 & {57{sel[3]}});
    result = result | (input_4 & {57{sel[4]}});
    MUX1HOT_v_57_5_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_4_2;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [3:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    MUX1HOT_v_5_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_5_2;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [4:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    MUX1HOT_v_5_5_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_6_2;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [5:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    MUX1HOT_v_5_6_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_11_2;
    input [5:0] input_10;
    input [5:0] input_9;
    input [5:0] input_8;
    input [5:0] input_7;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [10:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    result = result | (input_6 & {6{sel[6]}});
    result = result | (input_7 & {6{sel[7]}});
    result = result | (input_8 & {6{sel[8]}});
    result = result | (input_9 & {6{sel[9]}});
    result = result | (input_10 & {6{sel[10]}});
    MUX1HOT_v_6_11_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_5_2;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [4:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    MUX1HOT_v_6_5_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_6_2;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [5:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    MUX1HOT_v_6_6_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_9_2;
    input [5:0] input_8;
    input [5:0] input_7;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [8:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    result = result | (input_6 & {6{sel[6]}});
    result = result | (input_7 & {6{sel[7]}});
    result = result | (input_8 & {6{sel[8]}});
    MUX1HOT_v_6_9_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_3_2;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [2:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | (input_1 & {9{sel[1]}});
    result = result | (input_2 & {9{sel[2]}});
    MUX1HOT_v_9_3_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_5_2;
    input [8:0] input_4;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [4:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | (input_1 & {9{sel[1]}});
    result = result | (input_2 & {9{sel[2]}});
    result = result | (input_3 & {9{sel[3]}});
    result = result | (input_4 & {9{sel[4]}});
    MUX1HOT_v_9_5_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_8_2;
    input [8:0] input_7;
    input [8:0] input_6;
    input [8:0] input_5;
    input [8:0] input_4;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [7:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | (input_1 & {9{sel[1]}});
    result = result | (input_2 & {9{sel[2]}});
    result = result | (input_3 & {9{sel[3]}});
    result = result | (input_4 & {9{sel[4]}});
    result = result | (input_5 & {9{sel[5]}});
    result = result | (input_6 & {9{sel[6]}});
    result = result | (input_7 & {9{sel[7]}});
    MUX1HOT_v_9_8_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input  sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input  sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [12:0] MUX_v_13_2_2;
    input [12:0] input_0;
    input [12:0] input_1;
    input  sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input  sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [17:0] MUX_v_18_2_2;
    input [17:0] input_0;
    input [17:0] input_1;
    input  sel;
    reg [17:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_18_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [39:0] MUX_v_40_2_2;
    input [39:0] input_0;
    input [39:0] input_1;
    input  sel;
    reg [39:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_40_2_2 = result;
  end
  endfunction


  function automatic [41:0] MUX_v_42_2_2;
    input [41:0] input_0;
    input [41:0] input_1;
    input  sel;
    reg [41:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_42_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [49:0] MUX_v_50_2_2;
    input [49:0] input_0;
    input [49:0] input_1;
    input  sel;
    reg [49:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_50_2_2 = result;
  end
  endfunction


  function automatic [50:0] MUX_v_51_2_2;
    input [50:0] input_0;
    input [50:0] input_1;
    input  sel;
    reg [50:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_51_2_2 = result;
  end
  endfunction


  function automatic [51:0] MUX_v_52_2_2;
    input [51:0] input_0;
    input [51:0] input_1;
    input  sel;
    reg [51:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_52_2_2 = result;
  end
  endfunction


  function automatic [52:0] MUX_v_53_2_2;
    input [52:0] input_0;
    input [52:0] input_1;
    input  sel;
    reg [52:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_53_2_2 = result;
  end
  endfunction


  function automatic [55:0] MUX_v_56_2_2;
    input [55:0] input_0;
    input [55:0] input_1;
    input  sel;
    reg [55:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_56_2_2 = result;
  end
  endfunction


  function automatic [56:0] MUX_v_57_2_2;
    input [56:0] input_0;
    input [56:0] input_1;
    input  sel;
    reg [56:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_57_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [10:0] readslicef_12_11_1;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_12_11_1 = tmp[10:0];
  end
  endfunction


  function automatic [0:0] readslicef_12_1_11;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_12_1_11 = tmp[0:0];
  end
  endfunction


  function automatic [11:0] readslicef_13_12_1;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_13_12_1 = tmp[11:0];
  end
  endfunction


  function automatic [0:0] readslicef_13_1_12;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 12;
    readslicef_13_1_12 = tmp[0:0];
  end
  endfunction


  function automatic [12:0] readslicef_14_13_1;
    input [13:0] vector;
    reg [13:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_14_13_1 = tmp[12:0];
  end
  endfunction


  function automatic [16:0] readslicef_18_17_1;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_18_17_1 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_19_18_1;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_19_18_1 = tmp[17:0];
  end
  endfunction


  function automatic [15:0] readslicef_32_16_16;
    input [31:0] vector;
    reg [31:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_32_16_16 = tmp[15:0];
  end
  endfunction


  function automatic [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_53_1_52;
    input [52:0] vector;
    reg [52:0] tmp;
  begin
    tmp = vector >> 52;
    readslicef_53_1_52 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_54_1_53;
    input [53:0] vector;
    reg [53:0] tmp;
  begin
    tmp = vector >> 53;
    readslicef_54_1_53 = tmp[0:0];
  end
  endfunction


  function automatic [56:0] readslicef_58_57_1;
    input [57:0] vector;
    reg [57:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_58_57_1 = tmp[56:0];
  end
  endfunction


  function automatic [13:0] signext_14_13;
    input [12:0] vector;
  begin
    signext_14_13= {{1{vector[12]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2s_7_11 ;
    input [6:0]  vector ;
  begin
    conv_s2s_7_11 = {{4{vector[6]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_7_12 ;
    input [6:0]  vector ;
  begin
    conv_s2s_7_12 = {{5{vector[6]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_7_13 ;
    input [6:0]  vector ;
  begin
    conv_s2s_7_13 = {{6{vector[6]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_11_13 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_13 = {{2{vector[10]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_12_13 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_13 = {vector[11], vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [12:0] conv_s2u_7_13 ;
    input [6:0]  vector ;
  begin
    conv_s2u_7_13 = {{6{vector[6]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2u_8_12 ;
    input [7:0]  vector ;
  begin
    conv_s2u_8_12 = {{4{vector[7]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2u_8_13 ;
    input [7:0]  vector ;
  begin
    conv_s2u_8_13 = {{5{vector[7]}}, vector};
  end
  endfunction


  function automatic [13:0] conv_s2u_8_14 ;
    input [7:0]  vector ;
  begin
    conv_s2u_8_14 = {{6{vector[7]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [13:0] conv_s2u_12_14 ;
    input [11:0]  vector ;
  begin
    conv_s2u_12_14 = {{2{vector[11]}}, vector};
  end
  endfunction


  function automatic [13:0] conv_s2u_13_14 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_14 = {vector[12], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_19 = {vector[17], vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_23_24 ;
    input [22:0]  vector ;
  begin
    conv_s2u_23_24 = {vector[22], vector};
  end
  endfunction


  function automatic [12:0] conv_u2s_1_13 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_13 = {{12{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function automatic [15:0] conv_u2s_4_16 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_16 = {{12{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_10_12 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_12 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2s_11_13 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_13 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2s_12_13 ;
    input [11:0]  vector ;
  begin
    conv_u2s_12_13 =  {1'b0, vector};
  end
  endfunction


  function automatic [14:0] conv_u2s_14_15 ;
    input [13:0]  vector ;
  begin
    conv_u2s_14_15 =  {1'b0, vector};
  end
  endfunction


  function automatic [15:0] conv_u2s_14_16 ;
    input [13:0]  vector ;
  begin
    conv_u2s_14_16 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2s_16_17 =  {1'b0, vector};
  end
  endfunction


  function automatic [17:0] conv_u2s_16_18 ;
    input [15:0]  vector ;
  begin
    conv_u2s_16_18 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_1_12 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_12 = {{11{1'b0}}, vector};
  end
  endfunction


  function automatic [51:0] conv_u2u_1_52 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_52 = {{51{1'b0}}, vector};
  end
  endfunction


  function automatic [53:0] conv_u2u_1_54 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_54 = {{53{1'b0}}, vector};
  end
  endfunction


  function automatic [56:0] conv_u2u_1_57 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_57 = {{56{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_4_11 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_11 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_11_13 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_13 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_u2u_12_13 = {1'b0, vector};
  end
  endfunction


  function automatic [13:0] conv_u2u_12_14 ;
    input [11:0]  vector ;
  begin
    conv_u2u_12_14 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [14:0] conv_u2u_14_15 ;
    input [13:0]  vector ;
  begin
    conv_u2u_14_15 = {1'b0, vector};
  end
  endfunction


  function automatic [15:0] conv_u2u_14_16 ;
    input [13:0]  vector ;
  begin
    conv_u2u_14_16 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_14_17 ;
    input [13:0]  vector ;
  begin
    conv_u2u_14_17 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [17:0] conv_u2u_14_18 ;
    input [13:0]  vector ;
  begin
    conv_u2u_14_18 = {{4{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_17 = {1'b0, vector};
  end
  endfunction


  function automatic [17:0] conv_u2u_17_18 ;
    input [16:0]  vector ;
  begin
    conv_u2u_17_18 = {1'b0, vector};
  end
  endfunction


  function automatic [18:0] conv_u2u_17_19 ;
    input [16:0]  vector ;
  begin
    conv_u2u_17_19 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_30_32 ;
    input [29:0]  vector ;
  begin
    conv_u2u_30_32 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [52:0] conv_u2u_52_53 ;
    input [51:0]  vector ;
  begin
    conv_u2u_52_53 = {1'b0, vector};
  end
  endfunction


  function automatic [53:0] conv_u2u_53_54 ;
    input [52:0]  vector ;
  begin
    conv_u2u_53_54 = {1'b0, vector};
  end
  endfunction


  function automatic [56:0] conv_u2u_56_57 ;
    input [55:0]  vector ;
  begin
    conv_u2u_56_57 = {1'b0, vector};
  end
  endfunction


  function automatic [57:0] conv_u2u_57_58 ;
    input [56:0]  vector ;
  begin
    conv_u2u_57_58 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_struct
// ------------------------------------------------------------------


module stage_struct (
  clk, rst, arst_n, ap_start_rsc_dat, ap_start_rsc_vld, ap_start_rsc_rdy, ap_done_rsc_dat,
      ap_done_rsc_vld, ap_done_rsc_rdy, mode1_rsc_dat, mode1_triosy_lz, in_f_d_rsc_adr,
      in_f_d_rsc_d, in_f_d_rsc_we, in_f_d_rsc_q, in_f_d_rsc_en, in_f_d_triosy_lz,
      in_u_rsc_adr, in_u_rsc_d, in_u_rsc_we, in_u_rsc_q, in_u_rsc_en, in_u_triosy_lz,
      out_f_d_rsc_adr, out_f_d_rsc_d, out_f_d_rsc_we, out_f_d_rsc_q, out_f_d_rsc_en,
      out_f_d_triosy_lz, out_u_rsc_adr, out_u_rsc_d, out_u_rsc_we, out_u_rsc_q, out_u_rsc_en,
      out_u_triosy_lz, out1_rsc_dat_u, out1_rsc_dat_d, out1_rsc_vld, out1_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input [15:0] mode1_rsc_dat;
  output mode1_triosy_lz;
  output [9:0] in_f_d_rsc_adr;
  output [63:0] in_f_d_rsc_d;
  output in_f_d_rsc_we;
  input [63:0] in_f_d_rsc_q;
  output in_f_d_rsc_en;
  output in_f_d_triosy_lz;
  output [9:0] in_u_rsc_adr;
  output [15:0] in_u_rsc_d;
  output in_u_rsc_we;
  input [15:0] in_u_rsc_q;
  output in_u_rsc_en;
  output in_u_triosy_lz;
  output [9:0] out_f_d_rsc_adr;
  output [63:0] out_f_d_rsc_d;
  output out_f_d_rsc_we;
  input [63:0] out_f_d_rsc_q;
  output out_f_d_rsc_en;
  output out_f_d_triosy_lz;
  output [9:0] out_u_rsc_adr;
  output [15:0] out_u_rsc_d;
  output out_u_rsc_we;
  input [15:0] out_u_rsc_q;
  output out_u_rsc_en;
  output out_u_triosy_lz;
  output [15:0] out1_rsc_dat_u;
  output [63:0] out1_rsc_dat_d;
  output out1_rsc_vld;
  input out1_rsc_rdy;


  // Interconnect Declarations
  wire [9:0] in_f_d_rsci_adr_d;
  wire [63:0] in_f_d_rsci_d_d;
  wire in_f_d_rsci_en_d;
  wire [63:0] in_f_d_rsci_q_d;
  wire in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [9:0] in_u_rsci_adr_d;
  wire [15:0] in_u_rsci_d_d;
  wire in_u_rsci_en_d;
  wire [15:0] in_u_rsci_q_d;
  wire in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [9:0] out_f_d_rsci_adr_d;
  wire [63:0] out_f_d_rsci_d_d;
  wire out_f_d_rsci_en_d;
  wire [63:0] out_f_d_rsci_q_d;
  wire out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [9:0] out_u_rsci_adr_d;
  wire [15:0] out_u_rsci_d_d;
  wire out_u_rsci_en_d;
  wire [15:0] out_u_rsci_q_d;
  wire out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [9:0] BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr;
  wire [13:0] BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out;
  wire BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en;
  wire [13:0] BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out;
  wire BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en;
  wire [13:0] BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out;
  wire BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en;
  wire [13:0] BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out;
  wire BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en;
  wire [61:0] r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out;
  wire r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en;
  wire [63:0] BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out;
  wire [15:0] BUTTERFLY_i_div_cmp_a;
  wire [15:0] BUTTERFLY_i_div_cmp_b;
  wire [79:0] out1_rsc_dat;
  wire in_f_d_rsci_we_d_iff;
  wire in_u_rsci_we_d_iff;
  wire out_f_d_rsci_we_d_iff;
  wire out_u_rsci_we_d_iff;
  reg BUTTERFLY_i_div_cmp_z_15;
  reg BUTTERFLY_i_div_cmp_z_14;
  reg BUTTERFLY_i_div_cmp_z_13;
  reg BUTTERFLY_i_div_cmp_z_12;
  reg BUTTERFLY_i_div_cmp_z_11;
  reg BUTTERFLY_i_div_cmp_z_10;
  reg BUTTERFLY_i_div_cmp_z_9;
  reg BUTTERFLY_i_div_cmp_z_8;
  reg BUTTERFLY_i_div_cmp_z_7;
  reg BUTTERFLY_i_div_cmp_z_6;
  reg BUTTERFLY_i_div_cmp_z_5;
  reg BUTTERFLY_i_div_cmp_z_4;
  reg BUTTERFLY_i_div_cmp_z_3;
  reg BUTTERFLY_i_div_cmp_z_2;
  reg BUTTERFLY_i_div_cmp_z_1;
  reg BUTTERFLY_i_div_cmp_z_0;


  // Interconnect Declarations for Component Instantiations 
  wire [15:0] nl_stage_run_inst_BUTTERFLY_i_div_cmp_z;
  assign nl_stage_run_inst_BUTTERFLY_i_div_cmp_z = {BUTTERFLY_i_div_cmp_z_15 , BUTTERFLY_i_div_cmp_z_14
      , BUTTERFLY_i_div_cmp_z_13 , BUTTERFLY_i_div_cmp_z_12 , BUTTERFLY_i_div_cmp_z_11
      , BUTTERFLY_i_div_cmp_z_10 , BUTTERFLY_i_div_cmp_z_9 , BUTTERFLY_i_div_cmp_z_8
      , BUTTERFLY_i_div_cmp_z_7 , BUTTERFLY_i_div_cmp_z_6 , BUTTERFLY_i_div_cmp_z_5
      , BUTTERFLY_i_div_cmp_z_4 , BUTTERFLY_i_div_cmp_z_3 , BUTTERFLY_i_div_cmp_z_2
      , BUTTERFLY_i_div_cmp_z_1 , BUTTERFLY_i_div_cmp_z_0};
  
  `ifdef USE_PDK_ROM

    rom1_14m16h3v2 rom1_14(
      .CLK(clk),
      .CEN(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en),
      .A(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .Q(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out)
    );

    rom2_14m16h3v2 rom2_14(
      .CLK(clk),
      .CEN(BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en),
      .A(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .Q(BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out)
    );

    rom3_14m16h3v2 rom3_14(
      .CLK(clk),
      .CEN(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en),
      .A(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .Q(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out)
    );


    rom4_14m16h3v2 rom4_14(
      .CLK(clk),
      .CEN(BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en),
      .A(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .Q(BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out)
    );


    rom5_62m16h3v2 rom5_62(
      .CLK(clk),
      .CEN(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en),
      .A(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_addr),
      .Q(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out)
    );

    rom6_64m16h3v2 rom6_64(
      .CLK(clk),
      .CEN(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en),
      .A(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_addr),
      .Q(BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out)
    );
  
  
  `else
  stagemgc_rom_sync_regout_14_1024_14_1_0_0_1_0_1_0_0_0_1_60  BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp
      (
      .addr(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .data_out(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out),
      .clk(clk),
      .s_rst(rst),
      .a_rst(arst_n),
      .en(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en)
    );
  stagemgc_rom_sync_regout_13_1024_14_1_0_0_1_0_1_0_0_0_1_60  BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp
      (
      .addr(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .data_out(BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out),
      .clk(clk),
      .s_rst(rst),
      .a_rst(arst_n),
      .en(BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en)
    );
  stagemgc_rom_sync_regout_12_1024_14_1_0_0_1_0_1_0_0_0_1_60  BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp
      (
      .addr(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .data_out(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out),
      .clk(clk),
      .s_rst(rst),
      .a_rst(arst_n),
      .en(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en)
    );
  stagemgc_rom_sync_regout_11_1024_14_1_0_0_1_0_1_0_0_0_1_60  BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp
      (
      .addr(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .data_out(BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out),
      .clk(clk),
      .s_rst(rst),
      .a_rst(arst_n),
      .en(BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en)
    );
  stagemgc_rom_sync_regout_10_1024_62_1_0_0_1_0_1_0_0_0_1_60  r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp
      (
      .addr(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .data_out(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out),
      .clk(clk),
      .s_rst(rst),
      .a_rst(arst_n),
      .en(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en)
    );
  stagemgc_rom_sync_regout_9_1024_64_1_0_0_1_0_1_0_0_0_1_60  BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp
      (
      .addr(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .data_out(BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out),
      .clk(clk),
      .s_rst(rst),
      .a_rst(arst_n),
      .en(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en)
    );
  `endif
  stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_4_64_10_1024_1024_64_5_gen
      in_f_d_rsci (
      .en(in_f_d_rsc_en),
      .q(in_f_d_rsc_q),
      .we(in_f_d_rsc_we),
      .d(in_f_d_rsc_d),
      .adr(in_f_d_rsc_adr),
      .adr_d(in_f_d_rsci_adr_d),
      .d_d(in_f_d_rsci_d_d),
      .en_d(in_f_d_rsci_en_d),
      .we_d(in_f_d_rsci_we_d_iff),
      .q_d(in_f_d_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(in_f_d_rsci_we_d_iff)
    );
  stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_5_16_10_1024_1024_16_5_gen
      in_u_rsci (
      .en(in_u_rsc_en),
      .q(in_u_rsc_q),
      .we(in_u_rsc_we),
      .d(in_u_rsc_d),
      .adr(in_u_rsc_adr),
      .adr_d(in_u_rsci_adr_d),
      .d_d(in_u_rsci_d_d),
      .en_d(in_u_rsci_en_d),
      .we_d(in_u_rsci_we_d_iff),
      .q_d(in_u_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(in_u_rsci_we_d_iff)
    );
  stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_6_64_10_1024_1024_64_5_gen
      out_f_d_rsci (
      .en(out_f_d_rsc_en),
      .q(out_f_d_rsc_q),
      .we(out_f_d_rsc_we),
      .d(out_f_d_rsc_d),
      .adr(out_f_d_rsc_adr),
      .adr_d(out_f_d_rsci_adr_d),
      .d_d(out_f_d_rsci_d_d),
      .en_d(out_f_d_rsci_en_d),
      .we_d(out_f_d_rsci_we_d_iff),
      .q_d(out_f_d_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(out_f_d_rsci_we_d_iff)
    );
  stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_7_16_10_1024_1024_16_5_gen
      out_u_rsci (
      .en(out_u_rsc_en),
      .q(out_u_rsc_q),
      .we(out_u_rsc_we),
      .d(out_u_rsc_d),
      .adr(out_u_rsc_adr),
      .adr_d(out_u_rsci_adr_d),
      .d_d(out_u_rsci_d_d),
      .en_d(out_u_rsci_en_d),
      .we_d(out_u_rsci_we_d_iff),
      .q_d(out_u_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(out_u_rsci_we_d_iff)
    );
  stage_run stage_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .ap_start_rsc_dat(ap_start_rsc_dat),
      .ap_start_rsc_vld(ap_start_rsc_vld),
      .ap_start_rsc_rdy(ap_start_rsc_rdy),
      .ap_done_rsc_dat(ap_done_rsc_dat),
      .ap_done_rsc_vld(ap_done_rsc_vld),
      .ap_done_rsc_rdy(ap_done_rsc_rdy),
      .mode1_rsc_dat(mode1_rsc_dat),
      .mode1_triosy_lz(mode1_triosy_lz),
      .in_f_d_triosy_lz(in_f_d_triosy_lz),
      .in_u_triosy_lz(in_u_triosy_lz),
      .out_f_d_triosy_lz(out_f_d_triosy_lz),
      .out_u_triosy_lz(out_u_triosy_lz),
      .out1_rsc_dat(out1_rsc_dat),
      .out1_rsc_vld(out1_rsc_vld),
      .out1_rsc_rdy(out1_rsc_rdy),
      .in_f_d_rsci_adr_d(in_f_d_rsci_adr_d),
      .in_f_d_rsci_d_d(in_f_d_rsci_d_d),
      .in_f_d_rsci_en_d(in_f_d_rsci_en_d),
      .in_f_d_rsci_q_d(in_f_d_rsci_q_d),
      .in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .in_u_rsci_adr_d(in_u_rsci_adr_d),
      .in_u_rsci_d_d(in_u_rsci_d_d),
      .in_u_rsci_en_d(in_u_rsci_en_d),
      .in_u_rsci_q_d(in_u_rsci_q_d),
      .in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .out_f_d_rsci_adr_d(out_f_d_rsci_adr_d),
      .out_f_d_rsci_d_d(out_f_d_rsci_d_d),
      .out_f_d_rsci_en_d(out_f_d_rsci_en_d),
      .out_f_d_rsci_q_d(out_f_d_rsci_q_d),
      .out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .out_u_rsci_adr_d(out_u_rsci_adr_d),
      .out_u_rsci_d_d(out_u_rsci_d_d),
      .out_u_rsci_en_d(out_u_rsci_en_d),
      .out_u_rsci_q_d(out_u_rsci_q_d),
      .out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out),
      .BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en),
      .BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out(BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out),
      .BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en(BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en),
      .BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out),
      .BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en),
      .BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out(BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out),
      .BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en(BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en),
      .r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out),
      .r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en),
      .BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out(BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out),
      .BUTTERFLY_i_div_cmp_a(BUTTERFLY_i_div_cmp_a),
      .BUTTERFLY_i_div_cmp_b(BUTTERFLY_i_div_cmp_b),
      .BUTTERFLY_i_div_cmp_z(nl_stage_run_inst_BUTTERFLY_i_div_cmp_z[15:0]),
      .in_f_d_rsci_we_d_pff(in_f_d_rsci_we_d_iff),
      .in_u_rsci_we_d_pff(in_u_rsci_we_d_iff),
      .out_f_d_rsci_we_d_pff(out_f_d_rsci_we_d_iff),
      .out_u_rsci_we_d_pff(out_u_rsci_we_d_iff)
    );
  assign out1_rsc_dat_d = out1_rsc_dat[63:0];
  assign out1_rsc_dat_u = out1_rsc_dat[79:64];
  always @(BUTTERFLY_i_div_cmp_a or BUTTERFLY_i_div_cmp_b)
  begin : mgc_div_16_16_0_1_b0_line_26
    // Interconnect Declarations
    reg [16:0] divmod6449_2_diff_1;
    reg [16:0] divmod6449_2_diff_2;
    reg [16:0] divmod6449_2_diff_3;
    reg [16:0] divmod6449_2_diff_4;
    reg [16:0] divmod6449_2_diff_5;
    reg [16:0] divmod6449_2_diff_6;
    reg [16:0] divmod6449_2_diff_7;
    reg [16:0] divmod6449_2_diff_8;
    reg [16:0] divmod6449_2_diff_9;
    reg [16:0] divmod6449_2_diff_10;
    reg [16:0] divmod6449_2_diff_11;
    reg [16:0] divmod6449_2_diff_12;
    reg [16:0] divmod6449_2_diff_13;
    reg [16:0] divmod6449_2_diff_14;
    reg [16:0] divmod6449_2_diff_15;
    reg divmod6449_2_lbuf_29_15;
    reg divmod6449_2_lbuf_28_14;
    reg divmod6449_2_lbuf_28_15;
    reg divmod6449_2_lbuf_27_13;
    reg divmod6449_2_lbuf_27_14;
    reg divmod6449_2_lbuf_27_15;
    reg divmod6449_2_lbuf_26_12;
    reg divmod6449_2_lbuf_26_13;
    reg divmod6449_2_lbuf_26_14;
    reg divmod6449_2_lbuf_26_15;
    reg divmod6449_2_lbuf_25_11;
    reg divmod6449_2_lbuf_25_12;
    reg divmod6449_2_lbuf_25_13;
    reg divmod6449_2_lbuf_25_14;
    reg divmod6449_2_lbuf_25_15;
    reg divmod6449_2_lbuf_24_10;
    reg divmod6449_2_lbuf_24_11;
    reg divmod6449_2_lbuf_24_12;
    reg divmod6449_2_lbuf_24_13;
    reg divmod6449_2_lbuf_24_14;
    reg divmod6449_2_lbuf_24_15;
    reg divmod6449_2_lbuf_23_9;
    reg divmod6449_2_lbuf_23_10;
    reg divmod6449_2_lbuf_23_11;
    reg divmod6449_2_lbuf_23_12;
    reg divmod6449_2_lbuf_23_13;
    reg divmod6449_2_lbuf_23_14;
    reg divmod6449_2_lbuf_23_15;
    reg divmod6449_2_lbuf_22_8;
    reg divmod6449_2_lbuf_22_9;
    reg divmod6449_2_lbuf_22_10;
    reg divmod6449_2_lbuf_22_11;
    reg divmod6449_2_lbuf_22_12;
    reg divmod6449_2_lbuf_22_13;
    reg divmod6449_2_lbuf_22_14;
    reg divmod6449_2_lbuf_22_15;
    reg divmod6449_2_lbuf_21_7;
    reg divmod6449_2_lbuf_21_8;
    reg divmod6449_2_lbuf_21_9;
    reg divmod6449_2_lbuf_21_10;
    reg divmod6449_2_lbuf_21_11;
    reg divmod6449_2_lbuf_21_12;
    reg divmod6449_2_lbuf_21_13;
    reg divmod6449_2_lbuf_21_14;
    reg divmod6449_2_lbuf_21_15;
    reg divmod6449_2_lbuf_20_6;
    reg divmod6449_2_lbuf_20_7;
    reg divmod6449_2_lbuf_20_8;
    reg divmod6449_2_lbuf_20_9;
    reg divmod6449_2_lbuf_20_10;
    reg divmod6449_2_lbuf_20_11;
    reg divmod6449_2_lbuf_20_12;
    reg divmod6449_2_lbuf_20_13;
    reg divmod6449_2_lbuf_20_14;
    reg divmod6449_2_lbuf_20_15;
    reg divmod6449_2_lbuf_19_5;
    reg divmod6449_2_lbuf_19_6;
    reg divmod6449_2_lbuf_19_7;
    reg divmod6449_2_lbuf_19_8;
    reg divmod6449_2_lbuf_19_9;
    reg divmod6449_2_lbuf_19_10;
    reg divmod6449_2_lbuf_19_11;
    reg divmod6449_2_lbuf_19_12;
    reg divmod6449_2_lbuf_19_13;
    reg divmod6449_2_lbuf_19_14;
    reg divmod6449_2_lbuf_19_15;
    reg divmod6449_2_lbuf_18_4;
    reg divmod6449_2_lbuf_18_5;
    reg divmod6449_2_lbuf_18_6;
    reg divmod6449_2_lbuf_18_7;
    reg divmod6449_2_lbuf_18_8;
    reg divmod6449_2_lbuf_18_9;
    reg divmod6449_2_lbuf_18_10;
    reg divmod6449_2_lbuf_18_11;
    reg divmod6449_2_lbuf_18_12;
    reg divmod6449_2_lbuf_18_13;
    reg divmod6449_2_lbuf_18_14;
    reg divmod6449_2_lbuf_18_15;
    reg divmod6449_2_lbuf_17_3;
    reg divmod6449_2_lbuf_17_4;
    reg divmod6449_2_lbuf_17_5;
    reg divmod6449_2_lbuf_17_6;
    reg divmod6449_2_lbuf_17_7;
    reg divmod6449_2_lbuf_17_8;
    reg divmod6449_2_lbuf_17_9;
    reg divmod6449_2_lbuf_17_10;
    reg divmod6449_2_lbuf_17_11;
    reg divmod6449_2_lbuf_17_12;
    reg divmod6449_2_lbuf_17_13;
    reg divmod6449_2_lbuf_17_14;
    reg divmod6449_2_lbuf_17_15;
    reg divmod6449_2_lbuf_16_2;
    reg divmod6449_2_lbuf_16_3;
    reg divmod6449_2_lbuf_16_4;
    reg divmod6449_2_lbuf_16_5;
    reg divmod6449_2_lbuf_16_6;
    reg divmod6449_2_lbuf_16_7;
    reg divmod6449_2_lbuf_16_8;
    reg divmod6449_2_lbuf_16_9;
    reg divmod6449_2_lbuf_16_10;
    reg divmod6449_2_lbuf_16_11;
    reg divmod6449_2_lbuf_16_12;
    reg divmod6449_2_lbuf_16_13;
    reg divmod6449_2_lbuf_16_14;
    reg divmod6449_2_lbuf_16_15;
    reg [15:0] divmod6449_2_lbuf_15_0_1;
    reg divmod6449_2_lbuf_15;
    reg divmod6449_2_lbuf_15_1;
    reg divmod6449_2_lbuf_15_2;
    reg divmod6449_2_lbuf_15_3;
    reg divmod6449_2_lbuf_15_4;
    reg divmod6449_2_lbuf_15_5;
    reg divmod6449_2_lbuf_15_6;
    reg divmod6449_2_lbuf_15_7;
    reg divmod6449_2_lbuf_15_8;
    reg divmod6449_2_lbuf_15_9;
    reg divmod6449_2_lbuf_15_10;
    reg divmod6449_2_lbuf_15_11;
    reg divmod6449_2_lbuf_15_12;
    reg divmod6449_2_lbuf_15_13;

    reg[16:0] divmod6449_2_loop951_16_acc_1_nl;
    reg[18:0] nl_divmod6449_2_loop951_16_acc_1_nl;
    divmod6449_2_lbuf_15_0_1 = BUTTERFLY_i_div_cmp_a;
    divmod6449_2_diff_1 = conv_u2u_1_17(divmod6449_2_lbuf_15_0_1[15]) + ({1'b1 ,
        (~ BUTTERFLY_i_div_cmp_b)}) + 17'b00000000000000001;
    if ( divmod6449_2_diff_1[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_15_0_1[15] = divmod6449_2_diff_1[0];
    end
    divmod6449_2_lbuf_16_2 = divmod6449_2_lbuf_15_0_1[15];
    divmod6449_2_lbuf_15 = divmod6449_2_lbuf_15_0_1[14];
    divmod6449_2_diff_2 = conv_u2u_2_17(divmod6449_2_lbuf_15_0_1[15:14]) + ({1'b1
        , (~ BUTTERFLY_i_div_cmp_b)}) + 17'b00000000000000001;
    if ( divmod6449_2_diff_2[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_16_2 = divmod6449_2_diff_2[1];
      divmod6449_2_lbuf_15 = divmod6449_2_diff_2[0];
    end
    divmod6449_2_lbuf_17_3 = divmod6449_2_lbuf_16_2;
    divmod6449_2_lbuf_16_3 = divmod6449_2_lbuf_15;
    divmod6449_2_lbuf_15_1 = divmod6449_2_lbuf_15_0_1[13];
    divmod6449_2_diff_3 = conv_u2u_3_17({divmod6449_2_lbuf_16_2 , divmod6449_2_lbuf_15
        , (divmod6449_2_lbuf_15_0_1[13])}) + ({1'b1 , (~ BUTTERFLY_i_div_cmp_b)})
        + 17'b00000000000000001;
    if ( divmod6449_2_diff_3[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_17_3 = divmod6449_2_diff_3[2];
      divmod6449_2_lbuf_16_3 = divmod6449_2_diff_3[1];
      divmod6449_2_lbuf_15_1 = divmod6449_2_diff_3[0];
    end
    divmod6449_2_lbuf_18_4 = divmod6449_2_lbuf_17_3;
    divmod6449_2_lbuf_17_4 = divmod6449_2_lbuf_16_3;
    divmod6449_2_lbuf_16_4 = divmod6449_2_lbuf_15_1;
    divmod6449_2_lbuf_15_2 = divmod6449_2_lbuf_15_0_1[12];
    divmod6449_2_diff_4 = conv_u2u_4_17({divmod6449_2_lbuf_17_3 , divmod6449_2_lbuf_16_3
        , divmod6449_2_lbuf_15_1 , (divmod6449_2_lbuf_15_0_1[12])}) + ({1'b1 , (~
        BUTTERFLY_i_div_cmp_b)}) + 17'b00000000000000001;
    if ( divmod6449_2_diff_4[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_18_4 = divmod6449_2_diff_4[3];
      divmod6449_2_lbuf_17_4 = divmod6449_2_diff_4[2];
      divmod6449_2_lbuf_16_4 = divmod6449_2_diff_4[1];
      divmod6449_2_lbuf_15_2 = divmod6449_2_diff_4[0];
    end
    divmod6449_2_lbuf_19_5 = divmod6449_2_lbuf_18_4;
    divmod6449_2_lbuf_18_5 = divmod6449_2_lbuf_17_4;
    divmod6449_2_lbuf_17_5 = divmod6449_2_lbuf_16_4;
    divmod6449_2_lbuf_16_5 = divmod6449_2_lbuf_15_2;
    divmod6449_2_lbuf_15_3 = divmod6449_2_lbuf_15_0_1[11];
    divmod6449_2_diff_5 = conv_u2u_5_17({divmod6449_2_lbuf_18_4 , divmod6449_2_lbuf_17_4
        , divmod6449_2_lbuf_16_4 , divmod6449_2_lbuf_15_2 , (divmod6449_2_lbuf_15_0_1[11])})
        + ({1'b1 , (~ BUTTERFLY_i_div_cmp_b)}) + 17'b00000000000000001;
    if ( divmod6449_2_diff_5[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_19_5 = divmod6449_2_diff_5[4];
      divmod6449_2_lbuf_18_5 = divmod6449_2_diff_5[3];
      divmod6449_2_lbuf_17_5 = divmod6449_2_diff_5[2];
      divmod6449_2_lbuf_16_5 = divmod6449_2_diff_5[1];
      divmod6449_2_lbuf_15_3 = divmod6449_2_diff_5[0];
    end
    divmod6449_2_lbuf_20_6 = divmod6449_2_lbuf_19_5;
    divmod6449_2_lbuf_19_6 = divmod6449_2_lbuf_18_5;
    divmod6449_2_lbuf_18_6 = divmod6449_2_lbuf_17_5;
    divmod6449_2_lbuf_17_6 = divmod6449_2_lbuf_16_5;
    divmod6449_2_lbuf_16_6 = divmod6449_2_lbuf_15_3;
    divmod6449_2_lbuf_15_4 = divmod6449_2_lbuf_15_0_1[10];
    divmod6449_2_diff_6 = conv_u2u_6_17({divmod6449_2_lbuf_19_5 , divmod6449_2_lbuf_18_5
        , divmod6449_2_lbuf_17_5 , divmod6449_2_lbuf_16_5 , divmod6449_2_lbuf_15_3
        , (divmod6449_2_lbuf_15_0_1[10])}) + ({1'b1 , (~ BUTTERFLY_i_div_cmp_b)})
        + 17'b00000000000000001;
    if ( divmod6449_2_diff_6[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_20_6 = divmod6449_2_diff_6[5];
      divmod6449_2_lbuf_19_6 = divmod6449_2_diff_6[4];
      divmod6449_2_lbuf_18_6 = divmod6449_2_diff_6[3];
      divmod6449_2_lbuf_17_6 = divmod6449_2_diff_6[2];
      divmod6449_2_lbuf_16_6 = divmod6449_2_diff_6[1];
      divmod6449_2_lbuf_15_4 = divmod6449_2_diff_6[0];
    end
    divmod6449_2_lbuf_21_7 = divmod6449_2_lbuf_20_6;
    divmod6449_2_lbuf_20_7 = divmod6449_2_lbuf_19_6;
    divmod6449_2_lbuf_19_7 = divmod6449_2_lbuf_18_6;
    divmod6449_2_lbuf_18_7 = divmod6449_2_lbuf_17_6;
    divmod6449_2_lbuf_17_7 = divmod6449_2_lbuf_16_6;
    divmod6449_2_lbuf_16_7 = divmod6449_2_lbuf_15_4;
    divmod6449_2_lbuf_15_5 = divmod6449_2_lbuf_15_0_1[9];
    divmod6449_2_diff_7 = conv_u2u_7_17({divmod6449_2_lbuf_20_6 , divmod6449_2_lbuf_19_6
        , divmod6449_2_lbuf_18_6 , divmod6449_2_lbuf_17_6 , divmod6449_2_lbuf_16_6
        , divmod6449_2_lbuf_15_4 , (divmod6449_2_lbuf_15_0_1[9])}) + ({1'b1 , (~
        BUTTERFLY_i_div_cmp_b)}) + 17'b00000000000000001;
    if ( divmod6449_2_diff_7[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_21_7 = divmod6449_2_diff_7[6];
      divmod6449_2_lbuf_20_7 = divmod6449_2_diff_7[5];
      divmod6449_2_lbuf_19_7 = divmod6449_2_diff_7[4];
      divmod6449_2_lbuf_18_7 = divmod6449_2_diff_7[3];
      divmod6449_2_lbuf_17_7 = divmod6449_2_diff_7[2];
      divmod6449_2_lbuf_16_7 = divmod6449_2_diff_7[1];
      divmod6449_2_lbuf_15_5 = divmod6449_2_diff_7[0];
    end
    divmod6449_2_lbuf_22_8 = divmod6449_2_lbuf_21_7;
    divmod6449_2_lbuf_21_8 = divmod6449_2_lbuf_20_7;
    divmod6449_2_lbuf_20_8 = divmod6449_2_lbuf_19_7;
    divmod6449_2_lbuf_19_8 = divmod6449_2_lbuf_18_7;
    divmod6449_2_lbuf_18_8 = divmod6449_2_lbuf_17_7;
    divmod6449_2_lbuf_17_8 = divmod6449_2_lbuf_16_7;
    divmod6449_2_lbuf_16_8 = divmod6449_2_lbuf_15_5;
    divmod6449_2_lbuf_15_6 = divmod6449_2_lbuf_15_0_1[8];
    divmod6449_2_diff_8 = conv_u2u_8_17({divmod6449_2_lbuf_21_7 , divmod6449_2_lbuf_20_7
        , divmod6449_2_lbuf_19_7 , divmod6449_2_lbuf_18_7 , divmod6449_2_lbuf_17_7
        , divmod6449_2_lbuf_16_7 , divmod6449_2_lbuf_15_5 , (divmod6449_2_lbuf_15_0_1[8])})
        + ({1'b1 , (~ BUTTERFLY_i_div_cmp_b)}) + 17'b00000000000000001;
    if ( divmod6449_2_diff_8[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_22_8 = divmod6449_2_diff_8[7];
      divmod6449_2_lbuf_21_8 = divmod6449_2_diff_8[6];
      divmod6449_2_lbuf_20_8 = divmod6449_2_diff_8[5];
      divmod6449_2_lbuf_19_8 = divmod6449_2_diff_8[4];
      divmod6449_2_lbuf_18_8 = divmod6449_2_diff_8[3];
      divmod6449_2_lbuf_17_8 = divmod6449_2_diff_8[2];
      divmod6449_2_lbuf_16_8 = divmod6449_2_diff_8[1];
      divmod6449_2_lbuf_15_6 = divmod6449_2_diff_8[0];
    end
    divmod6449_2_lbuf_23_9 = divmod6449_2_lbuf_22_8;
    divmod6449_2_lbuf_22_9 = divmod6449_2_lbuf_21_8;
    divmod6449_2_lbuf_21_9 = divmod6449_2_lbuf_20_8;
    divmod6449_2_lbuf_20_9 = divmod6449_2_lbuf_19_8;
    divmod6449_2_lbuf_19_9 = divmod6449_2_lbuf_18_8;
    divmod6449_2_lbuf_18_9 = divmod6449_2_lbuf_17_8;
    divmod6449_2_lbuf_17_9 = divmod6449_2_lbuf_16_8;
    divmod6449_2_lbuf_16_9 = divmod6449_2_lbuf_15_6;
    divmod6449_2_lbuf_15_7 = divmod6449_2_lbuf_15_0_1[7];
    divmod6449_2_diff_9 = conv_u2u_9_17({divmod6449_2_lbuf_22_8 , divmod6449_2_lbuf_21_8
        , divmod6449_2_lbuf_20_8 , divmod6449_2_lbuf_19_8 , divmod6449_2_lbuf_18_8
        , divmod6449_2_lbuf_17_8 , divmod6449_2_lbuf_16_8 , divmod6449_2_lbuf_15_6
        , (divmod6449_2_lbuf_15_0_1[7])}) + ({1'b1 , (~ BUTTERFLY_i_div_cmp_b)})
        + 17'b00000000000000001;
    if ( divmod6449_2_diff_9[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_23_9 = divmod6449_2_diff_9[8];
      divmod6449_2_lbuf_22_9 = divmod6449_2_diff_9[7];
      divmod6449_2_lbuf_21_9 = divmod6449_2_diff_9[6];
      divmod6449_2_lbuf_20_9 = divmod6449_2_diff_9[5];
      divmod6449_2_lbuf_19_9 = divmod6449_2_diff_9[4];
      divmod6449_2_lbuf_18_9 = divmod6449_2_diff_9[3];
      divmod6449_2_lbuf_17_9 = divmod6449_2_diff_9[2];
      divmod6449_2_lbuf_16_9 = divmod6449_2_diff_9[1];
      divmod6449_2_lbuf_15_7 = divmod6449_2_diff_9[0];
    end
    divmod6449_2_lbuf_24_10 = divmod6449_2_lbuf_23_9;
    divmod6449_2_lbuf_23_10 = divmod6449_2_lbuf_22_9;
    divmod6449_2_lbuf_22_10 = divmod6449_2_lbuf_21_9;
    divmod6449_2_lbuf_21_10 = divmod6449_2_lbuf_20_9;
    divmod6449_2_lbuf_20_10 = divmod6449_2_lbuf_19_9;
    divmod6449_2_lbuf_19_10 = divmod6449_2_lbuf_18_9;
    divmod6449_2_lbuf_18_10 = divmod6449_2_lbuf_17_9;
    divmod6449_2_lbuf_17_10 = divmod6449_2_lbuf_16_9;
    divmod6449_2_lbuf_16_10 = divmod6449_2_lbuf_15_7;
    divmod6449_2_lbuf_15_8 = divmod6449_2_lbuf_15_0_1[6];
    divmod6449_2_diff_10 = conv_u2u_10_17({divmod6449_2_lbuf_23_9 , divmod6449_2_lbuf_22_9
        , divmod6449_2_lbuf_21_9 , divmod6449_2_lbuf_20_9 , divmod6449_2_lbuf_19_9
        , divmod6449_2_lbuf_18_9 , divmod6449_2_lbuf_17_9 , divmod6449_2_lbuf_16_9
        , divmod6449_2_lbuf_15_7 , (divmod6449_2_lbuf_15_0_1[6])}) + ({1'b1 , (~
        BUTTERFLY_i_div_cmp_b)}) + 17'b00000000000000001;
    if ( divmod6449_2_diff_10[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_23_10 = divmod6449_2_diff_10[8];
      divmod6449_2_lbuf_22_10 = divmod6449_2_diff_10[7];
      divmod6449_2_lbuf_24_10 = divmod6449_2_diff_10[9];
      divmod6449_2_lbuf_21_10 = divmod6449_2_diff_10[6];
      divmod6449_2_lbuf_20_10 = divmod6449_2_diff_10[5];
      divmod6449_2_lbuf_19_10 = divmod6449_2_diff_10[4];
      divmod6449_2_lbuf_18_10 = divmod6449_2_diff_10[3];
      divmod6449_2_lbuf_17_10 = divmod6449_2_diff_10[2];
      divmod6449_2_lbuf_16_10 = divmod6449_2_diff_10[1];
      divmod6449_2_lbuf_15_8 = divmod6449_2_diff_10[0];
    end
    divmod6449_2_lbuf_25_11 = divmod6449_2_lbuf_24_10;
    divmod6449_2_lbuf_24_11 = divmod6449_2_lbuf_23_10;
    divmod6449_2_lbuf_23_11 = divmod6449_2_lbuf_22_10;
    divmod6449_2_lbuf_22_11 = divmod6449_2_lbuf_21_10;
    divmod6449_2_lbuf_21_11 = divmod6449_2_lbuf_20_10;
    divmod6449_2_lbuf_20_11 = divmod6449_2_lbuf_19_10;
    divmod6449_2_lbuf_19_11 = divmod6449_2_lbuf_18_10;
    divmod6449_2_lbuf_18_11 = divmod6449_2_lbuf_17_10;
    divmod6449_2_lbuf_17_11 = divmod6449_2_lbuf_16_10;
    divmod6449_2_lbuf_16_11 = divmod6449_2_lbuf_15_8;
    divmod6449_2_lbuf_15_9 = divmod6449_2_lbuf_15_0_1[5];
    divmod6449_2_diff_11 = conv_u2u_11_17({divmod6449_2_lbuf_24_10 , divmod6449_2_lbuf_23_10
        , divmod6449_2_lbuf_22_10 , divmod6449_2_lbuf_21_10 , divmod6449_2_lbuf_20_10
        , divmod6449_2_lbuf_19_10 , divmod6449_2_lbuf_18_10 , divmod6449_2_lbuf_17_10
        , divmod6449_2_lbuf_16_10 , divmod6449_2_lbuf_15_8 , (divmod6449_2_lbuf_15_0_1[5])})
        + ({1'b1 , (~ BUTTERFLY_i_div_cmp_b)}) + 17'b00000000000000001;
    if ( divmod6449_2_diff_11[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_23_11 = divmod6449_2_diff_11[8];
      divmod6449_2_lbuf_22_11 = divmod6449_2_diff_11[7];
      divmod6449_2_lbuf_24_11 = divmod6449_2_diff_11[9];
      divmod6449_2_lbuf_21_11 = divmod6449_2_diff_11[6];
      divmod6449_2_lbuf_25_11 = divmod6449_2_diff_11[10];
      divmod6449_2_lbuf_20_11 = divmod6449_2_diff_11[5];
      divmod6449_2_lbuf_19_11 = divmod6449_2_diff_11[4];
      divmod6449_2_lbuf_18_11 = divmod6449_2_diff_11[3];
      divmod6449_2_lbuf_17_11 = divmod6449_2_diff_11[2];
      divmod6449_2_lbuf_16_11 = divmod6449_2_diff_11[1];
      divmod6449_2_lbuf_15_9 = divmod6449_2_diff_11[0];
    end
    divmod6449_2_lbuf_26_12 = divmod6449_2_lbuf_25_11;
    divmod6449_2_lbuf_25_12 = divmod6449_2_lbuf_24_11;
    divmod6449_2_lbuf_24_12 = divmod6449_2_lbuf_23_11;
    divmod6449_2_lbuf_23_12 = divmod6449_2_lbuf_22_11;
    divmod6449_2_lbuf_22_12 = divmod6449_2_lbuf_21_11;
    divmod6449_2_lbuf_21_12 = divmod6449_2_lbuf_20_11;
    divmod6449_2_lbuf_20_12 = divmod6449_2_lbuf_19_11;
    divmod6449_2_lbuf_19_12 = divmod6449_2_lbuf_18_11;
    divmod6449_2_lbuf_18_12 = divmod6449_2_lbuf_17_11;
    divmod6449_2_lbuf_17_12 = divmod6449_2_lbuf_16_11;
    divmod6449_2_lbuf_16_12 = divmod6449_2_lbuf_15_9;
    divmod6449_2_lbuf_15_10 = divmod6449_2_lbuf_15_0_1[4];
    divmod6449_2_diff_12 = conv_u2u_12_17({divmod6449_2_lbuf_25_11 , divmod6449_2_lbuf_24_11
        , divmod6449_2_lbuf_23_11 , divmod6449_2_lbuf_22_11 , divmod6449_2_lbuf_21_11
        , divmod6449_2_lbuf_20_11 , divmod6449_2_lbuf_19_11 , divmod6449_2_lbuf_18_11
        , divmod6449_2_lbuf_17_11 , divmod6449_2_lbuf_16_11 , divmod6449_2_lbuf_15_9
        , (divmod6449_2_lbuf_15_0_1[4])}) + ({1'b1 , (~ BUTTERFLY_i_div_cmp_b)})
        + 17'b00000000000000001;
    if ( divmod6449_2_diff_12[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_23_12 = divmod6449_2_diff_12[8];
      divmod6449_2_lbuf_22_12 = divmod6449_2_diff_12[7];
      divmod6449_2_lbuf_24_12 = divmod6449_2_diff_12[9];
      divmod6449_2_lbuf_21_12 = divmod6449_2_diff_12[6];
      divmod6449_2_lbuf_25_12 = divmod6449_2_diff_12[10];
      divmod6449_2_lbuf_20_12 = divmod6449_2_diff_12[5];
      divmod6449_2_lbuf_26_12 = divmod6449_2_diff_12[11];
      divmod6449_2_lbuf_19_12 = divmod6449_2_diff_12[4];
      divmod6449_2_lbuf_18_12 = divmod6449_2_diff_12[3];
      divmod6449_2_lbuf_17_12 = divmod6449_2_diff_12[2];
      divmod6449_2_lbuf_16_12 = divmod6449_2_diff_12[1];
      divmod6449_2_lbuf_15_10 = divmod6449_2_diff_12[0];
    end
    divmod6449_2_lbuf_27_13 = divmod6449_2_lbuf_26_12;
    divmod6449_2_lbuf_26_13 = divmod6449_2_lbuf_25_12;
    divmod6449_2_lbuf_25_13 = divmod6449_2_lbuf_24_12;
    divmod6449_2_lbuf_24_13 = divmod6449_2_lbuf_23_12;
    divmod6449_2_lbuf_23_13 = divmod6449_2_lbuf_22_12;
    divmod6449_2_lbuf_22_13 = divmod6449_2_lbuf_21_12;
    divmod6449_2_lbuf_21_13 = divmod6449_2_lbuf_20_12;
    divmod6449_2_lbuf_20_13 = divmod6449_2_lbuf_19_12;
    divmod6449_2_lbuf_19_13 = divmod6449_2_lbuf_18_12;
    divmod6449_2_lbuf_18_13 = divmod6449_2_lbuf_17_12;
    divmod6449_2_lbuf_17_13 = divmod6449_2_lbuf_16_12;
    divmod6449_2_lbuf_16_13 = divmod6449_2_lbuf_15_10;
    divmod6449_2_lbuf_15_11 = divmod6449_2_lbuf_15_0_1[3];
    divmod6449_2_diff_13 = conv_u2u_13_17({divmod6449_2_lbuf_26_12 , divmod6449_2_lbuf_25_12
        , divmod6449_2_lbuf_24_12 , divmod6449_2_lbuf_23_12 , divmod6449_2_lbuf_22_12
        , divmod6449_2_lbuf_21_12 , divmod6449_2_lbuf_20_12 , divmod6449_2_lbuf_19_12
        , divmod6449_2_lbuf_18_12 , divmod6449_2_lbuf_17_12 , divmod6449_2_lbuf_16_12
        , divmod6449_2_lbuf_15_10 , (divmod6449_2_lbuf_15_0_1[3])}) + ({1'b1 , (~
        BUTTERFLY_i_div_cmp_b)}) + 17'b00000000000000001;
    if ( divmod6449_2_diff_13[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_23_13 = divmod6449_2_diff_13[8];
      divmod6449_2_lbuf_22_13 = divmod6449_2_diff_13[7];
      divmod6449_2_lbuf_24_13 = divmod6449_2_diff_13[9];
      divmod6449_2_lbuf_21_13 = divmod6449_2_diff_13[6];
      divmod6449_2_lbuf_25_13 = divmod6449_2_diff_13[10];
      divmod6449_2_lbuf_20_13 = divmod6449_2_diff_13[5];
      divmod6449_2_lbuf_26_13 = divmod6449_2_diff_13[11];
      divmod6449_2_lbuf_19_13 = divmod6449_2_diff_13[4];
      divmod6449_2_lbuf_27_13 = divmod6449_2_diff_13[12];
      divmod6449_2_lbuf_18_13 = divmod6449_2_diff_13[3];
      divmod6449_2_lbuf_17_13 = divmod6449_2_diff_13[2];
      divmod6449_2_lbuf_16_13 = divmod6449_2_diff_13[1];
      divmod6449_2_lbuf_15_11 = divmod6449_2_diff_13[0];
    end
    divmod6449_2_lbuf_28_14 = divmod6449_2_lbuf_27_13;
    divmod6449_2_lbuf_27_14 = divmod6449_2_lbuf_26_13;
    divmod6449_2_lbuf_26_14 = divmod6449_2_lbuf_25_13;
    divmod6449_2_lbuf_25_14 = divmod6449_2_lbuf_24_13;
    divmod6449_2_lbuf_24_14 = divmod6449_2_lbuf_23_13;
    divmod6449_2_lbuf_23_14 = divmod6449_2_lbuf_22_13;
    divmod6449_2_lbuf_22_14 = divmod6449_2_lbuf_21_13;
    divmod6449_2_lbuf_21_14 = divmod6449_2_lbuf_20_13;
    divmod6449_2_lbuf_20_14 = divmod6449_2_lbuf_19_13;
    divmod6449_2_lbuf_19_14 = divmod6449_2_lbuf_18_13;
    divmod6449_2_lbuf_18_14 = divmod6449_2_lbuf_17_13;
    divmod6449_2_lbuf_17_14 = divmod6449_2_lbuf_16_13;
    divmod6449_2_lbuf_16_14 = divmod6449_2_lbuf_15_11;
    divmod6449_2_lbuf_15_12 = divmod6449_2_lbuf_15_0_1[2];
    divmod6449_2_diff_14 = conv_u2u_14_17({divmod6449_2_lbuf_27_13 , divmod6449_2_lbuf_26_13
        , divmod6449_2_lbuf_25_13 , divmod6449_2_lbuf_24_13 , divmod6449_2_lbuf_23_13
        , divmod6449_2_lbuf_22_13 , divmod6449_2_lbuf_21_13 , divmod6449_2_lbuf_20_13
        , divmod6449_2_lbuf_19_13 , divmod6449_2_lbuf_18_13 , divmod6449_2_lbuf_17_13
        , divmod6449_2_lbuf_16_13 , divmod6449_2_lbuf_15_11 , (divmod6449_2_lbuf_15_0_1[2])})
        + ({1'b1 , (~ BUTTERFLY_i_div_cmp_b)}) + 17'b00000000000000001;
    if ( divmod6449_2_diff_14[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_23_14 = divmod6449_2_diff_14[8];
      divmod6449_2_lbuf_22_14 = divmod6449_2_diff_14[7];
      divmod6449_2_lbuf_24_14 = divmod6449_2_diff_14[9];
      divmod6449_2_lbuf_21_14 = divmod6449_2_diff_14[6];
      divmod6449_2_lbuf_25_14 = divmod6449_2_diff_14[10];
      divmod6449_2_lbuf_20_14 = divmod6449_2_diff_14[5];
      divmod6449_2_lbuf_26_14 = divmod6449_2_diff_14[11];
      divmod6449_2_lbuf_19_14 = divmod6449_2_diff_14[4];
      divmod6449_2_lbuf_27_14 = divmod6449_2_diff_14[12];
      divmod6449_2_lbuf_18_14 = divmod6449_2_diff_14[3];
      divmod6449_2_lbuf_28_14 = divmod6449_2_diff_14[13];
      divmod6449_2_lbuf_17_14 = divmod6449_2_diff_14[2];
      divmod6449_2_lbuf_16_14 = divmod6449_2_diff_14[1];
      divmod6449_2_lbuf_15_12 = divmod6449_2_diff_14[0];
    end
    divmod6449_2_lbuf_29_15 = divmod6449_2_lbuf_28_14;
    divmod6449_2_lbuf_28_15 = divmod6449_2_lbuf_27_14;
    divmod6449_2_lbuf_27_15 = divmod6449_2_lbuf_26_14;
    divmod6449_2_lbuf_26_15 = divmod6449_2_lbuf_25_14;
    divmod6449_2_lbuf_25_15 = divmod6449_2_lbuf_24_14;
    divmod6449_2_lbuf_24_15 = divmod6449_2_lbuf_23_14;
    divmod6449_2_lbuf_23_15 = divmod6449_2_lbuf_22_14;
    divmod6449_2_lbuf_22_15 = divmod6449_2_lbuf_21_14;
    divmod6449_2_lbuf_21_15 = divmod6449_2_lbuf_20_14;
    divmod6449_2_lbuf_20_15 = divmod6449_2_lbuf_19_14;
    divmod6449_2_lbuf_19_15 = divmod6449_2_lbuf_18_14;
    divmod6449_2_lbuf_18_15 = divmod6449_2_lbuf_17_14;
    divmod6449_2_lbuf_17_15 = divmod6449_2_lbuf_16_14;
    divmod6449_2_lbuf_16_15 = divmod6449_2_lbuf_15_12;
    divmod6449_2_lbuf_15_13 = divmod6449_2_lbuf_15_0_1[1];
    divmod6449_2_diff_15 = conv_u2u_15_17({divmod6449_2_lbuf_28_14 , divmod6449_2_lbuf_27_14
        , divmod6449_2_lbuf_26_14 , divmod6449_2_lbuf_25_14 , divmod6449_2_lbuf_24_14
        , divmod6449_2_lbuf_23_14 , divmod6449_2_lbuf_22_14 , divmod6449_2_lbuf_21_14
        , divmod6449_2_lbuf_20_14 , divmod6449_2_lbuf_19_14 , divmod6449_2_lbuf_18_14
        , divmod6449_2_lbuf_17_14 , divmod6449_2_lbuf_16_14 , divmod6449_2_lbuf_15_12
        , (divmod6449_2_lbuf_15_0_1[1])}) + ({1'b1 , (~ BUTTERFLY_i_div_cmp_b)})
        + 17'b00000000000000001;
    if ( divmod6449_2_diff_15[16] ) begin
    end
    else begin
      divmod6449_2_lbuf_23_15 = divmod6449_2_diff_15[8];
      divmod6449_2_lbuf_22_15 = divmod6449_2_diff_15[7];
      divmod6449_2_lbuf_24_15 = divmod6449_2_diff_15[9];
      divmod6449_2_lbuf_21_15 = divmod6449_2_diff_15[6];
      divmod6449_2_lbuf_25_15 = divmod6449_2_diff_15[10];
      divmod6449_2_lbuf_20_15 = divmod6449_2_diff_15[5];
      divmod6449_2_lbuf_26_15 = divmod6449_2_diff_15[11];
      divmod6449_2_lbuf_19_15 = divmod6449_2_diff_15[4];
      divmod6449_2_lbuf_27_15 = divmod6449_2_diff_15[12];
      divmod6449_2_lbuf_18_15 = divmod6449_2_diff_15[3];
      divmod6449_2_lbuf_28_15 = divmod6449_2_diff_15[13];
      divmod6449_2_lbuf_17_15 = divmod6449_2_diff_15[2];
      divmod6449_2_lbuf_29_15 = divmod6449_2_diff_15[14];
      divmod6449_2_lbuf_16_15 = divmod6449_2_diff_15[1];
      divmod6449_2_lbuf_15_13 = divmod6449_2_diff_15[0];
    end
    BUTTERFLY_i_div_cmp_z_7 = ~ (divmod6449_2_diff_9[16]);
    BUTTERFLY_i_div_cmp_z_8 = ~ (divmod6449_2_diff_8[16]);
    BUTTERFLY_i_div_cmp_z_6 = ~ (divmod6449_2_diff_10[16]);
    BUTTERFLY_i_div_cmp_z_9 = ~ (divmod6449_2_diff_7[16]);
    BUTTERFLY_i_div_cmp_z_5 = ~ (divmod6449_2_diff_11[16]);
    BUTTERFLY_i_div_cmp_z_10 = ~ (divmod6449_2_diff_6[16]);
    BUTTERFLY_i_div_cmp_z_4 = ~ (divmod6449_2_diff_12[16]);
    BUTTERFLY_i_div_cmp_z_11 = ~ (divmod6449_2_diff_5[16]);
    BUTTERFLY_i_div_cmp_z_3 = ~ (divmod6449_2_diff_13[16]);
    BUTTERFLY_i_div_cmp_z_12 = ~ (divmod6449_2_diff_4[16]);
    BUTTERFLY_i_div_cmp_z_2 = ~ (divmod6449_2_diff_14[16]);
    BUTTERFLY_i_div_cmp_z_13 = ~ (divmod6449_2_diff_3[16]);
    BUTTERFLY_i_div_cmp_z_1 = ~ (divmod6449_2_diff_15[16]);
    BUTTERFLY_i_div_cmp_z_14 = ~ (divmod6449_2_diff_2[16]);
    nl_divmod6449_2_loop951_16_acc_1_nl = conv_u2u_16_17({divmod6449_2_lbuf_29_15
        , divmod6449_2_lbuf_28_15 , divmod6449_2_lbuf_27_15 , divmod6449_2_lbuf_26_15
        , divmod6449_2_lbuf_25_15 , divmod6449_2_lbuf_24_15 , divmod6449_2_lbuf_23_15
        , divmod6449_2_lbuf_22_15 , divmod6449_2_lbuf_21_15 , divmod6449_2_lbuf_20_15
        , divmod6449_2_lbuf_19_15 , divmod6449_2_lbuf_18_15 , divmod6449_2_lbuf_17_15
        , divmod6449_2_lbuf_16_15 , divmod6449_2_lbuf_15_13 , (divmod6449_2_lbuf_15_0_1[0])})
        + ({1'b1 , (~ BUTTERFLY_i_div_cmp_b)}) + 17'b00000000000000001;
    divmod6449_2_loop951_16_acc_1_nl = nl_divmod6449_2_loop951_16_acc_1_nl[16:0];
    BUTTERFLY_i_div_cmp_z_0 = ~ (readslicef_17_1_16(divmod6449_2_loop951_16_acc_1_nl));
    BUTTERFLY_i_div_cmp_z_15 = ~ (divmod6449_2_diff_1[16]);
  end


  function automatic [0:0] readslicef_17_1_16;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_17_1_16 = tmp[0:0];
  end
  endfunction


  function automatic [16:0] conv_u2u_1_17 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_17 = {{16{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_2_17 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_17 = {{15{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_3_17 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_17 = {{14{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_4_17 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_17 = {{13{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_5_17 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_17 = {{12{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_6_17 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_17 = {{11{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_7_17 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_17 = {{10{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_8_17 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_17 = {{9{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_9_17 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_17 = {{8{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_10_17 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_17 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_11_17 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_17 = {{6{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_12_17 ;
    input [11:0]  vector ;
  begin
    conv_u2u_12_17 = {{5{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_13_17 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_17 = {{4{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_14_17 ;
    input [13:0]  vector ;
  begin
    conv_u2u_14_17 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_15_17 ;
    input [14:0]  vector ;
  begin
    conv_u2u_15_17 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_17 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage
// ------------------------------------------------------------------


module stage (
  clk, rst, arst_n, ap_start_rsc_dat, ap_start_rsc_vld, ap_start_rsc_rdy, ap_done_rsc_dat,
      ap_done_rsc_vld, ap_done_rsc_rdy, mode1_rsc_dat, mode1_triosy_lz, in_f_d_rsc_adr,
      in_f_d_rsc_d, in_f_d_rsc_we, in_f_d_rsc_q, in_f_d_rsc_en, in_f_d_triosy_lz,
      in_u_rsc_adr, in_u_rsc_d, in_u_rsc_we, in_u_rsc_q, in_u_rsc_en, in_u_triosy_lz,
      out_f_d_rsc_adr, out_f_d_rsc_d, out_f_d_rsc_we, out_f_d_rsc_q, out_f_d_rsc_en,
      out_f_d_triosy_lz, out_u_rsc_adr, out_u_rsc_d, out_u_rsc_we, out_u_rsc_q, out_u_rsc_en,
      out_u_triosy_lz, out1_rsc_dat, out1_rsc_vld, out1_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input [15:0] mode1_rsc_dat;
  output mode1_triosy_lz;
  output [9:0] in_f_d_rsc_adr;
  output [63:0] in_f_d_rsc_d;
  output in_f_d_rsc_we;
  input [63:0] in_f_d_rsc_q;
  output in_f_d_rsc_en;
  output in_f_d_triosy_lz;
  output [9:0] in_u_rsc_adr;
  output [15:0] in_u_rsc_d;
  output in_u_rsc_we;
  input [15:0] in_u_rsc_q;
  output in_u_rsc_en;
  output in_u_triosy_lz;
  output [9:0] out_f_d_rsc_adr;
  output [63:0] out_f_d_rsc_d;
  output out_f_d_rsc_we;
  input [63:0] out_f_d_rsc_q;
  output out_f_d_rsc_en;
  output out_f_d_triosy_lz;
  output [9:0] out_u_rsc_adr;
  output [15:0] out_u_rsc_d;
  output out_u_rsc_we;
  input [15:0] out_u_rsc_q;
  output out_u_rsc_en;
  output out_u_triosy_lz;
  output [79:0] out1_rsc_dat;
  output out1_rsc_vld;
  input out1_rsc_rdy;


  // Interconnect Declarations
  wire [15:0] out1_rsc_dat_u;
  wire [63:0] out1_rsc_dat_d;


  // Interconnect Declarations for Component Instantiations 
  stage_struct stage_struct_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .ap_start_rsc_dat(ap_start_rsc_dat),
      .ap_start_rsc_vld(ap_start_rsc_vld),
      .ap_start_rsc_rdy(ap_start_rsc_rdy),
      .ap_done_rsc_dat(ap_done_rsc_dat),
      .ap_done_rsc_vld(ap_done_rsc_vld),
      .ap_done_rsc_rdy(ap_done_rsc_rdy),
      .mode1_rsc_dat(mode1_rsc_dat),
      .mode1_triosy_lz(mode1_triosy_lz),
      .in_f_d_rsc_adr(in_f_d_rsc_adr),
      .in_f_d_rsc_d(in_f_d_rsc_d),
      .in_f_d_rsc_we(in_f_d_rsc_we),
      .in_f_d_rsc_q(in_f_d_rsc_q),
      .in_f_d_rsc_en(in_f_d_rsc_en),
      .in_f_d_triosy_lz(in_f_d_triosy_lz),
      .in_u_rsc_adr(in_u_rsc_adr),
      .in_u_rsc_d(in_u_rsc_d),
      .in_u_rsc_we(in_u_rsc_we),
      .in_u_rsc_q(in_u_rsc_q),
      .in_u_rsc_en(in_u_rsc_en),
      .in_u_triosy_lz(in_u_triosy_lz),
      .out_f_d_rsc_adr(out_f_d_rsc_adr),
      .out_f_d_rsc_d(out_f_d_rsc_d),
      .out_f_d_rsc_we(out_f_d_rsc_we),
      .out_f_d_rsc_q(out_f_d_rsc_q),
      .out_f_d_rsc_en(out_f_d_rsc_en),
      .out_f_d_triosy_lz(out_f_d_triosy_lz),
      .out_u_rsc_adr(out_u_rsc_adr),
      .out_u_rsc_d(out_u_rsc_d),
      .out_u_rsc_we(out_u_rsc_we),
      .out_u_rsc_q(out_u_rsc_q),
      .out_u_rsc_en(out_u_rsc_en),
      .out_u_triosy_lz(out_u_triosy_lz),
      .out1_rsc_dat_u(out1_rsc_dat_u),
      .out1_rsc_dat_d(out1_rsc_dat_d),
      .out1_rsc_vld(out1_rsc_vld),
      .out1_rsc_rdy(out1_rsc_rdy)
    );
  assign out1_rsc_dat = {out1_rsc_dat_u , out1_rsc_dat_d};
endmodule



