module USER_PRJ1 #( parameter pUSER_PROJECT_SIDEBAND_WIDTH   = 5,
          parameter pADDR_WIDTH   = 12,
                   parameter pDATA_WIDTH   = 32
                 )
(
  output wire                        awready,
  output wire                        arready,
  output wire                        wready,
  output wire                        rvalid,
  output wire  [(pDATA_WIDTH-1) : 0] rdata,
  input  wire                        awvalid,
  input  wire                [11: 0] awaddr,
  input  wire                        arvalid,
  input  wire                [11: 0] araddr,
  input  wire                        wvalid,
  input  wire                 [3: 0] wstrb,
  input  wire  [(pDATA_WIDTH-1) : 0] wdata,
  input  wire                        rready,
  input  wire                        ss_tvalid,
  input  wire  [(pDATA_WIDTH-1) : 0] ss_tdata,
  input  wire                 [1: 0] ss_tuser,
    `ifdef USER_PROJECT_SIDEBAND_SUPPORT
  input  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] ss_tupsb,
  `endif
  input  wire                 [3: 0] ss_tstrb,
  input  wire                 [3: 0] ss_tkeep,
  input  wire                        ss_tlast,
  input  wire                        sm_tready,
  output wire                        ss_tready,
  output wire                        sm_tvalid,
  output wire  [(pDATA_WIDTH-1) : 0] sm_tdata,
  output wire                 [2: 0] sm_tid,
  `ifdef USER_PROJECT_SIDEBAND_SUPPORT
  output  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] sm_tupsb,
  `endif
  output wire                 [3: 0] sm_tstrb,
  output wire                 [3: 0] sm_tkeep,
  output wire                        sm_tlast,
  output wire                        low__pri_irq,
  output wire                        High_pri_req,
  output wire                [23: 0] la_data_o,
  input  wire                        axi_clk,
  input  wire                        axis_clk,
  input  wire                        axi_reset_n,
  input  wire                        axis_rst_n,
  input  wire                        user_clock2,
  input  wire                        uck2_rst_n
);

////////////////////////// axi- lite part


wire awvalid_in;
wire wvalid_in;

//write addr channel
assign awvalid_in	= awvalid; 
wire awready_out;
assign awready = awready_out;

//write data channel
assign 	wvalid_in	= wvalid;
wire wready_out;
assign wready = wready_out;

// if both awvalid_in=1 and wvalid_in=1 then output awready_out = 1 and wready_out = 1
assign awready_out = (awvalid_in && wvalid_in) ? 1 : 0;
assign wready_out = (awvalid_in && wvalid_in) ? 1 : 0;

wire ss_tready_out;
assign ss_tready=ss_tready_out;


wire sm_tvalid_out;
assign sm_tvalid = sm_tvalid_out;

wire [31:0] sm_tdata_out;
assign sm_tdata  = sm_tdata_out;

//write register   // to let RESET State go back to Command state
/*always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) begin
    reg_ap_control         <= 0;

  end else begin
    if ( awvalid_in && wvalid_in ) begin		//when awvalid_in=1 and wvalid_in=1 means awready_out=1 and wready_out=1
       if  (awaddr[11:0] == 12'h000 ) begin //offset 0
      
       end 
       else begin
       end
    end
  end
end
*/
localparam	RD_IDLE = 1'b0;
localparam	RD_ADDR_DONE = 1'b1;
localparam	Command   = 4'd0;
localparam	IN_COPY   = 4'd1;
localparam	OUT_COPY  = 4'd2;
localparam	RESET     = 4'd3;
localparam	F_WAIT1    = 4'd1;
localparam	F_OUT1     = 4'd2;
localparam	F_OUT2     = 4'd3;
localparam	U_OUT      = 4'd4;
reg [3:0] state,next_state;
//read register
reg [(pDATA_WIDTH-1) : 0] rdata_tmp;
assign arready = 1; //always assigned to 1, limitation: only support 1T in arvalid, if master issue 2T in arvalid then only 1st raddr is captured.
reg rvalid_out ;
assign rvalid = rvalid_out;
assign rdata =  rdata_tmp;
reg rd_state;
reg rd_next_state;
reg [pADDR_WIDTH-1:0] rd_addr;
reg [3:0] Out_state,next_Out_state;
////
always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) 
    rd_state <= RD_IDLE;
  else
    rd_state <= rd_next_state;
end



always@(*)begin
  case(rd_state)
    RD_IDLE:
      if(arvalid && arready) rd_next_state = RD_ADDR_DONE;
      else      rd_next_state = RD_IDLE;
    RD_ADDR_DONE:
      if(rready && rvalid_out) rd_next_state = RD_IDLE;
      else    rd_next_state = RD_ADDR_DONE;
    default:rd_next_state = RD_IDLE;
  endcase
end 

always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) begin
        rd_addr <= 0;
	      rvalid_out <= 0;
  end	
  else begin
    if (rd_state == RD_IDLE )
	  if(arvalid && arready) begin
		rd_addr <= araddr;
		rvalid_out <= 1;
	  end	
	if (rd_state == RD_ADDR_DONE ) 
	  if(rready && rvalid_out)
		rvalid_out <= 0;
  end	
end

////
always @* begin
  if      (rd_addr[11:0] == 12'h000) rdata_tmp = (state==RESET);
  else                               rdata_tmp = 0;
end


assign sm_tid        = 3'b0;
`ifdef USER_PROJECT_SIDEBAND_SUPPORT
  assign sm_tupsb      = 5'b0;
`endif
assign sm_tstrb      = 4'b0;
assign sm_tkeep      = 1'b0;
assign low__pri_irq  = 1'b0;
assign High_pri_req  = 1'b0;

// 24 bit 
// [23:16] for axi-lite interface; [15:12] for axi-stream interface; [11:8] for state; [7:4] for Out_state; [3:0] for data;
assign la_data_o[23:16] = {awvalid,awready_out,wvalid,wready_out,arvalid,1'b1,rready,rvalid_out};
assign la_data_o[15:12] = {ss_tvalid,ss_tready_out,sm_tvalid_out,sm_tready};
assign la_data_o[11:8]=state;
assign la_data_o[7:4]=Out_state;
assign la_data_o[3:0]={wdata[0],ss_tdata[0],sm_tdata_out[0],1'b0};

wire        in_ramf_en;
wire [63:0] in_ramf_q;
wire        in_ramf_we;
wire [63:0] in_ramf_d;
wire [9:0]  in_ramf_adr;

wire        in_ramu_en;
wire [15:0] in_ramu_q;
wire        in_ramu_we;
wire [15:0] in_ramu_d;
wire [9:0]  in_ramu_adr;

wire        out_ramf_en;
wire [63:0] out_ramf_q;
wire        out_ramf_we;
wire [63:0] out_ramf_d;
wire [9:0]  out_ramf_adr;

wire        out_ramu_en;
wire [15:0] out_ramu_q;
wire        out_ramu_we;
wire [15:0] out_ramu_d;
wire [9:0]  out_ramu_adr;

wire        ram0_en;
wire [63:0] ram0_q;
wire        ram0_we;
wire [63:0] ram0_d;
wire [9:0]  ram0_adr;

wire        ram1_en;
wire [63:0] ram1_q;
wire        ram1_we;
wire [63:0] ram1_d;
wire [9:0]  ram1_adr;

wire [63:0] In_data;
wire In_vld;
wire In_rdy;	
wire [9:0] Inram_adr;
wire [63:0] Inram_d;
wire Inram_we;
reg reg_rst_incpopy;
reg reg_rst_out_stage;
reg [31:0]regx_data;
reg [31:0]regy_data;
reg [15:0]reg_mode1_in;

assign ss_tready_out=(state==Command)?1'b1:(state==IN_COPY)?In_rdy:1'b0;
assign In_vld=(state==IN_COPY)?ss_tvalid:1'b0;

In_copy In_copy (
  .clk(axi_clk), 
  .rst(reg_rst_incpopy), 
  .arst_n(axi_reset_n),
  .in_data_rsc_dat(ss_tdata),
  .in_data_rsc_vld(In_vld), //I
  .in_data_rsc_rdy(In_rdy), 
  .qin_rsc_adr(Inram_adr),
  .qin_rsc_d(Inram_d),
  .qin_rsc_we(Inram_we),
  .qin_rsc_q(),
  .qin_rsc_en(Inram_en),
  .qin_triosy_lz(),
  .ap_done_rsc_dat(), 
  .ap_done_rsc_vld(In_copy_done),
  .ap_done_rsc_rdy(1'b1),
  .ap_start_rsc_dat(1'b1),
  .ap_start_rsc_vld(state==IN_COPY),
  .ap_start_rsc_rdy(),
  .mode_rsc_dat(reg_mode1_in==2||reg_mode1_in==3)
);

wire ap_done_vld;     
wire ap_done_rdy;     

wire Out_vld;

always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) begin
    state <= 4'b0;
  end
  else begin
    state <= next_state;
  end
end

wire Out_copy_done;

always@(*)begin
  case(state)
    Command:   
    	if(ss_tvalid && ss_tdata[3:2]==2'b01) next_state = IN_COPY;
   		else next_state = Command;
    IN_COPY:   
    	if(In_copy_done) next_state = OUT_COPY;
   		else next_state = IN_COPY;
    OUT_COPY:  
    	if(Out_copy_done) next_state=RESET;
   		else next_state=OUT_COPY;
    RESET:
    	if(awvalid_in && wvalid_in &&(awaddr[11:0] == 12'h000)&&(wdata[0]==1)) next_state=Command;
     	else next_state = RESET;
    default:next_state = Command;
  endcase
end 

reg reg_rst;

always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) begin
    reg_mode1_in <= 16'b0;
  end
  else begin
    if(state==Command)begin
      reg_mode1_in <= {14'b0,ss_tdata[1:0]};
    end
    else begin
      reg_mode1_in <=reg_mode1_in;
    end
  end
end

always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) begin 
    Out_state <= 2'b0;
  end
  else begin
  	Out_state <= next_Out_state;
  end
end

always@(*)begin
  case(Out_state)
    Command: 
    	if(ss_tvalid && ss_tdata[3:2]==2'b01 && (ss_tdata[1:0]==2'd0 || ss_tdata[1:0]== 2'd1))  next_Out_state = F_WAIT1;
    	else if(ss_tvalid && ss_tdata[3:2]==2'b01 && (ss_tdata[1:0]==2'd2 || ss_tdata[1:0]==2'd3))  next_Out_state = U_OUT;
    	else next_Out_state=Command;
    	
    F_WAIT1:
    	if(Out_copy_done)next_Out_state = Command;
			else if(Out_vld)next_Out_state = F_OUT1;
    	else next_Out_state = F_WAIT1;
    	
    F_OUT1: 
    	if(sm_tready) next_Out_state = F_OUT2;
    	else next_Out_state = F_OUT1;
    	
    F_OUT2: 
    	if(sm_tready) next_Out_state = F_WAIT1;
    	else next_Out_state = F_OUT2;
    	
    U_OUT:    
    	if(Out_copy_done)next_Out_state = Command;
    	else next_Out_state = U_OUT;
    	
    default:next_Out_state=Command;
  endcase
end 

wire [79:0] Out_data;

always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) begin
		regx_data <= 32'b0;
		regy_data <= 32'b0;
  end
  else begin
  	if(Out_state==F_WAIT1 && Out_vld)begin
			regx_data <= Out_data[31:0];
			regy_data <= Out_data[63:32];
 	  end
 	  else begin
      regx_data <= regx_data;
			regy_data <= regy_data;
 	  end
  end
end

/********** sm_tlast ***********/

reg [11:0] last_cnt;
always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) begin
		last_cnt <= 12'b0;
  end
  else begin
    if(state==RESET) last_cnt <= 12'b0;
    else begin
      if(((Out_state==U_OUT) ? Out_vld : (Out_state==F_OUT1||Out_state==F_OUT2))&sm_tready) last_cnt<=last_cnt+12'b1;
      else last_cnt<=last_cnt;
 	  end
  end
end




assign sm_tlast  = (reg_mode1_in[1])  ? ((last_cnt==12'd1023) ? 1 : 0) : ((last_cnt==12'd2047) ? 1 : 0);
assign sm_tvalid_out=(Out_state==U_OUT) ? Out_vld : (Out_state==F_OUT1||Out_state==F_OUT2);
assign sm_tdata_out=(Out_state==U_OUT) ? {16'b0,Out_data[79:64]} : ((Out_state==F_OUT1)?regx_data:regy_data);
assign Out_rdy   = (Out_state==U_OUT||Out_state==F_OUT2) ? sm_tready : 0;




fiFFNTT fiFFNTT(
.clk(axi_clk),          // I
.rst(reg_rst),          // I
.arst_n(axi_reset_n),   // I
.ap_start_rsc_dat(1'b1),// I
.ap_start_rsc_vld(state==OUT_COPY),    // I
.ap_start_rsc_rdy(),    // O
.ap_done_rsc_dat(),     // O
.ap_done_rsc_vld(Out_copy_done), // O
.ap_done_rsc_rdy(1'b1),     // I
.mode1_rsc_dat(reg_mode1_in),  //I 16
.mode1_triosy_lz(), 
.in_f_d_rsc_adr(in_ramf_adr),  // O 10
.in_f_d_rsc_d(in_ramf_d),    // O 64
.in_f_d_rsc_we(in_ramf_we),   // O 1 
.in_f_d_rsc_q(in_ramf_q),    // I 64
.in_f_d_rsc_en(in_ramf_en),   // O 1
.in_f_d_triosy_lz(), 
.in_u_rsc_adr(in_ramu_adr), // O 10
.in_u_rsc_d(in_ramu_d),   // O 16
.in_u_rsc_we(in_ramu_we),  // O
.in_u_rsc_q(in_ramu_q),   // I 16
.in_u_rsc_en(in_ramu_en),  // O 
.in_u_triosy_lz(),
.out_f_d_rsc_adr(out_ramf_adr),
.out_f_d_rsc_d(out_ramf_d),
.out_f_d_rsc_we(out_ramf_we),
.out_f_d_rsc_q(out_ramf_q), 
.out_f_d_rsc_en(out_ramf_en),
.out_f_d_triosy_lz(),
.out_u_rsc_adr(out_ramu_adr), 
.out_u_rsc_d(out_ramu_d),
.out_u_rsc_we(out_ramu_we), 
.out_u_rsc_q(out_ramu_q),
.out_u_rsc_en(out_ramu_en),
.out_u_triosy_lz(),
.out1_rsc_dat(Out_data),//O,80 bit{16'b,64'b},
.out1_rsc_vld(Out_vld),//O;
.out1_rsc_rdy(Out_rdy)
);






wire mux_state;
assign mux_state=!(reg_mode1_in==2||reg_mode1_in==3);
assign ram0_en   = (state==IN_COPY)?Inram_en  : ((mux_state)? in_ramf_en:in_ramu_en);
assign ram0_we   = (state==IN_COPY)?Inram_we  : ((mux_state)? in_ramf_we:in_ramu_we);
assign ram0_adr  = (state==IN_COPY)?Inram_adr : ((mux_state)? in_ramf_adr:in_ramu_adr);
assign ram0_d    = (state==IN_COPY)?Inram_d   : ((mux_state)? in_ramf_d:{48'b0,in_ramu_d});
assign in_ramu_q = ram0_q[15:0];
assign in_ramf_q = ram0_q;


assign ram1_en  	= (mux_state) ? out_ramf_en  : out_ramu_en;
assign ram1_we  	= (mux_state) ? out_ramf_we  : out_ramu_we;
assign ram1_adr 	= (mux_state) ? out_ramf_adr : out_ramu_adr;
assign ram1_d   	= (mux_state) ? out_ramf_d   : {48'b0,out_ramu_d};
assign out_ramu_q = ram1_q[15:0];
assign out_ramf_q = ram1_q;
`ifdef USE_PDK_SRAM
ralshd1024x64m4h3v2 SRAM0(
  .CLK(axi_clk),
  .WEN(~ram0_we),
  .OEN(1'b0),
  .CEN(~ram0_en),
  .A(ram0_adr),
  .D(ram0_d),
  .Q(ram0_q)
);

ralshd1024x64m4h3v2 SRAM1(
  .CLK(axi_clk),
  .WEN(~ram1_we),
  .OEN(1'b0),
  .CEN(~ram1_en),
  .A(ram1_adr),
  .D(ram1_d),
  .Q(ram1_q)
);

`else
SRAM1RW1024x8 S1(
.CE(axi_clk),
.WEB(~ram0_we),
.OEB(1'b0),
.CSB(~ram0_en),

.A(ram0_adr),
.I(ram0_d[7:0]),
.O(ram0_q[7:0])
);
SRAM1RW1024x8 S2(
.CE(axi_clk),
.WEB(~ram0_we),
.OEB(1'b0),
.CSB(~ram0_en),

.A(ram0_adr),
.I(ram0_d[15:8]),
.O(ram0_q[15:8])
);

SRAM1RW1024x8 S3(
.CE(axi_clk),
.WEB(~ram0_we),
.OEB(1'b0),
.CSB(~ram0_en),

.A(ram0_adr),
.I(ram0_d[23:16]),
.O(ram0_q[23:16])
);

SRAM1RW1024x8 S4(
.CE(axi_clk),
.WEB(~ram0_we),
.OEB(1'b0),
.CSB(~ram0_en),

.A(ram0_adr),
.I(ram0_d[31:24]),
.O(ram0_q[31:24])
);

SRAM1RW1024x8 S5(
.CE(axi_clk),
.WEB(~ram0_we),
.OEB(1'b0),
.CSB(~ram0_en),

.A(ram0_adr),
.I(ram0_d[39:32]),
.O(ram0_q[39:32])
);

SRAM1RW1024x8 S6(
.CE(axi_clk),
.WEB(~ram0_we),
.OEB(1'b0),
.CSB(~ram0_en),

.A(ram0_adr),
.I(ram0_d[47:40]),
.O(ram0_q[47:40])
);


SRAM1RW1024x8 S7(
.CE(axi_clk),
.WEB(~ram0_we),
.OEB(1'b0),
.CSB(~ram0_en),

.A(ram0_adr),
.I(ram0_d[55:48]),
.O(ram0_q[55:48])
);

SRAM1RW1024x8 S8(
.CE(axi_clk),
.WEB(~ram0_we),
.OEB(1'b0),
.CSB(~ram0_en),

.A(ram0_adr),
.I(ram0_d[63:56]),
.O(ram0_q[63:56])
);



SRAM1RW1024x8 S11(
.CE(axi_clk),
.WEB(~ram1_we),
.OEB(1'b0),
.CSB(~ram1_en),

.A(ram1_adr),
.I(ram1_d[7:0]),
.O(ram1_q[7:0])
);
SRAM1RW1024x8 S12(
.CE(axi_clk),
.WEB(~ram1_we),
.OEB(1'b0),
.CSB(~ram1_en),

.A(ram1_adr),
.I(ram1_d[15:8]),
.O(ram1_q[15:8])
);

SRAM1RW1024x8 S13(
.CE(axi_clk),
.WEB(~ram1_we),
.OEB(1'b0),
.CSB(~ram1_en),

.A(ram1_adr),
.I(ram1_d[23:16]),
.O(ram1_q[23:16])
);

SRAM1RW1024x8 S14(
.CE(axi_clk),
.WEB(~ram1_we),
.OEB(1'b0),
.CSB(~ram1_en),

.A(ram1_adr),
.I(ram1_d[31:24]),
.O(ram1_q[31:24])
);

SRAM1RW1024x8 S15(
.CE(axi_clk),
.WEB(~ram1_we),
.OEB(1'b0),
.CSB(~ram1_en),

.A(ram1_adr),
.I(ram1_d[39:32]),
.O(ram1_q[39:32])
);

SRAM1RW1024x8 S16(
.CE(axi_clk),
.WEB(~ram1_we),
.OEB(1'b0),
.CSB(~ram1_en),

.A(ram1_adr),
.I(ram1_d[47:40]),
.O(ram1_q[47:40])
);


SRAM1RW1024x8 S17(
.CE(axi_clk),
.WEB(~ram1_we),
.OEB(1'b0),
.CSB(~ram1_en),

.A(ram1_adr),
.I(ram1_d[55:48]),
.O(ram1_q[55:48])
);

SRAM1RW1024x8 S18(
.CE(axi_clk),
.WEB(~ram1_we),
.OEB(1'b0),
.CSB(~ram1_en),

.A(ram1_adr),
.I(ram1_d[63:56]),
.O(ram1_q[63:56])
);
`endif
endmodule 


`define numAddr 10
`define numWords 1024
`define wordLength 8


module SRAM1RW1024x8 (A,CE,WEB,OEB,CSB,I,O);

input 				CE;
input 				WEB;
input 				OEB;
input 				CSB;

input 	[`numAddr-1:0] 		A;
input 	[`wordLength-1:0] 	I;
output 	[`wordLength-1:0] 	O;

/*reg   [`wordLength-1:0]   	memory[`numWords-1:0];*/
/*reg  	[`wordLength-1:0]	data_out;*/
wire 	[`wordLength-1:0] 	O;

wire 				RE;
wire 				WE;

SRAM1RW1024x8_1bit sram_IO0 ( CE, WEB,  A, OEB, CSB, I[0], O[0]);
SRAM1RW1024x8_1bit sram_IO1 ( CE, WEB,  A, OEB, CSB, I[1], O[1]);
SRAM1RW1024x8_1bit sram_IO2 ( CE, WEB,  A, OEB, CSB, I[2], O[2]);
SRAM1RW1024x8_1bit sram_IO3 ( CE, WEB,  A, OEB, CSB, I[3], O[3]);
SRAM1RW1024x8_1bit sram_IO4 ( CE, WEB,  A, OEB, CSB, I[4], O[4]);
SRAM1RW1024x8_1bit sram_IO5 ( CE, WEB,  A, OEB, CSB, I[5], O[5]);
SRAM1RW1024x8_1bit sram_IO6 ( CE, WEB,  A, OEB, CSB, I[6], O[6]);
SRAM1RW1024x8_1bit sram_IO7 ( CE, WEB,  A, OEB, CSB, I[7], O[7]);


endmodule


module SRAM1RW1024x8_1bit (CE_i, WEB_i,  A_i, OEB_i, CSB_i, I_i, O_i);

input CSB_i;
input OEB_i;
input CE_i;
input WEB_i;

input 	[`numAddr-1:0] 	A_i;
input 	[0:0] I_i;

output 	[0:0] O_i;

reg 	[0:0]O_i;
reg    	[0:0]  	memory[`numWords-1:0];
reg  	[0:0]	data_out;


// Write Mode
and u1 (RE, ~CSB_i,  WEB_i);
and u2 (WE, ~CSB_i, ~WEB_i);


always @ (posedge CE_i) 
	if (RE)
		data_out = memory[A_i];
always @ (posedge CE_i) 
	if (WE)
		memory[A_i] = I_i;
		

always @ (data_out or OEB_i)
	if (!OEB_i) 
		O_i = data_out;
	else
		O_i =  1'bz;


endmodule
