//===========================================================
// Modified by Vic Chen
// Oct 5, 2024
//===========================================================

//`ifndef __GLOBAL_DEFINE_H
// Global parameters
`define __GLOBAL_DEFINE_H

`define MPRJ_IO_PADS_1 19	/* number of user GPIO pads on user1 side */
`define MPRJ_IO_PADS_2 19	/* number of user GPIO pads on user2 side */
`define MPRJ_IO_PADS (`MPRJ_IO_PADS_1 + `MPRJ_IO_PADS_2)

`define MPRJ_PWR_PADS_1 2	/* vdda1, vccd1 enable/disable control */
`define MPRJ_PWR_PADS_2 2	/* vdda2, vccd2 enable/disable control */
`define MPRJ_PWR_PADS (`MPRJ_PWR_PADS_1 + `MPRJ_PWR_PADS_2)

// Analog pads are only used by the "caravan" module and associated
// modules such as user_analog_project_wrapper and chip_io_alt.

`define ANALOG_PADS_1 5
`define ANALOG_PADS_2 6

`define ANALOG_PADS (`ANALOG_PADS_1 + `ANALOG_PADS_2)

// Number of GPIO pads defined in the caravel openframe layout
`define OPENFRAME_IO_PADS 44

// Size of soc_mem_synth

// Type and size of soc_mem
// `define USE_OPENRAM
`define USE_CUSTOM_DFFRAM
// don't change the following without double checking addr widths
`define MEM_WORDS 256

// Number of columns in the custom memory; takes one of three values:
// 1 column : 1 KB, 2 column: 2 KB, 4 column: 4KB
`define DFFRAM_WSIZE 4
`define DFFRAM_USE_LATCH 0

// not really parameterized but just to easily keep track of the number
// of ram_block across different modules
`define RAM_BLOCKS 1

// Clock divisor default value
`define CLK_DIV 3'b010

// GPIO control default mode and enable for most I/Os
// Most I/Os set to be user input pins on startup.
// NOTE:  To be modified, with GPIOs 5 to 35 being set from a build-time-
// programmable block.
`define MGMT_INIT 1'b0
`define OENB_INIT 1'b0
`define DM_INIT 3'b001

//`define TOP_ROUTING 1
`define REMOVE_LEVEL_SHIFT   1 //tony_debug
`define NO_POR_PAD 1 //tony_debug
`define REMOVE_sky130_ef_sc_hd__decap_12 1 //tony_debug
`define REMOVE_sky130_ef_io__corner_pad 1 //tony_debug
`define REMOVE_spare_logic_block 1 //tony_debug
`define REMOVE_sky130_fd_sc_hd__macro_sparecell 1 //tony_debug
`define SINGLE_POWER_DOMAIN 1 //tony_debug
`define REMOVE_PLL 1 //tony_debug
`define REMOVE_POWER_PAD //tony_debug
//`endif // __GLOBAL_DEFINE_H
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype wire

//`ifndef __USER_DEFINES_H
// User GPIO initial configuration parameters
`define __USER_DEFINES_H

// Useful GPIO mode values.  These match the names used in defs.h.
`define GPIO_MODE_MGMT_STD_INPUT_NOPULL    13'h0403
`define GPIO_MODE_MGMT_STD_INPUT_PULLDOWN  13'h0c01
`define GPIO_MODE_MGMT_STD_INPUT_PULLUP    13'h0801
`define GPIO_MODE_MGMT_STD_OUTPUT          13'h1809
`define GPIO_MODE_MGMT_STD_BIDIRECTIONAL   13'h1801
`define GPIO_MODE_MGMT_STD_ANALOG          13'h000b

`define GPIO_MODE_USER_STD_INPUT_NOPULL    13'h0402
`define GPIO_MODE_USER_STD_INPUT_PULLDOWN  13'h0c00
`define GPIO_MODE_USER_STD_INPUT_PULLUP    13'h0800
`define GPIO_MODE_USER_STD_OUTPUT          13'h1808
`define GPIO_MODE_USER_STD_BIDIRECTIONAL   13'h1800
`define GPIO_MODE_USER_STD_OUT_MONITORED   13'h1802
`define GPIO_MODE_USER_STD_ANALOG          13'h000a

// The power-on configuration for GPIO 0 to 4 is fixed and cannot be
// modified (allowing the SPI and debug to always be accessible unless
// overridden by a flash program).

// The values below can be any of the standard types defined above,
// or they can be any 13-bit value if the user wants a non-standard
// startup state for the GPIO.  By default, every GPIO from 5 to 37
// is set to power up as an input controlled by the management SoC.
// Users may want to redefine these so that the user project powers
// up in a state that can be used immediately without depending on
// the management SoC to run a startup program to configure the GPIOs.

`define USER_CONFIG_GPIO_5_INIT  `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_6_INIT  `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_7_INIT  `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_8_INIT  `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_9_INIT  `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_10_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_11_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_12_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_13_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL

// Configurations of GPIO 14 to 24 are used on caravel but not caravan.
`define USER_CONFIG_GPIO_14_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_15_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_16_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_17_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_18_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_19_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_20_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_21_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_22_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_23_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_24_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL

`define USER_CONFIG_GPIO_25_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_26_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_27_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_28_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_29_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_30_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_31_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_32_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_33_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_34_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_35_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_36_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL
`define USER_CONFIG_GPIO_37_INIT `GPIO_MODE_MGMT_STD_INPUT_NOPULL

//`endif // __USER_DEFINES_H
//===========================================================
// Author: Vic Chen
// Email: s179038@gmail.com
// Date:  Sep 27, 2024
//===========================================================
`default_nettype wire

// IO signal
//==========================
// 0:  mprj[0] - JTAG ---- I
// 1:  mprj[1] - SDO ----- O
// 2:  mprj[2] - SDI ----- I
// 3:  mprj[3] - CSB ----- I
// 4:  mprj[4] - SCK ----- I
// 5:  mprj[5] - ser_rx -- I
// 6:  mprj[6] - ser_tx -- O
// 7:  mprj[7] - irq ----- I
//--------------------------
// 8 ~ 21:
//     mprj[20:8] - RXD -- I
//     mprj[21] - RXCLK -- I
//--------------------------
// 22 ~ 35:
//     mprj[34:22] - TXD - O
//     mprj[35] - TXCLK -- O
//--------------------------
// 36: mprj[36] - IOCLK -- I
// 37: mprj[37] - NOTUSE - I
//==========================
// 38: clock ------------- I
// 39: flash_csb --------- O
// 40: flash_clk --------- O
// 41: flash_io0 --------- O
// 42: flash_io1 --------- I
// 43: gpio -------------- I

module pads_config (
    input         clk,
    input         resetb, // reset, active low
    // Wishbone Slave ports
    input         wb_clk_i,
    input         wb_rst_i,
    input         wbs_stb_i,
    input         wbs_cyc_i,
    input         wbs_we_i,
    input   [3:0] wbs_sel_i,
    input  [31:0] wbs_dat_i,
    input  [31:0] wbs_adr_i,
    output        wbs_ack_o,
    output [31:0] wbs_dat_o,
    // Output REN/OEN
    output        re_n,
    output [37:0] oe_n
);

    reg [37:0] r_OEN;
    reg        ACK;

    wire [37:0] cnfg_en; // Configure Enable
    wire        cnfg_decode; // Check target address
    wire        cnfg_vld;
  
    assign cnfg_decode = (wbs_adr_i[31:12] == 20'h3000_6)? 1'b1 : 1'b0;
    assign cnfg_vld = wbs_cyc_i & wbs_stb_i;

    assign wbs_ack_o = ACK;

    // Initially, set all ports to INPUT
    // Pull-up/down Resistor Enable: 0: Enable, 1: Disable
    // Reset period, force ren=0, i.e. enable pull-up/down resistors
    assign re_n = 1'b1 & resetb;
    generate
        genvar i;
        for (i = 0; i < 38; i = i + 1) begin : AND_RST_OEN
            assign oe_n[i] = r_OEN[i] | (~resetb);
        end
    endgenerate

    // Caravel FSIC initial IO state when reset
    always @(posedge clk or negedge resetb) begin
        if (~resetb) begin
            r_OEN[0]     <=   {{1'b1}};  // JTAG
            r_OEN[1]     <=   {{1'b0}};  // SDO
            r_OEN[5:2]   <=  {4{1'b1}};  // SDI, CSB, SCK, ser_rx
            r_OEN[6]     <=   {{1'b0}};  // ser_tx
            r_OEN[21:7]  <= {15{1'b1}};  // irq, RXD, RXCLK
            r_OEN[35:22] <= {14{1'b0}};  // TXD, TXCLK
            r_OEN[36]    <=   {{1'b1}};  // IOCLK
            r_OEN[37]    <=   {{1'b1}};  // mprj[37]
        end else begin
            integer i;
            for (i = 0; i < 38; i = i + 1) begin
                if (cnfg_en[i]) r_OEN[i] <= wbs_dat_i[0];
            end
        end
    end

    always @(posedge wb_clk_i or posedge wb_rst_i) begin
        if (wb_rst_i) begin
            ACK <= 0;
        end else begin
            if (cnfg_decode & cnfg_vld)
                ACK <= 1;
            else
                ACK <= 0;
        end
    end

    // WRITE
    assign cnfg_en[0]  = ((wbs_adr_i[7:0] == 8'h00) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[1]  = ((wbs_adr_i[7:0] == 8'h01) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[2]  = ((wbs_adr_i[7:0] == 8'h02) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[3]  = ((wbs_adr_i[7:0] == 8'h03) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[4]  = ((wbs_adr_i[7:0] == 8'h04) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[5]  = ((wbs_adr_i[7:0] == 8'h05) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[6]  = ((wbs_adr_i[7:0] == 8'h06) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[7]  = ((wbs_adr_i[7:0] == 8'h07) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[8]  = ((wbs_adr_i[7:0] == 8'h08) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[9]  = ((wbs_adr_i[7:0] == 8'h09) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[10] = ((wbs_adr_i[7:0] == 8'h0a) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[11] = ((wbs_adr_i[7:0] == 8'h0b) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[12] = ((wbs_adr_i[7:0] == 8'h0c) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[13] = ((wbs_adr_i[7:0] == 8'h0d) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[14] = ((wbs_adr_i[7:0] == 8'h0e) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[15] = ((wbs_adr_i[7:0] == 8'h0f) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[16] = ((wbs_adr_i[7:0] == 8'h10) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[17] = ((wbs_adr_i[7:0] == 8'h11) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[18] = ((wbs_adr_i[7:0] == 8'h12) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[19] = ((wbs_adr_i[7:0] == 8'h13) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[20] = ((wbs_adr_i[7:0] == 8'h14) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[21] = ((wbs_adr_i[7:0] == 8'h15) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[22] = ((wbs_adr_i[7:0] == 8'h16) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[23] = ((wbs_adr_i[7:0] == 8'h17) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[24] = ((wbs_adr_i[7:0] == 8'h18) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[25] = ((wbs_adr_i[7:0] == 8'h19) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[26] = ((wbs_adr_i[7:0] == 8'h1a) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[27] = ((wbs_adr_i[7:0] == 8'h1b) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[28] = ((wbs_adr_i[7:0] == 8'h1c) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[29] = ((wbs_adr_i[7:0] == 8'h1d) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[30] = ((wbs_adr_i[7:0] == 8'h1e) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[31] = ((wbs_adr_i[7:0] == 8'h1f) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[32] = ((wbs_adr_i[7:0] == 8'h20) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[33] = ((wbs_adr_i[7:0] == 8'h21) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[34] = ((wbs_adr_i[7:0] == 8'h22) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[35] = ((wbs_adr_i[7:0] == 8'h23) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[36] = ((wbs_adr_i[7:0] == 8'h24) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;
    assign cnfg_en[37] = ((wbs_adr_i[7:0] == 8'h25) && wbs_we_i & (cnfg_decode & cnfg_vld))? 1'b1 : 1'b0;

    // READ
    assign wbs_dat_o = ((wbs_adr_i[7:0] == 8'h00) && (!wbs_we_i))? r_OEN[0] :
                       ((wbs_adr_i[7:0] == 8'h01) && (!wbs_we_i))? r_OEN[1] :
                       ((wbs_adr_i[7:0] == 8'h02) && (!wbs_we_i))? r_OEN[2] :
                       ((wbs_adr_i[7:0] == 8'h03) && (!wbs_we_i))? r_OEN[3] :
                       ((wbs_adr_i[7:0] == 8'h04) && (!wbs_we_i))? r_OEN[4] :
                       ((wbs_adr_i[7:0] == 8'h05) && (!wbs_we_i))? r_OEN[5] :
                       ((wbs_adr_i[7:0] == 8'h06) && (!wbs_we_i))? r_OEN[6] :
                       ((wbs_adr_i[7:0] == 8'h07) && (!wbs_we_i))? r_OEN[7] :
                       ((wbs_adr_i[7:0] == 8'h08) && (!wbs_we_i))? r_OEN[8] :
                       ((wbs_adr_i[7:0] == 8'h09) && (!wbs_we_i))? r_OEN[9] :
                       ((wbs_adr_i[7:0] == 8'h0a) && (!wbs_we_i))? r_OEN[10] :
                       ((wbs_adr_i[7:0] == 8'h0b) && (!wbs_we_i))? r_OEN[11] :
                       ((wbs_adr_i[7:0] == 8'h0c) && (!wbs_we_i))? r_OEN[12] :
                       ((wbs_adr_i[7:0] == 8'h0d) && (!wbs_we_i))? r_OEN[13] :
                       ((wbs_adr_i[7:0] == 8'h0e) && (!wbs_we_i))? r_OEN[14] :
                       ((wbs_adr_i[7:0] == 8'h0f) && (!wbs_we_i))? r_OEN[15] :
                       ((wbs_adr_i[7:0] == 8'h10) && (!wbs_we_i))? r_OEN[16] :
                       ((wbs_adr_i[7:0] == 8'h11) && (!wbs_we_i))? r_OEN[17] :
                       ((wbs_adr_i[7:0] == 8'h12) && (!wbs_we_i))? r_OEN[18] :
                       ((wbs_adr_i[7:0] == 8'h13) && (!wbs_we_i))? r_OEN[19] :
                       ((wbs_adr_i[7:0] == 8'h14) && (!wbs_we_i))? r_OEN[20] :
                       ((wbs_adr_i[7:0] == 8'h15) && (!wbs_we_i))? r_OEN[21] :
                       ((wbs_adr_i[7:0] == 8'h16) && (!wbs_we_i))? r_OEN[22] :
                       ((wbs_adr_i[7:0] == 8'h17) && (!wbs_we_i))? r_OEN[23] :
                       ((wbs_adr_i[7:0] == 8'h18) && (!wbs_we_i))? r_OEN[24] :
                       ((wbs_adr_i[7:0] == 8'h19) && (!wbs_we_i))? r_OEN[25] :
                       ((wbs_adr_i[7:0] == 8'h1a) && (!wbs_we_i))? r_OEN[26] :
                       ((wbs_adr_i[7:0] == 8'h1b) && (!wbs_we_i))? r_OEN[27] :
                       ((wbs_adr_i[7:0] == 8'h1c) && (!wbs_we_i))? r_OEN[28] :
                       ((wbs_adr_i[7:0] == 8'h1d) && (!wbs_we_i))? r_OEN[29] :
                       ((wbs_adr_i[7:0] == 8'h1e) && (!wbs_we_i))? r_OEN[30] :
                       ((wbs_adr_i[7:0] == 8'h1f) && (!wbs_we_i))? r_OEN[31] :
                       ((wbs_adr_i[7:0] == 8'h20) && (!wbs_we_i))? r_OEN[32] :
                       ((wbs_adr_i[7:0] == 8'h21) && (!wbs_we_i))? r_OEN[33] :
                       ((wbs_adr_i[7:0] == 8'h22) && (!wbs_we_i))? r_OEN[34] :
                       ((wbs_adr_i[7:0] == 8'h23) && (!wbs_we_i))? r_OEN[35] :
                       ((wbs_adr_i[7:0] == 8'h24) && (!wbs_we_i))? r_OEN[36] :
                       ((wbs_adr_i[7:0] == 8'h25) && (!wbs_we_i))? r_OEN[37] :
                                                                   32'd0;

    
endmodule
module RAM256 #(parameter USE_LATCH = 1,
    WSIZE     = 4
)
(

    input   wire                 CLK,    // FO: 2
    input   wire [WSIZE-1:0]     WE0,     // FO: 2
    input   wire                 EN0,     // FO: 2
    input   wire [7:0]           A0,      // FO: 5
    input   wire [(WSIZE*8-1):0] Di0,     // FO: 2
    output  wire [(WSIZE*8-1):0] Do0
    );
    
    wire [1:0]             SEL0;
    wire [(WSIZE*8-1):0]    Do0_pre[1:0]; 
    assign SEL0[0] = EN0 && (~A0[7]);
    assign SEL0[1] = EN0 && ( A0[7]);
    
    generate
        genvar i;
        for (i=0; i< 2; i=i+1) begin : BANK128
            RAM128 RAM128 ( .CLK(CLK), .EN0(SEL0[i]), .WE0(WE0), .Di0(Di0), .Do0(Do0_pre[i]), .A0(A0[6:0]) );        
        end
    endgenerate
    
    assign Do0 = A0[7]? Do0_pre[1]:Do0_pre[0];
                                                                                                                                                          
endmodule
//`include "fsic_defines.v"

module RAM128 #(parameter USE_LATCH = 1,
                          WSIZE     = 4
)
(
    input   wire                 CLK,   
    input   wire [WSIZE-1:0]     WE0,   
    input   wire                 EN0,   
    input   wire [6:0]           A0,    
    input   wire [(WSIZE*8-1):0] Di0,   
    output  wire [(WSIZE*8-1):0] Do0
    );
    wire [(WSIZE*8-1):0]    Do0_pre[1:0]; 
    wire we;
    assign we = (WE0[3] && WE0[2] && WE0[1] && WE0[0]);
    ra1shd128x32m4h3v2 RAM128x32 ( .CLK(CLK), .CEN(~EN0), .WEN(~we), .OEN(1'b0), .D(Di0), .Q(Do0), .A(A0[6:0]) );

  
endmodule
//===========================================================
// Modified by Vic Chen
// Oct 5, 2024
//===========================================================

/* Copyright (C) 1991-2020 Free Software Foundation, Inc.
   This file is part of the GNU C Library.

   The GNU C Library is free software; you can redistribute it and/or
   modify it under the terms of the GNU Lesser General Public
   License as published by the Free Software Foundation; either
   version 2.1 of the License, or (at your option) any later version.

   The GNU C Library is distributed in the hope that it will be useful,
   but WITHOUT ANY WARRANTY; without even the implied warranty of
   MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
   Lesser General Public License for more details.

   You should have received a copy of the GNU Lesser General Public
   License along with the GNU C Library; if not, see
   <https://www.gnu.org/licenses/>.  */

/* This header is separate from features.h so that the compiler can
   include it implicitly at the start of every compilation.  It must
   not itself include <features.h> or any other header that includes
   <features.h> because the implicit include comes before any feature
   test macros that may be defined in a source file before it first
   explicitly includes a system header.  GCC knows the name of this
   header in order to preinclude it.  */

/* glibc's intent is to support the IEC 559 math functionality, real
   and complex.  If the GCC (4.9 and later) predefined macros
   specifying compiler intent are available, use them to determine
   whether the overall intent is to support these features; otherwise,
   presume an older compiler has intent to support these features and
   define these macros by default.  */
/* wchar_t uses Unicode 10.0.0.  Version 10.0 of the Unicode Standard is
   synchronized with ISO/IEC 10646:2017, fifth edition, plus
   the following additions from Amendment 1 to the fifth edition:
   - 56 emoji characters
   - 285 hentaigana
   - 3 additional Zanabazar Square characters */
 

// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/*--------------------------------------------------------------*/
/* caravel, a project harness for the Google/SkyWater sky130	*/
/* fabrication process and open source PDK			*/
/*                                                          	*/
/* Copyright 2020 efabless, Inc.                            	*/
/* Written by Tim Edwards, December 2019                    	*/
/* and Mohamed Shalan, August 2020			    	*/
/* This file is open source hardware released under the     	*/
/* Apache 2.0 license.  See file LICENSE.                   	*/
/*								*/
/* Updated 10/15/2021:  Revised using the housekeeping module	*/
/* from housekeeping.v (refactoring a number of functions from	*/
/* the management SoC).						*/
/*                                                          	*/
/*--------------------------------------------------------------*/
module caravel_top (
    inout [`MPRJ_IO_PADS-1:0]  mprj_io,

    //Willy debug - e
    input clock, // CMOS core clock input, not a crystal
    input resetb, // Reset input (sense inverted)

    // Note that only two flash data pins are dedicated to the
    // management SoC wrapper.  The management SoC exports the
    // quad SPI mode status to make use of the top two mprj_io
    // pins for io2 and io3.

    output flash_csb,
    output flash_clk,
    output flash_io0,
    input  flash_io1, //Willy debug

    inout gpio // Used for external LDO control
);


    //------------------------------------------------------------
    // This value is uniquely defined for each user project.
    //------------------------------------------------------------
    parameter USER_PROJECT_ID = 32'h00000000;

    /*
     *--------------------------------------------------------------------
     *
     * These pins are overlaid on mprj_io space.  They have the function
     * below when the management processor is in reset, or in the default
     * configuration.  They are assigned to uses in the user space by the
     * configuration program running off of the SPI flash.  Note that even
     * when the user has taken control of these pins, they can be restored
     * to the original use by setting the resetb pin low.  The SPI pins and
     * UART pins can be connected directly to an FTDI chip as long as the
     * FTDI chip sets these lines to high impedence (input function) at
     * all times except when holding the chip in reset.
     *
     * JTAG       = mprj_io[0]		(inout)
     * SDO 	  = mprj_io[1]		(output)
     * SDI 	  = mprj_io[2]		(input)
     * CSB 	  = mprj_io[3]		(input)
     * SCK	  = mprj_io[4]		(input)
     * ser_rx     = mprj_io[5]		(input)
     * ser_tx     = mprj_io[6]		(output)
     * irq 	  = mprj_io[7]		(input)
     *
     * spi_sck    = mprj_io[32]		(output)
     * spi_csb    = mprj_io[33]		(output)
     * spi_sdi    = mprj_io[34]		(input)
     * spi_sdo    = mprj_io[35]		(output)
     * flash_io2  = mprj_io[36]		(inout) 
     * flash_io3  = mprj_io[37]		(inout) 
     *
     * These pins are reserved for any project that wants to incorporate
     * its own processor and flash controller.  While a user project can
     * technically use any available I/O pins for the purpose, these
     * four pins connect to a pass-through mode from the SPI slave (pins
     * 1-4 above) so that any SPI flash connected to these specific pins
     * can be accessed through the SPI slave even when the processor is in
     * reset.
     *
     * user_flash_csb = mprj_io[8]
     * user_flash_sck = mprj_io[9]
     * user_flash_io0 = mprj_io[10]
     * user_flash_io1 = mprj_io[11]
     *
     *--------------------------------------------------------------------
     */
    //Willy debug - s
    //wire [`MPRJ_IO_PADS-1:0] mprj_io;
    //Willy debug - e


    // One-bit GPIO dedicated to management SoC (outside of user control)
    wire gpio_out_core;
    wire gpio_in_core;
    wire gpio_mode0_core;
    wire gpio_mode1_core;
    wire gpio_outenb_core;
    wire gpio_inenb_core;

    // User Project Control (pad-facing)
    wire [`MPRJ_IO_PADS-1:0] mprj_io_inp_dis;
    wire [`MPRJ_IO_PADS-1:0] mprj_io_oeb;
    wire [`MPRJ_IO_PADS-1:0] mprj_io_ib_mode_sel;
    wire [`MPRJ_IO_PADS-1:0] mprj_io_vtrip_sel;
    wire [`MPRJ_IO_PADS-1:0] mprj_io_slow_sel;
    wire [`MPRJ_IO_PADS-1:0] mprj_io_holdover;
    wire [`MPRJ_IO_PADS-1:0] mprj_io_analog_en;
    wire [`MPRJ_IO_PADS-1:0] mprj_io_analog_sel;
    wire [`MPRJ_IO_PADS-1:0] mprj_io_analog_pol;
    wire [`MPRJ_IO_PADS*3-1:0] mprj_io_dm;
    wire [`MPRJ_IO_PADS-1:0] mprj_io_in;
    wire [`MPRJ_IO_PADS-1:0] mprj_io_out;
    wire [`MPRJ_IO_PADS-1:0] mprj_io_one;

    // User Project Control (user-facing)
    wire [`MPRJ_IO_PADS-1:0] user_io_oeb;
    wire [`MPRJ_IO_PADS-1:0] user_io_in;
    wire [`MPRJ_IO_PADS-1:0] user_io_out;
    wire [`MPRJ_IO_PADS-10:0] user_analog_io;

    /* Padframe control signals */
    wire [`MPRJ_IO_PADS_1-1:0] gpio_serial_link_1;
    wire [`MPRJ_IO_PADS_2-1:0] gpio_serial_link_2;
    wire mprj_io_loader_resetn;
    wire mprj_io_loader_clock;
    wire mprj_io_loader_strobe;
    wire mprj_io_loader_data_1; /* user1 side serial loader */
    wire mprj_io_loader_data_2; /* user2 side serial loader */

    // User Project Control management I/O
    // There are two types of GPIO connections:
    // (1) Full Bidirectional: Management connects to in, out, and oeb
    //     Uses:  JTAG and SDO
    // (2) Selectable bidirectional:  Management connects to in and out,
    //	   which are tied together.  oeb is grounded (oeb from the
    //	   configuration is used)

    // SDI 	 = mprj_io[2]		(input)
    // CSB 	 = mprj_io[3]		(input)
    // SCK	 = mprj_io[4]		(input)
    // ser_rx    = mprj_io[5]		(input)
    // ser_tx    = mprj_io[6]		(output)
    // irq 	 = mprj_io[7]		(input)

    wire [`MPRJ_IO_PADS-1:0] mgmt_io_in; /* two- and three-pin data in	*/
    wire [`MPRJ_IO_PADS-1:0] mgmt_io_out; /* two- and three-pin data out	*/
    wire [`MPRJ_IO_PADS-1:0] mgmt_io_oeb; /* output enable, used only by	*/
      /* the three-pin interfaces	*/
    wire [`MPRJ_PWR_PADS-1:0] pwr_ctrl_nc; /* no-connects */

    /* Buffers are placed between housekeeping and gpio_control_block		*/
    /* instances to mitigate timing issues on very long (> 1.5mm) wires.	*/
    wire [`MPRJ_IO_PADS-1:0] mgmt_io_in_hk; /* mgmt_io_in at housekeeping	*/
    wire [`MPRJ_IO_PADS-1:0] mgmt_io_out_hk; /* mgmt_io_out at housekeeping	*/
    wire [`MPRJ_IO_PADS-1:0] mgmt_io_oeb_hk; /* mgmt_io_oeb at housekeeping	*/

    wire clock_core;

    // Power-on-reset signal.  The reset pad generates the sense-inverted
    // reset at 3.3V.  The 1.8V signal and the inverted 1.8V signal are
    // derived.

    wire porb_h;
    wire porb_l;
    wire por_l;

    wire rstb_h;
    wire rstb_l;

    // Flash SPI communication (management SoC to housekeeping)
    wire flash_clk_core, flash_csb_core;
    wire flash_clk_oeb_core, flash_csb_oeb_core;
    wire flash_io0_oeb_core, flash_io1_oeb_core;
    wire flash_io2_oeb_core, flash_io3_oeb_core;
    wire flash_io0_ieb_core, flash_io1_ieb_core;
    wire flash_io2_ieb_core, flash_io3_ieb_core;
    wire flash_io0_do_core, flash_io1_do_core;
    wire flash_io2_do_core, flash_io3_do_core;
    wire flash_io0_di_core, flash_io1_di_core;
    wire flash_io2_di_core, flash_io3_di_core;

    // Flash SPI communication (
    wire flash_clk_frame;
    wire flash_csb_frame;
    wire flash_clk_oeb, flash_csb_oeb;
    wire flash_clk_ieb, flash_csb_ieb;
    wire flash_io0_oeb, flash_io1_oeb;
    wire flash_io0_ieb, flash_io1_ieb;
    wire flash_io0_do, flash_io1_do;
    wire flash_io0_di, flash_io1_di;

 // Flash buffered signals
    wire flash_clk_frame_buf;
    wire flash_csb_frame_buf;
    wire flash_clk_ieb_buf, flash_csb_ieb_buf;
    wire flash_io0_oeb_buf, flash_io1_oeb_buf;
    wire flash_io0_ieb_buf, flash_io1_ieb_buf;
    wire flash_io0_do_buf, flash_io1_do_buf;
    wire flash_io0_di_buf, flash_io1_di_buf;

   // Clock and reset buffered signals
   wire caravel_clk_buf;
   wire caravel_rstn_buf;
   wire clock_core_buf;

 // SoC pass through buffered signals
 wire mprj_io_loader_clock_buf;
 wire mprj_io_loader_strobe_buf;
 wire mprj_io_loader_resetn_buf;
 wire mprj_io_loader_data_2_buf;
 wire rstb_l_buf;
 wire por_l_buf;
 wire porb_h_buf;


    // SoC core
    wire caravel_clk;
    wire caravel_clk2;
    wire caravel_rstn;
    
//Willy debug - s
//assign mprj_o = mprj_io_out;
//assign mprj_en = mprj_io_oeb;
//assign mprj_io_in = mprj_i;

   //================ Start of Padframe ================//
   //================= IO Configure ====================//
   // Input:  OEN = 1, REN = 0 during reset operation
   //         OEN = 1, REN = 1 during normal operation
   //---------------------------------------------------//
   // Output: OEN = 1, REN = 1 during reset operation
   //         OEN = 0, REN = 1 during normal operation
   //===================================================//
   wire        REN;
   wire [37:0] mprj_oen;


    // Input Pad for MPRJ
    `define INPAD_MPRJ(n) \
        PDDWDGZ iopad_MPRJ``n(  \
            .C(mprj_io_in[n]),  \
            .PAD(mprj_io[n]),   \
            .REN(REN)           \
        );

    `define IOPAD_MPRJ(n)         \
        PDUW04DGZ iopad_MPRJ``n(  \
            .I(mprj_io_out[n]),   \
            .C(mprj_io_in[n]),    \
            .OEN(mprj_oen[n]),    \
            .PAD(mprj_io[n]),     \
            .REN(REN)             \
        );

    PDDWDGZ iopad_CLK(
        .PAD(clock), 
        .C(clock_core),
        .REN(REN)
    );
    PDISDGZ iopad_RST(
        .C(resetb_core),
        .PAD(resetb)
    );

    wire fcsb_oen, fclk_oen, fio0_oen, fio1_oen;
    assign fclk_oen = 1'b0 | (~resetb_core);
    assign fcsb_oen = 1'b0 | (~resetb_core);
    assign fio0_oen = 1'b0 | (~resetb_core);
    assign fio1_oen = 1'b1 | (~resetb_core);
    assign gpio_oen = 1'b1 | (~resetb_core);

    PDUW04DGZ iopad_FCSB(
        .PAD(flash_csb), 
        .I(flash_csb_frame_buf), 
        .C(), 
        .OEN(fcsb_oen), 
        .REN(REN)
    );
    PDUW04DGZ iopad_FCLK(
        .PAD(flash_clk), 
        .I(flash_clk_frame_buf), 
        .C(), 
        .OEN(fclk_oen), 
        .REN(REN)
    );
    PDUW04DGZ iopad_FIO0(
        .PAD(flash_io0), 
        .I(flash_io0_do_buf), 
    	  .C(flash_io0_di), 
        .OEN(fio0_oen), 
        .REN(REN)
    );
    PDUW04DGZ iopad_FIO1(
        .PAD(flash_io1), 
        .I(flash_io1_do_buf), 
    	  .C(flash_io1_di), 
        .OEN(fio1_oen), 
        .REN(REN)
    );
    // Management GPIO pad
    PDUW04DGZ iopad_GPIO(
        .PAD(gpio), 
        .I(gpio_out_core), 
        .C(gpio_in_core), 
        .OEN(gpio_oen), 
        .REN(REN)
    );
    // Instance 38 MPRJ Pads
    `IOPAD_MPRJ(0)   // JTAG
    `IOPAD_MPRJ(1)   // SDO
    `IOPAD_MPRJ(2)   // SDI
    `IOPAD_MPRJ(3)   // CSB
    `IOPAD_MPRJ(4)   // SCK
    `IOPAD_MPRJ(5)   // ser_rx
    `IOPAD_MPRJ(6)   // ser_tx
    `INPAD_MPRJ(7)   // irq
    
    `INPAD_MPRJ(8)   // RXD[0]
    `INPAD_MPRJ(9)   // RXD[1]
    `INPAD_MPRJ(10)  // RXD[2]
    `INPAD_MPRJ(11)  // RXD[3]
    `INPAD_MPRJ(12)  // RXD[4]
    `INPAD_MPRJ(13)  // RXD[5]
    `INPAD_MPRJ(14)  // RXD[6]
    `INPAD_MPRJ(15)  // RXD[7]
    `INPAD_MPRJ(16)  // RXD[8]
    `INPAD_MPRJ(17)  // RXD[9]
    `INPAD_MPRJ(18)  // RXD[10]
    `INPAD_MPRJ(19)  // RXD[11]
    `INPAD_MPRJ(20)  // RXD[12]
    `INPAD_MPRJ(21)  // RXCLK
    
    `IOPAD_MPRJ(22)  // TXD[0]
    `IOPAD_MPRJ(23)  // TXD[1]
    `IOPAD_MPRJ(24)  // TXD[2]
    `IOPAD_MPRJ(25)  // TXD[3]
    `IOPAD_MPRJ(26)  // TXD[4]
    `IOPAD_MPRJ(27)  // TXD[5]
    `IOPAD_MPRJ(28)  // TXD[6]
    `IOPAD_MPRJ(29)  // TXD[7]
    `IOPAD_MPRJ(30)  // TXD[8]
    `IOPAD_MPRJ(31)  // TXD[9]
    `IOPAD_MPRJ(32)  // TXD[10]
    `IOPAD_MPRJ(33)  // TXD[11]
    `IOPAD_MPRJ(34)  // TXD[12]
    `IOPAD_MPRJ(35)  // TXCLK
    
    `INPAD_MPRJ(36)  // IOCLK
    `IOPAD_MPRJ(37)  // NOT USE


//Willy debug - e
    
    
 // FPGA - Remove module buff_flash_clkrst - bypass the buffer
 //  .A({in_n, in_s}), 
 //	.X({out_s, out_n})); 
 assign {caravel_clk_buf,
  caravel_rstn_buf,
  flash_clk_frame_buf,
  flash_csb_frame_buf,
  flash_clk_oeb_buf,
  flash_csb_oeb_buf,
  flash_io0_oeb_buf,
  flash_io1_oeb_buf,
  flash_io0_ieb_buf,
  flash_io1_ieb_buf,
  flash_io0_do_buf,
  flash_io1_do_buf } =
  {
  caravel_clk,
  caravel_rstn,
  flash_clk_frame,
  flash_csb_frame,
  flash_clk_oeb,
  flash_csb_oeb,
  flash_io0_oeb,
  flash_io1_oeb,
  flash_io0_ieb,
  flash_io1_ieb,
  flash_io0_do,
  flash_io1_do };
 assign
 {
  clock_core_buf,
  flash_io1_di_buf,
  flash_io0_di_buf } =
 {
  clock_core,
  flash_io1_di,
  flash_io0_di };
// end of module buff_flash_clkrst 




  /* NOTE: The first 7 GPIO are unbuffered, and all
		 * OEB lines except the last three are unbuffered
		 * (most of these end up being no-connects from
		 * housekeeping).
		 */
  assign mgmt_io_in_hk[6:0] = mgmt_io_in[6:0];
  assign mgmt_io_out[6:0] = mgmt_io_out_hk[6:0];
  assign mgmt_io_oeb[34:0] = mgmt_io_oeb_hk[34:0];
// FPGA Remove module gpio_signal_buffering
  assign mgmt_io_in_hk[37:7] = mgmt_io_in[37:7];
         assign mgmt_io_out[37:7] = mgmt_io_out_hk[37:7];
  assign mgmt_io_oeb[37:35] = mgmt_io_oeb_hk[37:35];


/*
 chip_io padframe(
// FPGA: Remove vdd, vss, ports
 // Core Side Pins
 .gpio(gpio),
 .mprj_io(mprj_io),
 .clock(clock),
 .resetb(resetb),
 .flash_csb(flash_csb),
 .flash_clk(flash_clk),
 .flash_io0(flash_io0),
 .flash_io1(flash_io1),
 // SoC Core Interface
 .porb_h(porb_h),
 .por(por_l_buf),
 .resetb_core_h(rstb_h),
 .clock_core(clock_core),
 .gpio_out_core(gpio_out_core),
 .gpio_in_core(gpio_in_core),
 .gpio_mode0_core(gpio_mode0_core),
 .gpio_mode1_core(gpio_mode1_core),
 .gpio_outenb_core(gpio_outenb_core),
 .gpio_inenb_core(gpio_inenb_core),
 .flash_csb_core(flash_csb_frame_buf),
 .flash_clk_core(flash_clk_frame_buf),
 .flash_csb_oeb_core(flash_csb_oeb_buf),
 .flash_clk_oeb_core(flash_clk_oeb_buf),
 .flash_io0_oeb_core(flash_io0_oeb_buf),
 .flash_io1_oeb_core(flash_io1_oeb_buf),
 .flash_io0_ieb_core(flash_io0_ieb_buf),
 .flash_io1_ieb_core(flash_io1_ieb_buf),
 .flash_io0_do_core(flash_io0_do_buf),
 .flash_io1_do_core(flash_io1_do_buf),
 .flash_io0_di_core(flash_io0_di),
 .flash_io1_di_core(flash_io1_di),
 .mprj_io_one(mprj_io_one),
//Willy debug .mprj_io_in(mprj_io_in),
 .mprj_io_out(mprj_io_out),
 .mprj_io_oeb(mprj_io_oeb),
 .mprj_io_inp_dis(mprj_io_inp_dis),
 .mprj_io_ib_mode_sel(mprj_io_ib_mode_sel),
 .mprj_io_vtrip_sel(mprj_io_vtrip_sel),
 .mprj_io_slow_sel(mprj_io_slow_sel),
 .mprj_io_holdover(mprj_io_holdover),
 .mprj_io_analog_en(mprj_io_analog_en),
 .mprj_io_analog_sel(mprj_io_analog_sel),
 .mprj_io_analog_pol(mprj_io_analog_pol),
 .mprj_io_dm(mprj_io_dm),
 .mprj_analog_io(user_analog_io)
    );
*/

    // Logic analyzer signals
    wire [127:0] la_data_in_user; // From CPU to MPRJ
    wire [127:0] la_data_in_mprj; // From MPRJ to CPU
    wire [127:0] la_data_out_mprj; // From CPU to MPRJ
    wire [127:0] la_data_out_user; // From MPRJ to CPU
    wire [127:0] la_oenb_user; // From CPU to MPRJ
    wire [127:0] la_oenb_mprj; // From CPU to MPRJ
    wire [127:0] la_iena_mprj; // From CPU only

    wire [2:0] user_irq; // From MRPJ to CPU
    wire [2:0] user_irq_core;
    wire [2:0] user_irq_ena;
    wire [2:0] irq_spi; // From SPI and external pins

    // Exported Wishbone Bus (processor facing)
    wire mprj_iena_wb;
    wire mprj_cyc_o_core;
    wire mprj_stb_o_core;
    wire mprj_we_o_core;
    wire [3:0] mprj_sel_o_core;
    wire [31:0] mprj_adr_o_core;
    wire [31:0] mprj_dat_o_core;
    wire mprj_ack_i_core;
    wire [31:0] mprj_dat_i_core;

    wire [31:0] hk_dat_i;
    wire hk_ack_i;
    wire hk_stb_o;
    wire hk_cyc_o;

    // Exported Wishbone Bus (user area facing)
    wire mprj_cyc_o_user;
    wire mprj_stb_o_user;
    wire mprj_we_o_user;
    wire [3:0] mprj_sel_o_user;
    wire [31:0] mprj_adr_o_user;
    wire [31:0] mprj_dat_o_user;
    wire [31:0] mprj_dat_i_user;
    wire mprj_ack_i_user;

    // Mask revision
    wire [31:0] mask_rev;

    wire mprj_clock;
    wire mprj_clock2;
    wire mprj_reset;

    // Power monitoring 


    // Management processor (wrapper).  Any management core
    // implementation must match this pinout.

    // Pass thru clock and reset
    wire clk_passthru;
    wire resetn_passthru;

 // NC passthru signal porb_h 
 //wire porb_h_in_nc;
 //wire porb_h_out_nc;

    mgmt_core_wrapper soc (

	    // SoC pass through buffered signals
	    .serial_clock_in(mprj_io_loader_clock),
	    .serial_clock_out(mprj_io_loader_clock_buf),
	    .serial_load_in(mprj_io_loader_strobe),
	    .serial_load_out(mprj_io_loader_strobe_buf),
	    .serial_resetn_in(mprj_io_loader_resetn),
	    .serial_resetn_out(mprj_io_loader_resetn_buf),
	    .serial_data_2_in(mprj_io_loader_data_2),
	    .serial_data_2_out(mprj_io_loader_data_2_buf),
	    .rstb_l_in(rstb_l),
	    .rstb_l_out(rstb_l_buf),

		 // [Vic]: POR is useless here
	    //.porb_h_in(porb_h_in_nc),
	    //.porb_h_out(porb_h_out_nc),
	    //.por_l_in(por_l),
	    //.por_l_out(por_l_buf),
    
	    // Clock and reset
	    .core_clk(caravel_clk_buf),
	    .core_rstn(caravel_rstn_buf),
    
        // Pass thru Clock and reset
	    .clk_in(caravel_clk_buf),
	    .resetn_in(caravel_rstn_buf),
	    .clk_out(clk_passthru),
	    .resetn_out(resetn_passthru),
    
	    // GPIO (1 pin)
	    .gpio_out_pad(gpio_out_core),
	    .gpio_in_pad(gpio_in_core),
	    .gpio_mode0_pad(gpio_mode0_core),
	    .gpio_mode1_pad(gpio_mode1_core),
	    .gpio_outenb_pad(gpio_outenb_core),
	    .gpio_inenb_pad(gpio_inenb_core),
    
	    // Primary SPI flash controller
	    .flash_csb(flash_csb_core),
	    .flash_clk(flash_clk_core),
	    .flash_io0_oeb(flash_io0_oeb_core),
	    .flash_io0_di(flash_io0_di_core),
	    .flash_io0_do(flash_io0_do_core),
	    .flash_io1_oeb(flash_io1_oeb_core),
	    .flash_io1_di(flash_io1_di_core),
	    .flash_io1_do(flash_io1_do_core),
	    .flash_io2_oeb(flash_io2_oeb_core),
	    .flash_io2_di(flash_io2_di_core),
	    .flash_io2_do(flash_io2_do_core),
	    .flash_io3_oeb(flash_io3_oeb_core),
	    .flash_io3_di(flash_io3_di_core),
	    .flash_io3_do(flash_io3_do_core),
    
	    // Exported Wishbone Bus
	    .mprj_wb_iena(mprj_iena_wb),
	    .mprj_cyc_o(mprj_cyc_o_core),
	    .mprj_stb_o(mprj_stb_o_core),
	    .mprj_we_o(mprj_we_o_core),
	    .mprj_sel_o(mprj_sel_o_core),
	    .mprj_adr_o(mprj_adr_o_core),
	    .mprj_dat_o(mprj_dat_o_core),
	    .mprj_ack_i(mprj_ack_i_core),
	    .mprj_dat_i(mprj_dat_i_core),
    
	    .hk_stb_o(hk_stb_o),
	    .hk_cyc_o(hk_cyc_o),
	    .hk_dat_i(hk_dat_i),
	    .hk_ack_i(hk_ack_i),
    
	    // IRQ
	    .irq({irq_spi, user_irq}),
	    .user_irq_ena(user_irq_ena),
    
	    // Module status (these may or may not be implemented)
	    .qspi_enabled(qspi_enabled),
	    .uart_enabled(uart_enabled),
	    .spi_enabled(spi_enabled),
	    .debug_mode(debug_mode),
    
	    // Module I/O (these may or may not be implemented)
	    // UART
	    .ser_tx(ser_tx),
	    .ser_rx(ser_rx),
	    // SPI master
	    .spi_sdi(spi_sdi),
	    .spi_csb(spi_csb),
	    .spi_sck(spi_sck),
	    .spi_sdo(spi_sdo),
	    .spi_sdoenb(spi_sdoenb),
	    // Debug
	    .debug_in(debug_in),
	    .debug_out(debug_out),
	    .debug_oeb(debug_oeb),
	    // Logic analyzer
	    .la_input(la_data_in_mprj),
	    .la_output(la_data_out_mprj),
	    .la_oenb(la_oenb_mprj),
	    .la_iena(la_iena_mprj),
    
    	// Trap status
    	.trap(trap)
    );

    /* Clock and reset to user space are passed through a tristate	*/
    /* buffer like the above, but since they are intended to be		*/
    /* always active, connect the enable to the logic-1 output from	*/
    /* the vccd1 domain.						*/
// FPGA : Remove mgmt_protect module, passthrough


 assign la_data_in_mprj = la_data_out_user;
 assign la_data_in_user = la_data_out_mprj;
 assign la_oenb_user = la_oenb_mprj;

   assign mprj_clock = clk_passthru;
   assign mprj_clock2 = caravel_clk2;
   assign mprj_reset = ~resetn_passthru; // Note: it is inversted - mprj_reset is active high
   assign mprj_cyc_o_user = mprj_cyc_o_core;
   assign mprj_stb_o_user = mprj_stb_o_core;
   assign mprj_we_o_user = mprj_we_o_core;
   assign mprj_sel_o_user = mprj_sel_o_core;
   assign mprj_adr_o_user = mprj_adr_o_core;
   assign mprj_dat_o_user = mprj_dat_o_core;
   assign mprj_dat_i_core = mprj_dat_i_user;
   assign mprj_ack_i_core = mprj_ack_i_user;
   assign user_irq = user_irq_core;

   assign user1_vcc_powergood = 1'b1;
   assign user2_vcc_powergood = 1'b1;
   assign user1_vdd_powergood = 1'b1;
   assign user2_vdd_powergood = 1'b1;

    /*--------------------------------------------------*/
    /* Wrapper module around the user project 		*/
    /*--------------------------------------------------*/
   wire        uspj_cyc; // CYC
   wire        uspj_ack;
   wire [31:0] uspj_dat;

   user_project_wrapper mprj (

      .wb_clk_i(mprj_clock),
      .wb_rst_i(mprj_reset),

      // Management SoC Wishbone bus (exported)
      .wbs_cyc_i(uspj_cyc),
      .wbs_stb_i(mprj_stb_o_user),
      .wbs_we_i(mprj_we_o_user),
      .wbs_sel_i(mprj_sel_o_user),
      .wbs_adr_i(mprj_adr_o_user),
      .wbs_dat_i(mprj_dat_o_user),
      .wbs_ack_o(uspj_ack),
      .wbs_dat_o(uspj_dat),

      // GPIO pad 3-pin interface (plus analog)
      .io_in (user_io_in),
      .io_out(user_io_out),
      .io_oeb(user_io_oeb),
      //.analog_io(user_analog_io),

      // Logic analyzer
      .la_data_in(la_data_in_user),
      .la_data_out(la_data_out_user),
      .la_oenb(la_oenb_user),

      // Independent clock
      .user_clock2(mprj_clock2),

      // IRQ
      .user_irq(user_irq_core)
   );

   //======================================================//
   // [Vic]: PAD IOs should also be flexible
   //======================================================//
   wire        wb_mux;
   wire        io_cnfg_cyc;
   wire        io_cnfg_ack;
   wire [31:0] io_cnfg_dat;

   pads_config PAD_IO_CNFG (
  	   .clk(clock_core),
	   .resetb(resetb_core),
	   .wb_clk_i(mprj_clock),
	   .wb_rst_i(mprj_reset),
	   .wbs_cyc_i(io_cnfg_cyc),
	   .wbs_stb_i(mprj_stb_o_user),
	   .wbs_we_i(mprj_we_o_user),
	   .wbs_sel_i(mprj_sel_o_user),
	   .wbs_adr_i(mprj_adr_o_user),
	   .wbs_dat_i(mprj_dat_o_user),
	   .wbs_ack_o(io_cnfg_ack),
	   .wbs_dat_o(io_cnfg_dat),
	   .re_n(REN),
	   .oe_n(mprj_oen)
   );
   // IO configuration area: 3000_6000 ~ 3000_6025
   assign wb_mux = (mprj_adr_o_user[31:12] == 20'h3000_6)? 1'b1 : 1'b0;
   assign uspj_cyc    = (wb_mux)? 0 : mprj_cyc_o_user;
   assign io_cnfg_cyc = (wb_mux)? mprj_cyc_o_user : 0;
   assign mprj_ack_i_user = (wb_mux)? io_cnfg_ack : uspj_ack;
   assign mprj_dat_i_user = (wb_mux)? io_cnfg_dat : uspj_dat;
   //======================================================//


    wire [`MPRJ_IO_PADS_1-1:0] gpio_serial_link_1_shifted;
    wire [`MPRJ_IO_PADS_2-1:0] gpio_serial_link_2_shifted;

    assign gpio_serial_link_1_shifted = {gpio_serial_link_1[`MPRJ_IO_PADS_1-2:0],
      mprj_io_loader_data_1};
    // Note that serial_link_2 is backwards compared to serial_link_1, so it
    // shifts in the other direction.
    assign gpio_serial_link_2_shifted = {mprj_io_loader_data_2_buf,
      gpio_serial_link_2[`MPRJ_IO_PADS_2-1:1]};

    // Propagating clock and reset to mitigate timing and fanout issues
    wire [`MPRJ_IO_PADS_1-1:0] gpio_clock_1;
    wire [`MPRJ_IO_PADS_2-1:0] gpio_clock_2;
    wire [`MPRJ_IO_PADS_1-1:0] gpio_resetn_1;
    wire [`MPRJ_IO_PADS_2-1:0] gpio_resetn_2;
    wire [`MPRJ_IO_PADS_1-1:0] gpio_load_1;
    wire [`MPRJ_IO_PADS_2-1:0] gpio_load_2;
    wire [`MPRJ_IO_PADS_1-1:0] gpio_clock_1_shifted;
    wire [`MPRJ_IO_PADS_2-1:0] gpio_clock_2_shifted;
    wire [`MPRJ_IO_PADS_1-1:0] gpio_resetn_1_shifted;
    wire [`MPRJ_IO_PADS_2-1:0] gpio_resetn_2_shifted;
    wire [`MPRJ_IO_PADS_1-1:0] gpio_load_1_shifted;
    wire [`MPRJ_IO_PADS_2-1:0] gpio_load_2_shifted;

    assign gpio_clock_1_shifted = {gpio_clock_1[`MPRJ_IO_PADS_1-2:0],
      mprj_io_loader_clock};
    assign gpio_clock_2_shifted = {mprj_io_loader_clock_buf,
     gpio_clock_2[`MPRJ_IO_PADS_2-1:1]};
    assign gpio_resetn_1_shifted = {gpio_resetn_1[`MPRJ_IO_PADS_1-2:0],
      mprj_io_loader_resetn};
    assign gpio_resetn_2_shifted = {mprj_io_loader_resetn_buf,
     gpio_resetn_2[`MPRJ_IO_PADS_2-1:1]};
    assign gpio_load_1_shifted = {gpio_load_1[`MPRJ_IO_PADS_1-2:0],
      mprj_io_loader_strobe};
    assign gpio_load_2_shifted = {mprj_io_loader_strobe_buf,
     gpio_load_2[`MPRJ_IO_PADS_2-1:1]};

    wire [2:0] spi_pll_sel;
    wire [2:0] spi_pll90_sel;
    wire [4:0] spi_pll_div;
    wire [25:0] spi_pll_trim;
    wire  ext_reset;
// FPGA Remove module caravel_clocking: clock/reset directly from IO pad
    assign caravel_clk = clock_core_buf;
    assign caravel_clk2 = clock_core_buf;
    assign caravel_rstn = rstb_l_buf // original design : sync rstb_l_buf 3T 
                          & ~ext_reset;

   // DCO/Digital Locked Loop
   // FPGA: Remove digital_pll

   // Housekeeping interface

   housekeeping housekeeping (
         .wb_clk_i(caravel_clk),
         .wb_rstn_i(caravel_rstn),
 
         .wb_adr_i(mprj_adr_o_core),
         .wb_dat_i(mprj_dat_o_core),
         .wb_sel_i(mprj_sel_o_core),
         .wb_we_i(mprj_we_o_core),
         .wb_cyc_i(hk_cyc_o),
         .wb_stb_i(hk_stb_o),
         .wb_ack_o(hk_ack_i),
         .wb_dat_o(hk_dat_i),
 
         .porb(porb_l),
 
         .pll_ena(spi_pll_ena),
         .pll_dco_ena(spi_pll_dco_ena),
         .pll_div(spi_pll_div),
         .pll_sel(spi_pll_sel),
         .pll90_sel(spi_pll90_sel),
         .pll_trim(spi_pll_trim),
         .pll_bypass(ext_clk_sel),
 
  .qspi_enabled(qspi_enabled),
  .uart_enabled(uart_enabled),
  .spi_enabled(spi_enabled),
  .debug_mode(debug_mode),
 
  .ser_tx(ser_tx),
  .ser_rx(ser_rx),
 
  .spi_sdi(spi_sdi),
  .spi_csb(spi_csb),
  .spi_sck(spi_sck),
  .spi_sdo(spi_sdo),
  .spi_sdoenb(spi_sdoenb),
 
  .debug_in(debug_in),
  .debug_out(debug_out),
  .debug_oeb(debug_oeb),
 
         .irq(irq_spi),
         .reset(ext_reset),
 
         .serial_clock(mprj_io_loader_clock),
         .serial_load(mprj_io_loader_strobe),
         .serial_resetn(mprj_io_loader_resetn),
         .serial_data_1(mprj_io_loader_data_1),
         .serial_data_2(mprj_io_loader_data_2),
 
  .mgmt_gpio_in(mgmt_io_in_hk),
  .mgmt_gpio_out(mgmt_io_out_hk),
  .mgmt_gpio_oeb(mgmt_io_oeb_hk),
 
  .pwr_ctrl_out(pwr_ctrl_nc), /* Not used in this version */
 
         .trap(trap),
 
  .user_clock(caravel_clk2),
 
         .mask_rev_in(mask_rev),
 
  .spimemio_flash_csb(flash_csb_core),
  .spimemio_flash_clk(flash_clk_core),
  .spimemio_flash_io0_oeb(flash_io0_oeb_core),
  .spimemio_flash_io1_oeb(flash_io1_oeb_core),
  .spimemio_flash_io2_oeb(flash_io2_oeb_core),
  .spimemio_flash_io3_oeb(flash_io3_oeb_core),
  .spimemio_flash_io0_do(flash_io0_do_core),
  .spimemio_flash_io1_do(flash_io1_do_core),
  .spimemio_flash_io2_do(flash_io2_do_core),
  .spimemio_flash_io3_do(flash_io3_do_core),
  .spimemio_flash_io0_di(flash_io0_di_core),
  .spimemio_flash_io1_di(flash_io1_di_core),
  .spimemio_flash_io2_di(flash_io2_di_core),
  .spimemio_flash_io3_di(flash_io3_di_core),
 
  .pad_flash_csb(flash_csb_frame),
  .pad_flash_csb_oeb(flash_csb_oeb),
  .pad_flash_clk(flash_clk_frame),
  .pad_flash_clk_oeb(flash_clk_oeb),
  .pad_flash_io0_oeb(flash_io0_oeb),
  .pad_flash_io1_oeb(flash_io1_oeb),
  .pad_flash_io0_ieb(flash_io0_ieb),
  .pad_flash_io1_ieb(flash_io1_ieb),
  .pad_flash_io0_do(flash_io0_do),
  .pad_flash_io1_do(flash_io1_do),
  .pad_flash_io0_di(flash_io0_di_buf),
  .pad_flash_io1_di(flash_io1_di_buf),


   .usr1_vcc_pwrgood(user1_vcc_powergood),
   .usr2_vcc_pwrgood(user2_vcc_powergood),
   .usr1_vdd_pwrgood(user1_vdd_powergood),
   .usr2_vdd_pwrgood(user2_vdd_powergood)
    );

    // [Vic]: Remove GPIO configuration logics
    assign mprj_io_out = user_io_out;
    assign user_io_in  = mprj_io_in;
    assign mgmt_io_in  = mprj_io_in;

// FPGA: Remove module user_id_programming
    assign mask_rev = USER_PROJECT_ID;


   // Power-on-reset circuit
   // FPGA: Remove module "simple_por", "xres_buf"
   // Hack por equal to resetb
   assign porb_h = resetb_core;
   assign porb_l = resetb_core;
   assign por_l = ~porb_l;
// rstb_l is a level-shift version of rstb_h
    assign rstb_l = resetb_core;
// FPGA: remove module spare_logic_block


endmodule
// `default_nettype wire
//===========================================================
// Modified by Vic Chen
// July 26, 2024
//===========================================================

// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

//-----------------------------------------------------------
// Housekeeping interface for Caravel
//-----------------------------------------------------------
// Written by Tim Edwards
// efabless, inc. September 27, 2020
//-----------------------------------------------------------

//-----------------------------------------------------------
// This is a standalone slave SPI for the caravel chip that is
// intended to be independent of the picosoc and independent
// of all IP blocks except the power-on-reset.  This SPI has
// register outputs controlling the functions that critically
// affect operation of the picosoc and so cannot be accessed
// from the picosoc itself.  This includes the PLL enables,
// mode, and trim.  It also has a general reset for the picosoc,
// an IRQ input, a bypass for the entire crystal oscillator
// and PLL chain, the manufacturer and product IDs and product
// revision number.
//
// Updated and revised, 10/13/2021:
// This module now comprises what was previously split into
// the housekeeping SPI, the mprj_ctrl block (control over
// the GPIO), and sysctrl (redirection of certain internal
// signals to the GPIO);  and additionally manages the SPI
// flash signals and pass-through mode.  Essentially all
// aspects of the system related to the use and configuration
// of the GPIO has been shifted to this module.  This allows
// GPIO to be configured from either the management SoC
// through the wishbone interface, or externally through the
// SPI interface.  It allows essentially any processor to
// take the place of the PicoRV32 as long as that processor
// can access memory-mapped space via the wishbone bus.
//-----------------------------------------------------------

//------------------------------------------------------------
// Caravel defined registers (by SPI address):
// See:  doc/memory_map.txt
//------------------------------------------------------------

module housekeeping #(
    parameter GPIO_BASE_ADR = 32'h2600_0000,
    parameter SPI_BASE_ADR = 32'h2610_0000,
    parameter SYS_BASE_ADR = 32'h2620_0000,
    parameter IO_CTRL_BITS = 13
) (
    inout wire VPWR,
    inout wire VGND,

    // Wishbone interface to management SoC
    input wire wb_clk_i,
    input wire wb_rstn_i,
    input wire [31:0] wb_adr_i,
    input wire [31:0] wb_dat_i,
    input wire [3:0] wb_sel_i,
    input wire wb_we_i,
    input wire wb_cyc_i,
    input wire wb_stb_i,
    output reg wb_ack_o,
    output reg [31:0] wb_dat_o,

    // Primary reset
    input wire porb,

	/////////////////////////////
	//// [Vic]: PLL is unsed ////
	// Clocking control parameters
    output reg pll_ena,
    output reg pll_dco_ena,
    output reg [4:0] pll_div,
    output reg [2:0] pll_sel,
    output reg [2:0] pll90_sel,
    output reg [25:0] pll_trim,
    output reg pll_bypass,
	/////////////////////////////

    // Module enable status from SoC
    input wire qspi_enabled,
    input wire uart_enabled,
    input wire spi_enabled,
    input wire debug_mode,
    
    // UART interface to/from SoC
    input wire ser_tx,
    output wire ser_rx,

    // SPI master interface to/from SoC
    output wire spi_sdi,
    input wire spi_csb,
    input wire spi_sck,
    input wire spi_sdo,
    input wire spi_sdoenb,

    // External (originating from SPI and pad) IRQ and reset
    output wire [2:0] irq,
    output wire reset,

    // GPIO serial loader programming interface
    output wire serial_clock,
    output wire serial_load,
    output wire serial_resetn,
    output wire serial_data_1,
    output wire serial_data_2,

    // GPIO data management (to padframe)---three-pin interface
    input wire [`MPRJ_IO_PADS-1:0] mgmt_gpio_in,
    output wire [`MPRJ_IO_PADS-1:0] mgmt_gpio_out,
    output wire [`MPRJ_IO_PADS-1:0] mgmt_gpio_oeb,

    // Power control output (reserved for future use with LDOs)
    output reg [`MPRJ_PWR_PADS-1:0] pwr_ctrl_out,

    // CPU trap state status (for system monitoring)
    input wire trap,

    // User clock (for system monitoring)
    input wire user_clock,

    // Mask revision/User project ID
    input wire [31:0] mask_rev_in,

    // SPI flash management (management SoC side)
    input wire spimemio_flash_csb,
    input wire spimemio_flash_clk,
    input wire spimemio_flash_io0_oeb,
    input wire spimemio_flash_io1_oeb,
    input wire spimemio_flash_io2_oeb,
    input wire spimemio_flash_io3_oeb,
    input wire spimemio_flash_io0_do,
    input wire spimemio_flash_io1_do,
    input wire spimemio_flash_io2_do,
    input wire spimemio_flash_io3_do,
    output wire spimemio_flash_io0_di,
    output wire spimemio_flash_io1_di,
    output wire spimemio_flash_io2_di,
    output wire spimemio_flash_io3_di,

    // Debug interface (routes to first GPIO) from management SoC
    output wire debug_in,
    input wire debug_out,
    input wire debug_oeb,

    // SPI flash management (padframe side)
    // (io2 and io3 are part of GPIO array, not dedicated pads)
    output wire pad_flash_csb,
    output wire pad_flash_csb_oeb,
    output wire pad_flash_clk,
    output wire pad_flash_clk_oeb,
    output wire pad_flash_io0_oeb,
    output wire pad_flash_io1_oeb,
    output wire pad_flash_io0_ieb,
    output wire pad_flash_io1_ieb,
    output wire pad_flash_io0_do,
    output wire pad_flash_io1_do,
    input wire pad_flash_io0_di,
    input wire pad_flash_io1_di,
    

    // System signal monitoring
    input wire usr1_vcc_pwrgood,
    input wire usr2_vcc_pwrgood,
    input wire usr1_vdd_pwrgood,
    input wire usr2_vdd_pwrgood
);

    localparam OEB = 1;		// Offset of output enable (bar) in shift register
    localparam INP_DIS = 3;	// Offset of input disable in shift register

    reg reset_reg;
    reg irq_spi;
    reg serial_bb_clock;
    reg serial_bb_load;
    reg serial_bb_resetn;
    reg serial_bb_data_1;
    reg serial_bb_data_2;
    reg serial_bb_enable;
    reg serial_xfer;
    reg hkspi_disable;

    reg clk1_output_dest;
    reg clk2_output_dest;
    reg trap_output_dest;
    reg irq_1_inputsrc;
    reg irq_2_inputsrc;

    reg [IO_CTRL_BITS-1:0] gpio_configure [`MPRJ_IO_PADS-1:0];
    reg [`MPRJ_IO_PADS-1:0] mgmt_gpio_data;

    /* mgmt_gpio_data_buf holds the lower bits during a back-door
     * write to GPIO data so that all 32 bits can update at once.
     */
    reg [23:0] mgmt_gpio_data_buf;


    wire [7:0] odata;
    wire [7:0] idata;
    wire [7:0] iaddr;

    wire rdstb;
    wire wrstb;
    wire pass_thru_mgmt;		// Mode detected by housekeeping_spi
    wire pass_thru_mgmt_delay;
    wire pass_thru_user;		// Mode detected by housekeeping_spi
    wire pass_thru_user_delay;
    wire pass_thru_mgmt_reset;
    wire pass_thru_user_reset;
    wire sdo;
    wire sdo_enb;

    wire [7:0]	caddr;	// Combination of SPI address and back door address
    wire [7:0]	cdata;	// Combination of SPI data and back door data
    wire	cwstb;	// Combination of SPI write strobe and back door write strobe
    wire	csclk;	// Combination of SPI SCK and back door access trigger


	// Output clock signals buffer wires
	wire mgmt_gpio_out_9_prebuff, mgmt_gpio_out_14_prebuff, mgmt_gpio_out_15_prebuff, pad_flash_clk_prebuff;



    // Pass-through mode handling.  Signals may only be applied when the
    // core processor is in reset.

    assign reset = (pass_thru_mgmt_reset) ? 1'b1 : reset_reg;

	// Invert wb_rstn_i
	wire wb_rst_i;
	assign wb_rst_i = ~wb_rstn_i;
	
    // Pass-through mode.  Housekeeping SPI signals get inserted
    // between the management SoC and the flash SPI I/O.
    assign pad_flash_csb = (pass_thru_mgmt_delay) ? mgmt_gpio_in[3] : spimemio_flash_csb;
    assign pad_flash_csb_oeb = (pass_thru_mgmt_delay) ? 1'b0 : (~porb ? 1'b1 : 1'b0);
    assign pad_flash_clk_prebuff = (pass_thru_mgmt) ? mgmt_gpio_in[4] : spimemio_flash_clk;
    assign pad_flash_clk_oeb = (pass_thru_mgmt) ? 1'b0 : (~porb ? 1'b1 : 1'b0);
    assign pad_flash_io0_oeb = (pass_thru_mgmt_delay) ? 1'b0 : spimemio_flash_io0_oeb;
    assign pad_flash_io1_oeb = (pass_thru_mgmt) ? 1'b1 : spimemio_flash_io1_oeb;
    assign pad_flash_io0_ieb = (pass_thru_mgmt_delay) ? 1'b1 : ~spimemio_flash_io0_oeb;
    assign pad_flash_io1_ieb = (pass_thru_mgmt) ? 1'b0 : ~spimemio_flash_io1_oeb;
    assign pad_flash_io0_do = (pass_thru_mgmt_delay) ? mgmt_gpio_in[2] : spimemio_flash_io0_do;
    assign pad_flash_io1_do = spimemio_flash_io1_do;
    assign spimemio_flash_io0_di = (pass_thru_mgmt_delay) ? 1'b0 : pad_flash_io0_di;
    assign spimemio_flash_io1_di = (pass_thru_mgmt) ? 1'b0 : pad_flash_io1_di;

(* keep *) vic_buff_inst pad_flashh_clk_buff_inst (
	.A(pad_flash_clk_prebuff),
    .X(pad_flash_clk));

    wire [11:0] mfgr_id;
    wire [7:0]  prod_id;
    wire [31:0] mask_rev;

    reg serial_busy;

    // Wishbone bus "back door" to SPI registers.  This section of code
    // (1) Maps SPI byte addresses to memory map 32-bit addresses
    // (2) Applies signals to the housekeeping SPI to mux in the SPI address,
    //	   clock, and write strobe.  This is done carefully and slowly to
    //	   avoid glitching on the SCK line and to avoid forcing the
    //	   housekeeping module to keep up with the core clock timing.

    wire      	sys_select;	// System monitoring memory map address selected
    wire      	gpio_select;	// GPIO configuration memory map address selected
    wire      	spi_select;	// SPI back door memory map address selected

    // Wishbone Back Door.  This is a simple interface making use of the
    // housekeeping SPI protocol.  The housekeeping SPI uses byte-wide
    // data, so this interface will stall the processor by holding wb_ack_o
    // low until all bytes have been transferred between the processor and
    // housekeeping SPI.

    reg [3:0] wbbd_state;
    reg [7:0] wbbd_addr;	/* SPI address translated from WB */
    reg [7:0] wbbd_data;	/* SPI data translated from WB */
    reg       wbbd_sck;	    /* wishbone access trigger (back-door clock) */
    reg       wbbd_write;	/* wishbone write trigger (back-door strobe) */
    reg       wbbd_busy;	/* Raised during a wishbone read or write */

    // This defines a state machine that accesses the SPI registers through
    // the back door wishbone interface.  The process is relatively slow
    // since the SPI data are byte-wide, so four individual accesses are
    // made to read 4 bytes from the SPI to fill data on the wishbone bus
    // before sending ACK and letting the processor continue.

    `define WBBD_IDLE	4'h0	/* Back door access is idle */
    `define WBBD_SETUP0	4'h1	/* Apply address and data for byte 1 of 4 */
    `define WBBD_RW0	4'h2	/* Latch data for byte 1 of 4 */
    `define WBBD_SETUP1	4'h3	/* Apply address and data for byte 2 of 4 */
    `define WBBD_RW1	4'h4	/* Latch data for byte 2 of 4 */
    `define WBBD_SETUP2	4'h5	/* Apply address and data for byte 3 of 4 */
    `define WBBD_RW2	4'h6	/* Latch data for byte 3 of 4 */
    `define WBBD_SETUP3	4'h7	/* Apply address and data for byte 4 of 4 */
    `define WBBD_RW3	4'h8	/* Latch data for byte 4 of 4 */
    `define WBBD_DONE	4'h9	/* Send ACK back to wishbone */
    `define WBBD_RESET	4'ha	/* Clock once to reset the transfer bit */

    assign sys_select = (wb_adr_i[31:8] == SYS_BASE_ADR[31:8]);
    assign gpio_select = (wb_adr_i[31:8] == GPIO_BASE_ADR[31:8]);
    assign spi_select = (wb_adr_i[31:8] == SPI_BASE_ADR[31:8]);

    /* Register bit to SPI address mapping */

    function [7:0] fdata(input [7:0] address);
	begin
	case (address)
	    /* Housekeeping SPI Protocol */
	    8'h00 : fdata = 8'h00;			// SPI status (fixed) 

	    /* Status and Identification */
	    8'h01 : fdata = {4'h0, mfgr_id[11:8]};	// Manufacturer ID (fixed)
	    8'h02 : fdata = mfgr_id[7:0];		// Manufacturer ID (fixed)
	    8'h03 : fdata = prod_id;			// Product ID (fixed)
	    8'h04 : fdata = mask_rev[31:24];		// Mask rev (via programmed)
	    8'h05 : fdata = mask_rev[23:16];		// Mask rev (via programmed)
	    8'h06 : fdata = mask_rev[15:8];		// Mask rev (via programmed)
	    8'h07 : fdata = mask_rev[7:0];		// Mask rev (via programmed)

		// [Vic]: Remove PLL signals
	    /* Clocking control */
	    //8'h08 : fdata = {6'b000000, pll_dco_ena, pll_ena};
	    //8'h09 : fdata = {7'b0000000, pll_bypass};
	    8'h0a : fdata = {7'b0000000, irq_spi};
	    8'h0b : fdata = {7'b0000000, reset};
	    8'h0c : fdata = {7'b0000000, trap};		// CPU trap state
	    //8'h0d : fdata = pll_trim[7:0];
	    //8'h0e : fdata = pll_trim[15:8];
	    //8'h0f : fdata = pll_trim[23:16];
	    //8'h10 : fdata = {6'b000000, pll_trim[25:24]};
	    //8'h11 : fdata = {2'b00, pll90_sel, pll_sel};
	    //8'h12 : fdata = {3'b000, pll_div};

	    // GPIO Control (bit bang and automatic)
	    // NOTE: "serial_busy" is the read-back signal occupying the same
	    // address/bit as "serial_xfer".
	    8'h13 : fdata = {1'b0, serial_data_2, serial_data_1, serial_bb_clock,
				serial_bb_load, serial_bb_resetn, serial_bb_enable,
				serial_busy};
		
		default: fdata = 8'h00;


	    /* System monitoring */
	    8'h1a : fdata = {4'b0000, usr1_vcc_pwrgood, usr2_vcc_pwrgood,
				usr1_vdd_pwrgood, usr2_vdd_pwrgood};
	    8'h1b : fdata = {5'b00000, clk1_output_dest, clk2_output_dest,
				trap_output_dest};
	    8'h1c : fdata = {6'b000000, irq_2_inputsrc, irq_1_inputsrc};

	    /* GPIO Configuration */
	    8'h1d : fdata = {3'b000, gpio_configure[0][12:8]};
	    8'h1e : fdata = gpio_configure[0][7:0];
	    8'h1f : fdata = {3'b000, gpio_configure[1][12:8]};
	    8'h20 : fdata = gpio_configure[1][7:0];
	    8'h21 : fdata = {3'b000, gpio_configure[2][12:8]};
	    8'h22 : fdata = gpio_configure[2][7:0];
	    8'h23 : fdata = {3'b000, gpio_configure[3][12:8]};
	    8'h24 : fdata = gpio_configure[3][7:0];
	    8'h25 : fdata = {3'b000, gpio_configure[4][12:8]};
	    8'h26 : fdata = gpio_configure[4][7:0];
	    8'h27 : fdata = {3'b000, gpio_configure[5][12:8]};
	    8'h28 : fdata = gpio_configure[5][7:0];
	    8'h29 : fdata = {3'b000, gpio_configure[6][12:8]};
	    8'h2a : fdata = gpio_configure[6][7:0];
	    8'h2b : fdata = {3'b000, gpio_configure[7][12:8]};
	    8'h2c : fdata = gpio_configure[7][7:0];
	    8'h2d : fdata = {3'b000, gpio_configure[8][12:8]};
	    8'h2e : fdata = gpio_configure[8][7:0];
	    8'h2f : fdata = {3'b000, gpio_configure[9][12:8]};
	    8'h30 : fdata = gpio_configure[9][7:0];
	    8'h31 : fdata = {3'b000, gpio_configure[10][12:8]};
	    8'h32 : fdata = gpio_configure[10][7:0];
	    8'h33 : fdata = {3'b000, gpio_configure[11][12:8]};
	    8'h34 : fdata = gpio_configure[11][7:0];
	    8'h35 : fdata = {3'b000, gpio_configure[12][12:8]};
	    8'h36 : fdata = gpio_configure[12][7:0];
	    8'h37 : fdata = {3'b000, gpio_configure[13][12:8]};
	    8'h38 : fdata = gpio_configure[13][7:0];
	    8'h39 : fdata = {3'b000, gpio_configure[14][12:8]};
	    8'h3a : fdata = gpio_configure[14][7:0];
	    8'h3b : fdata = {3'b000, gpio_configure[15][12:8]};
	    8'h3c : fdata = gpio_configure[15][7:0];
	    8'h3d : fdata = {3'b000, gpio_configure[16][12:8]};
	    8'h3e : fdata = gpio_configure[16][7:0];
	    8'h3f : fdata = {3'b000, gpio_configure[17][12:8]};
	    8'h40 : fdata = gpio_configure[17][7:0];
	    8'h41 : fdata = {3'b000, gpio_configure[18][12:8]};
	    8'h42 : fdata = gpio_configure[18][7:0];
	    8'h43 : fdata = {3'b000, gpio_configure[19][12:8]};
	    8'h44 : fdata = gpio_configure[19][7:0];
	    8'h45 : fdata = {3'b000, gpio_configure[20][12:8]};
	    8'h46 : fdata = gpio_configure[20][7:0];
	    8'h47 : fdata = {3'b000, gpio_configure[21][12:8]};
	    8'h48 : fdata = gpio_configure[21][7:0];
	    8'h49 : fdata = {3'b000, gpio_configure[22][12:8]};
	    8'h4a : fdata = gpio_configure[22][7:0];
	    8'h4b : fdata = {3'b000, gpio_configure[23][12:8]};
	    8'h4c : fdata = gpio_configure[23][7:0];
	    8'h4d : fdata = {3'b000, gpio_configure[24][12:8]};
	    8'h4e : fdata = gpio_configure[24][7:0];
	    8'h4f : fdata = {3'b000, gpio_configure[25][12:8]};
	    8'h50 : fdata = gpio_configure[25][7:0];
	    8'h51 : fdata = {3'b000, gpio_configure[26][12:8]};
	    8'h52 : fdata = gpio_configure[26][7:0];
	    8'h53 : fdata = {3'b000, gpio_configure[27][12:8]};
	    8'h54 : fdata = gpio_configure[27][7:0];
	    8'h55 : fdata = {3'b000, gpio_configure[28][12:8]};
	    8'h56 : fdata = gpio_configure[28][7:0];
	    8'h57 : fdata = {3'b000, gpio_configure[29][12:8]};
	    8'h58 : fdata = gpio_configure[29][7:0];
	    8'h59 : fdata = {3'b000, gpio_configure[30][12:8]};
	    8'h5a : fdata = gpio_configure[30][7:0];
	    8'h5b : fdata = {3'b000, gpio_configure[31][12:8]};
	    8'h5c : fdata = gpio_configure[31][7:0];
	    8'h5d : fdata = {3'b000, gpio_configure[32][12:8]};
	    8'h5e : fdata = gpio_configure[32][7:0];
	    8'h5f : fdata = {3'b000, gpio_configure[33][12:8]};
	    8'h60 : fdata = gpio_configure[33][7:0];
	    8'h61 : fdata = {3'b000, gpio_configure[34][12:8]};
	    8'h62 : fdata = gpio_configure[34][7:0];
	    8'h63 : fdata = {3'b000, gpio_configure[35][12:8]};
	    8'h64 : fdata = gpio_configure[35][7:0];
	    8'h65 : fdata = {3'b000, gpio_configure[36][12:8]};
	    8'h66 : fdata = gpio_configure[36][7:0];
	    8'h67 : fdata = {3'b000, gpio_configure[37][12:8]};
	    8'h68 : fdata = gpio_configure[37][7:0];

	    // GPIO Data
	    8'h69 : fdata = {2'b00, mgmt_gpio_in[`MPRJ_IO_PADS-1:32]};
	    8'h6a : fdata = mgmt_gpio_in[31:24];
	    8'h6b : fdata = mgmt_gpio_in[23:16];
	    8'h6c : fdata = mgmt_gpio_in[15:8];
	    8'h6d : fdata = mgmt_gpio_in[7:0];

	    // Power Control (reserved)
	    8'h6e : fdata = {4'b0000, pwr_ctrl_out};

	    // Housekeeping SPI system disable
	    8'h6f : fdata = {7'b0000000, hkspi_disable};

	endcase
	end
    endfunction

    /* Memory map address to SPI address translation for back door access */
    /* (see doc/memory_map.txt)						  */

    wire [11:0] gpio_adr = GPIO_BASE_ADR[23:12];
    wire [11:0] sys_adr = SYS_BASE_ADR[23:12];
    wire [11:0] spi_adr = SPI_BASE_ADR[23:12];

    function [7:0] spiaddr(input [31:0] wbaddress);
	begin
	/* Address taken from lower 8 bits and upper 4 bits of the 32-bit */
	/* wishbone address.						  */
	case ({wbaddress[23:20], wbaddress[7:0]})
	    spi_adr  | 12'h000 : spiaddr = 8'h00;	// SPI status (reserved)
	    spi_adr  | 12'h004 : spiaddr = 8'h03;	// product ID
	    spi_adr  | 12'h005 : spiaddr = 8'h02;	// Manufacturer ID (low)
	    spi_adr  | 12'h006 : spiaddr = 8'h01;	// Manufacturer ID (high)
	    spi_adr  | 12'h008 : spiaddr = 8'h07;	// User project ID (low)
	    spi_adr  | 12'h009 : spiaddr = 8'h06;	// User project ID .
	    spi_adr  | 12'h00a : spiaddr = 8'h05;	// User project ID .
	    spi_adr  | 12'h00b : spiaddr = 8'h04;	// User project ID (high)

	    spi_adr  | 12'h00c : spiaddr = 8'h08;	// PLL enables
	    spi_adr  | 12'h010 : spiaddr = 8'h09;	// PLL bypass
	    spi_adr  | 12'h014 : spiaddr = 8'h0a;	// IRQ
	    spi_adr  | 12'h018 : spiaddr = 8'h0b;	// Reset
	    spi_adr  | 12'h028 : spiaddr = 8'h0c;	// CPU trap state
	    spi_adr  | 12'h01f : spiaddr = 8'h10;	// PLL trim
	    spi_adr  | 12'h01e : spiaddr = 8'h0f;	// PLL trim
	    spi_adr  | 12'h01d : spiaddr = 8'h0e;	// PLL trim
	    spi_adr  | 12'h01c : spiaddr = 8'h0d;	// PLL trim
	    spi_adr  | 12'h020 : spiaddr = 8'h11;	// PLL source
	    spi_adr  | 12'h024 : spiaddr = 8'h12;	// PLL divider

	    spi_adr  | 12'h02c : spiaddr = 8'h19;	// SRAM read-only data
	    spi_adr  | 12'h02d : spiaddr = 8'h18;	// SRAM read-only data
	    spi_adr  | 12'h02e : spiaddr = 8'h17;	// SRAM read-only data
	    spi_adr  | 12'h02f : spiaddr = 8'h16;	// SRAM read-only data
	    spi_adr  | 12'h030 : spiaddr = 8'h15;	// SRAM read-only address
	    spi_adr  | 12'h034 : spiaddr = 8'h14;	// SRAM read-only control

	    gpio_adr | 12'h000 : spiaddr = 8'h13;	// GPIO control

	    sys_adr  | 12'h000 : spiaddr = 8'h1a;	// Power monitor
	    sys_adr  | 12'h004 : spiaddr = 8'h1b;	// Output redirect
	    sys_adr  | 12'h00c : spiaddr = 8'h1c;	// Input redirect

	    gpio_adr | 12'h025 : spiaddr = 8'h1d;	// GPIO configuration
	    gpio_adr | 12'h024 : spiaddr = 8'h1e;
	    gpio_adr | 12'h029 : spiaddr = 8'h1f;
	    gpio_adr | 12'h028 : spiaddr = 8'h20;
	    gpio_adr | 12'h02d : spiaddr = 8'h21;
	    gpio_adr | 12'h02c : spiaddr = 8'h22;
	    gpio_adr | 12'h031 : spiaddr = 8'h23;
	    gpio_adr | 12'h030 : spiaddr = 8'h24;
	    gpio_adr | 12'h035 : spiaddr = 8'h25;
	    gpio_adr | 12'h034 : spiaddr = 8'h26;
	    gpio_adr | 12'h039 : spiaddr = 8'h27;
	    gpio_adr | 12'h038 : spiaddr = 8'h28;
	    gpio_adr | 12'h03d : spiaddr = 8'h29;
	    gpio_adr | 12'h03c : spiaddr = 8'h2a;
	    gpio_adr | 12'h041 : spiaddr = 8'h2b;
	    gpio_adr | 12'h040 : spiaddr = 8'h2c;
	    gpio_adr | 12'h045 : spiaddr = 8'h2d;
	    gpio_adr | 12'h044 : spiaddr = 8'h2e;
	    gpio_adr | 12'h049 : spiaddr = 8'h2f;
	    gpio_adr | 12'h048 : spiaddr = 8'h30;
	    gpio_adr | 12'h04d : spiaddr = 8'h31;
	    gpio_adr | 12'h04c : spiaddr = 8'h32;
	    gpio_adr | 12'h051 : spiaddr = 8'h33;
	    gpio_adr | 12'h050 : spiaddr = 8'h34;
	    gpio_adr | 12'h055 : spiaddr = 8'h35;
	    gpio_adr | 12'h054 : spiaddr = 8'h36;
	    gpio_adr | 12'h059 : spiaddr = 8'h37;
	    gpio_adr | 12'h058 : spiaddr = 8'h38;
	    gpio_adr | 12'h05d : spiaddr = 8'h39;
	    gpio_adr | 12'h05c : spiaddr = 8'h3a;
	    gpio_adr | 12'h061 : spiaddr = 8'h3b;
	    gpio_adr | 12'h060 : spiaddr = 8'h3c;
	    gpio_adr | 12'h065 : spiaddr = 8'h3d;
	    gpio_adr | 12'h064 : spiaddr = 8'h3e;
	    gpio_adr | 12'h069 : spiaddr = 8'h3f;
	    gpio_adr | 12'h068 : spiaddr = 8'h40;
	    gpio_adr | 12'h06d : spiaddr = 8'h41;
	    gpio_adr | 12'h06c : spiaddr = 8'h42;
	    gpio_adr | 12'h071 : spiaddr = 8'h43;
	    gpio_adr | 12'h070 : spiaddr = 8'h44;
	    gpio_adr | 12'h075 : spiaddr = 8'h45;
	    gpio_adr | 12'h074 : spiaddr = 8'h46;
	    gpio_adr | 12'h079 : spiaddr = 8'h47;
	    gpio_adr | 12'h078 : spiaddr = 8'h48;
	    gpio_adr | 12'h07d : spiaddr = 8'h49;
	    gpio_adr | 12'h07c : spiaddr = 8'h4a;
	    gpio_adr | 12'h081 : spiaddr = 8'h4b;
	    gpio_adr | 12'h080 : spiaddr = 8'h4c;
	    gpio_adr | 12'h085 : spiaddr = 8'h4d;
	    gpio_adr | 12'h084 : spiaddr = 8'h4e;
	    gpio_adr | 12'h089 : spiaddr = 8'h4f;
	    gpio_adr | 12'h088 : spiaddr = 8'h50;
	    gpio_adr | 12'h08d : spiaddr = 8'h51;
	    gpio_adr | 12'h08c : spiaddr = 8'h52;
	    gpio_adr | 12'h091 : spiaddr = 8'h53;
	    gpio_adr | 12'h090 : spiaddr = 8'h54;
	    gpio_adr | 12'h095 : spiaddr = 8'h55;
	    gpio_adr | 12'h094 : spiaddr = 8'h56;
	    gpio_adr | 12'h099 : spiaddr = 8'h57;
	    gpio_adr | 12'h098 : spiaddr = 8'h58;
	    gpio_adr | 12'h09d : spiaddr = 8'h59;
	    gpio_adr | 12'h09c : spiaddr = 8'h5a;
	    gpio_adr | 12'h0a1 : spiaddr = 8'h5b;
	    gpio_adr | 12'h0a0 : spiaddr = 8'h5c;
	    gpio_adr | 12'h0a5 : spiaddr = 8'h5d;
	    gpio_adr | 12'h0a4 : spiaddr = 8'h5e;
	    gpio_adr | 12'h0a9 : spiaddr = 8'h5f;
	    gpio_adr | 12'h0a8 : spiaddr = 8'h60;
	    gpio_adr | 12'h0ad : spiaddr = 8'h61;
	    gpio_adr | 12'h0ac : spiaddr = 8'h62;
	    gpio_adr | 12'h0b1 : spiaddr = 8'h63;
	    gpio_adr | 12'h0b0 : spiaddr = 8'h64;
	    gpio_adr | 12'h0b5 : spiaddr = 8'h65;
	    gpio_adr | 12'h0b4 : spiaddr = 8'h66;
	    gpio_adr | 12'h0b9 : spiaddr = 8'h67;
	    gpio_adr | 12'h0b8 : spiaddr = 8'h68;

	    gpio_adr | 12'h010 : spiaddr = 8'h69;	// GPIO data (h)

	    gpio_adr | 12'h00f : spiaddr = 8'h6a;	// GPIO data (l)
	    gpio_adr | 12'h00e : spiaddr = 8'h6b;	// GPIO data (l)
	    gpio_adr | 12'h00d : spiaddr = 8'h6c;	// GPIO data (l)
	    gpio_adr | 12'h00c : spiaddr = 8'h6d;	// GPIO data (l)

	    gpio_adr | 12'h004 : spiaddr = 8'h6e;	// Power control

	    sys_adr  | 12'h010 : spiaddr = 8'h6f;	// Housekeeping SPI disable

	    default : spiaddr = 8'h00;
	endcase
	end
    endfunction
	
    // SPI is considered active when the GPIO for CSB is set to input and
    // CSB is low.  SPI is considered "busy" when rdstb or wrstb are high,
    // indicating that the SPI will read or write a byte on the next SCK
    // transition.

    wire spi_is_enabled = (~gpio_configure[3][INP_DIS]) & (~hkspi_disable);
    wire spi_is_active = spi_is_enabled && (mgmt_gpio_in[3] == 1'b0);
    wire spi_is_busy = spi_is_active && (rdstb || wrstb);

    /* Wishbone back-door state machine and address translation */

    always @(posedge wb_clk_i or posedge wb_rst_i) begin
	if (wb_rst_i) begin
	    wbbd_sck <= 1'b0;
	    wbbd_write <= 1'b0;
	    wbbd_addr <= 8'd0;
	    wbbd_data <= 8'd0;
	    wbbd_busy <= 1'b0;
	    wb_ack_o <= 1'b0;
	    wbbd_state <= `WBBD_IDLE;
	end else begin
	    case (wbbd_state)
		`WBBD_IDLE: begin
		    wbbd_sck <= 1'b0;
		    wbbd_busy <= 1'b0;
		    if ((sys_select | gpio_select | spi_select) &&
	    	    		 wb_cyc_i && wb_stb_i) begin
			wb_ack_o <= 1'b0;
			wbbd_state <= `WBBD_SETUP0;
		    end
		end
		`WBBD_SETUP0: begin
		    wbbd_sck <= 1'b0;
		    wbbd_addr <= spiaddr(wb_adr_i);
		    if (wb_sel_i[0] & wb_we_i) begin
		    	wbbd_data <= wb_dat_i[7:0];
		    end
		    wbbd_write <= wb_sel_i[0] & wb_we_i;
		    wbbd_busy <= 1'b1;

		    // If the SPI is being accessed and about to read or
		    // write a byte, then stall until the SPI is ready.
		    if (!spi_is_busy) begin
		        wbbd_state <= `WBBD_RW0;
		    end
		end
		`WBBD_RW0: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b1;
		    wb_dat_o[7:0] <= odata;
		    wbbd_state <= `WBBD_SETUP1;
		end
		`WBBD_SETUP1: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b0;
		    wbbd_addr <= spiaddr(wb_adr_i + 1);
		    if (wb_sel_i[1] & wb_we_i) begin
		    	wbbd_data <= wb_dat_i[15:8];
		    end
		    wbbd_write <= wb_sel_i[1] & wb_we_i;
		    if (!spi_is_busy) begin
		        wbbd_state <= `WBBD_RW1;
		    end
		end
		`WBBD_RW1: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b1;
		    wb_dat_o[15:8] <= odata;
		    wbbd_state <= `WBBD_SETUP2;
		end
		`WBBD_SETUP2: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b0;
		    wbbd_addr <= spiaddr(wb_adr_i + 2);
		    if (wb_sel_i[2] & wb_we_i) begin
		    	wbbd_data <= wb_dat_i[23:16];
		    end
		    wbbd_write <= wb_sel_i[2] & wb_we_i;
		    if (!spi_is_busy) begin
		        wbbd_state <= `WBBD_RW2;
		    end
		end
		`WBBD_RW2: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b1;
		    wb_dat_o[23:16] <= odata;
		    wbbd_state <= `WBBD_SETUP3;
		end
		`WBBD_SETUP3: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b0;
		    wbbd_addr <= spiaddr(wb_adr_i + 3);
		    if (wb_sel_i[3] & wb_we_i) begin
		    	wbbd_data <= wb_dat_i[31:24];
		    end
		    wbbd_write <= wb_sel_i[3] & wb_we_i;
		    if (!spi_is_busy) begin
		        wbbd_state <= `WBBD_RW3;
		    end
		end
		`WBBD_RW3: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b1;
		    wb_dat_o[31:24] <= odata;
		    wb_ack_o <= 1'b1;	// Release hold on wishbone bus
		    wbbd_state <= `WBBD_DONE;
		end
		`WBBD_DONE: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b0;
		    wb_ack_o <= 1'b0;	// Reset for next access
		    wbbd_write <= 1'b0;
		    wbbd_state <= `WBBD_RESET;
		end
		`WBBD_RESET: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b1;
		    wb_ack_o <= 1'b0;
		    wbbd_write <= 1'b0;
		    wbbd_state <= `WBBD_IDLE;
		end
	    endcase
	end
    end

    // Instantiate the SPI interface protocol module

    housekeeping_spi hkspi (
		.reset(~porb),
    	.SCK(mgmt_gpio_in[4]),
    	.SDI(mgmt_gpio_in[2]),
    	.CSB((spi_is_enabled) ? mgmt_gpio_in[3] : 1'b1),
    	.SDO(sdo),
    	.sdoenb(sdo_enb),
    	.idata(odata),
    	.odata(idata),
    	.oaddr(iaddr),
    	.rdstb(rdstb),
    	.wrstb(wrstb),
    	.pass_thru_mgmt(pass_thru_mgmt),
    	.pass_thru_mgmt_delay(pass_thru_mgmt_delay),
    	.pass_thru_user(pass_thru_user),
    	.pass_thru_user_delay(pass_thru_user_delay),
    	.pass_thru_mgmt_reset(pass_thru_mgmt_reset),
    	.pass_thru_user_reset(pass_thru_user_reset)
    );



    // GPIO data handling to and from the management SoC

    assign mgmt_gpio_out[37] = (qspi_enabled) ? spimemio_flash_io3_do :
		mgmt_gpio_data[37];
    assign mgmt_gpio_out[36] = (qspi_enabled) ? spimemio_flash_io2_do :
		mgmt_gpio_data[36];

    assign mgmt_gpio_oeb[37] = (qspi_enabled) ? spimemio_flash_io3_oeb :
		~gpio_configure[37][INP_DIS];
    assign mgmt_gpio_oeb[36] = (qspi_enabled) ? spimemio_flash_io2_oeb :
		~gpio_configure[36][INP_DIS];
    assign mgmt_gpio_oeb[35] = (spi_enabled) ? spi_sdoenb :
		~gpio_configure[35][INP_DIS];

    // NOTE:  Ignored by spimemio module when QSPI disabled, so they do not
    // need any exception when qspi_enabled == 1.
    assign spimemio_flash_io3_di = mgmt_gpio_in[37];
    assign spimemio_flash_io2_di = mgmt_gpio_in[36];

    // SPI master is assigned to the other 4 bits of the data high word.
    assign mgmt_gpio_out[32] = (spi_enabled) ? spi_sck : mgmt_gpio_data[32];
    assign mgmt_gpio_out[33] = (spi_enabled) ? spi_csb : mgmt_gpio_data[33];
    assign mgmt_gpio_out[34] = mgmt_gpio_data[34];
    assign mgmt_gpio_out[35] = (spi_enabled) ? spi_sdo : mgmt_gpio_data[35];

    assign mgmt_gpio_out[31:16] = mgmt_gpio_data[31:16];
    assign mgmt_gpio_out[12:11] = mgmt_gpio_data[12:11];

    assign mgmt_gpio_out[10] = (pass_thru_user_delay) ? mgmt_gpio_in[2]
			: mgmt_gpio_data[10];
    assign mgmt_gpio_out_9_prebuff = (pass_thru_user) ? mgmt_gpio_in[4]
			: mgmt_gpio_data[9];

(* keep *) vic_buff_inst mgmt_gpio_9_buff_inst (
	.A(mgmt_gpio_out_9_prebuff),
    .X(mgmt_gpio_out[9]));

    assign mgmt_gpio_out[8] = (pass_thru_user_delay) ? mgmt_gpio_in[3]
			: mgmt_gpio_data[8];

    assign mgmt_gpio_out[7] = mgmt_gpio_data[7];
    assign mgmt_gpio_out[6] = (uart_enabled) ? ser_tx : mgmt_gpio_data[6];
    assign mgmt_gpio_out[5:2] = mgmt_gpio_data[5:2];

    // In pass-through modes, route SDO from the respective flash (user or
    // management SoC) to the dedicated SDO pin (GPIO[1])

    assign mgmt_gpio_out[1] = (pass_thru_mgmt) ? pad_flash_io1_di :
		 (pass_thru_user) ? mgmt_gpio_in[11] :
		 (spi_is_active) ? sdo : mgmt_gpio_data[1];
    assign mgmt_gpio_out[0] = (debug_mode) ? debug_out : mgmt_gpio_data[0];

    assign mgmt_gpio_oeb[1] = (spi_is_active) ? sdo_enb : ~gpio_configure[1][INP_DIS];
    assign mgmt_gpio_oeb[0] = (debug_mode) ? debug_oeb : ~gpio_configure[0][INP_DIS];

    assign ser_rx = (uart_enabled) ? mgmt_gpio_in[5] : 1'b0;
    assign spi_sdi = (spi_enabled) ? mgmt_gpio_in[34] : 1'b0;
    assign debug_in = (debug_mode) ? mgmt_gpio_in[0] : 1'b0;

    genvar i;

    /* These are disconnected, but apply a meaningful signal anyway */
    generate
	for (i = 2; i < `MPRJ_IO_PADS-3; i = i + 1) begin
	    assign mgmt_gpio_oeb[i] = ~gpio_configure[i][INP_DIS];
	end
    endgenerate

    // System monitoring.  Multiplex the clock and trap
    // signals to the associated pad, and multiplex the irq signals
    // from the associated pad, when the redirection is enabled.  Note
    // that the redirection is upstream of the user/managment multiplexing,
    // so the pad being under control of the user area takes precedence
    // over the system monitoring function.

    assign mgmt_gpio_out_15_prebuff = (clk2_output_dest == 1'b1) ? user_clock
		: mgmt_gpio_data[15];

(* keep *) vic_buff_inst mgmt_gpio_15_buff_inst (
	.A(mgmt_gpio_out_15_prebuff),
    .X(mgmt_gpio_out[15]));

    assign mgmt_gpio_out_14_prebuff = (clk1_output_dest == 1'b1) ? wb_clk_i
		: mgmt_gpio_data[14];

(* keep *) vic_buff_inst mgmt_gpio_14_buff_inst (
	.A(mgmt_gpio_out_14_prebuff),
    .X(mgmt_gpio_out[14]));

    assign mgmt_gpio_out[13] = (trap_output_dest == 1'b1) ? trap
		: mgmt_gpio_data[13];

    assign irq[0] = irq_spi;
    assign irq[1] = (irq_1_inputsrc == 1'b1) ? mgmt_gpio_in[7] : 1'b0;
    assign irq[2] = (irq_2_inputsrc == 1'b1) ? mgmt_gpio_in[12] : 1'b0;

    // GPIO serial loader and GPIO management control

`define GPIO_IDLE	2'b00
`define GPIO_START	2'b01
`define GPIO_XBYTE	2'b10
`define GPIO_LOAD	2'b11

    reg [3:0]	xfer_count;
    reg [4:0]	pad_count_1;
    reg [5:0]	pad_count_2;
    reg [1:0]	xfer_state;

    reg serial_clock_pre;
    reg serial_resetn_pre;
    reg serial_load_pre;
    reg [IO_CTRL_BITS-1:0] serial_data_staging_1;
    reg [IO_CTRL_BITS-1:0] serial_data_staging_2;

    assign serial_clock = (serial_bb_enable == 1'b1) ?
			serial_bb_clock : serial_clock_pre;
    assign serial_resetn = (serial_bb_enable == 1'b1) ?
			serial_bb_resetn : serial_resetn_pre;
    assign serial_load = (serial_bb_enable == 1'b1) ?
			serial_bb_load : serial_load_pre;

    assign serial_data_1 = (serial_bb_enable == 1'b1) ?
			serial_bb_data_1 : serial_data_staging_1[IO_CTRL_BITS-1];
    assign serial_data_2 = (serial_bb_enable == 1'b1) ?
			serial_bb_data_2 : serial_data_staging_2[IO_CTRL_BITS-1];

    always @(posedge wb_clk_i or negedge porb) begin
	if (porb == 1'b0) begin
	    xfer_state <= `GPIO_IDLE;
	    xfer_count <= 4'd0;
            /* NOTE:  This assumes that MPRJ_IO_PADS_1 and MPRJ_IO_PADS_2 are
             * equal, because they get clocked the same number of cycles by
             * the same clock signal.  pad_count_2 gates the count for both.
             */
	    pad_count_1 <= `MPRJ_IO_PADS_1 - 1;
	    pad_count_2 <= `MPRJ_IO_PADS_1;
	    serial_resetn_pre <= 1'b0;
	    serial_clock_pre <= 1'b0;
	    serial_load_pre <= 1'b0;
	    serial_data_staging_1 <= 0;
	    serial_data_staging_2 <= 0;
	    serial_busy <= 1'b0;

	end else begin

            serial_resetn_pre <= 1'b1;
	    case (xfer_state)
		`GPIO_IDLE: begin
		    pad_count_1 <= `MPRJ_IO_PADS_1 - 1;
                    pad_count_2 <= `MPRJ_IO_PADS_1;
                    serial_clock_pre <= 1'b0;
                    serial_load_pre <= 1'b0;
                    if (serial_xfer == 1'b1) begin
                        xfer_state <= `GPIO_START;
	    	    	serial_busy <= 1'b1;
                    end else begin
	    	    	serial_busy <= 1'b0;
		    end
		end
		`GPIO_START: begin
                    serial_clock_pre <= 1'b0;
                    serial_load_pre <= 1'b0;
                    xfer_count <= 6'd0;
                    pad_count_1 <= pad_count_1 - 1;
                    pad_count_2 <= pad_count_2 + 1;
                    xfer_state <= `GPIO_XBYTE;
                    serial_data_staging_1 <= gpio_configure[pad_count_1];
                    serial_data_staging_2 <= gpio_configure[pad_count_2];
		end
		`GPIO_XBYTE: begin
                    serial_clock_pre <= ~serial_clock;
                    serial_load_pre <= 1'b0;
                    if (serial_clock == 1'b0) begin
                        if (xfer_count == IO_CTRL_BITS - 1) begin
                            xfer_count <= 4'd0;
                            if (pad_count_2 == `MPRJ_IO_PADS) begin
                                xfer_state <= `GPIO_LOAD;
                            end else begin
                                xfer_state <= `GPIO_START;
                            end
                        end else begin
                            xfer_count <= xfer_count + 1;
                        end
                    end else begin
                        serial_data_staging_1 <=
				{serial_data_staging_1[IO_CTRL_BITS-2:0], 1'b0};
                        serial_data_staging_2 <=
				{serial_data_staging_2[IO_CTRL_BITS-2:0], 1'b0};
                    end
		end
		`GPIO_LOAD: begin
                    xfer_count <= xfer_count + 1;

                    /* Load sequence:  Pulse clock for final data shift in;
                     * Pulse the load strobe.
                     * Return to idle mode.
                     */
                    if (xfer_count == 4'd0) begin
                        serial_clock_pre <= 1'b0;
                        serial_load_pre <= 1'b0;
                    end else if (xfer_count == 4'd1) begin
                        serial_clock_pre <= 1'b0;
                        serial_load_pre <= 1'b1;
                    end else if (xfer_count == 4'd2) begin
	    	    	serial_busy <= 1'b0;
                        serial_clock_pre <= 1'b0;
                        serial_load_pre <= 1'b0;
                        xfer_state <= `GPIO_IDLE;
		    end
                end
            endcase
	end
    end

    // SPI Identification

    assign mfgr_id = 12'h456;		// Hard-coded
    assign prod_id = 8'h11;		// Hard-coded
    assign mask_rev = mask_rev_in;	// Copy in to out.

    // SPI Data transfer protocol.  The wishbone back door may only be
    // used if the front door is closed (CSB is high or the CSB pin is
    // not an input).  The time to apply values for the back door access
    // is limited to the clock cycle around the read or write from the
    // wbbd state machine (see below).

    assign caddr = (wbbd_busy) ? wbbd_addr : iaddr;
    //assign csclk = (wbbd_busy) ? wbbd_sck : ((spi_is_active) ? mgmt_gpio_in[4] : 1'b0); // synopsys infer_mux
    //(* keep = "ture" *) assign csclk = (wbbd_busy) ? wbbd_sck : ((spi_is_active) ? mgmt_gpio_in[4] : 1'b0);
    //assign csclk = (wbbd_busy) ? wbbd_sck : ((spi_is_active) ? mgmt_gpio_in[4] : 1'b0);

    // use a MUX instance for create_generated_clock in sdc
    wire tmp_hkspi_clk;
    assign tmp_hkspi_clk = (spi_is_active) ? mgmt_gpio_in[4] : 1'b0;
    //assign csclk = (wbbd_busy) ? wbbd_sck : tmp_hkspi_clk;
   
	clkmux csclk_MUX_dont_touch (
        .A(tmp_hkspi_clk),
        .B(wbbd_sck),
        .S0(wbbd_busy),
        .Y(csclk)
	);

    assign cdata = (wbbd_busy) ? wbbd_data : idata;
    assign cwstb = (wbbd_busy) ? wbbd_write : wrstb;

    assign odata = fdata(caddr);

    // Register mapping and I/O to SPI interface module

    integer j;

    always @(posedge csclk or negedge porb) begin
	if (porb == 1'b0) begin
            // Set trim for PLL at (almost) slowest rate (~90MHz).  However,
            // pll_trim[12] must be set to zero for proper startup.
			///////////////////////////////////////////////////////////////////////
			// [Vic]: Remove PLL signals
            // pll_trim <= 26'b11111111111110111111111111;
            // pll_sel <= 3'b010;		// Default output divider divide-by-2
            // pll90_sel <= 3'b010;	// Default secondary output divider divide-by-2
            // pll_div <= 5'b00100;	// Default feedback divider divide-by-8
            // pll_dco_ena <= 1'b1;	// Default free-running PLL
            // pll_ena <= 1'b0;		// Default PLL turned off
            // pll_bypass <= 1'b1;		// Default bypass mode (don't use PLL)
			///////////////////////////////////////////////////////////////////////
            irq_spi <= 1'b0;
            reset_reg <= 1'b0;

	    // System monitoring signals
	    clk1_output_dest <= 1'b0;
	    clk2_output_dest <= 1'b0;
	    trap_output_dest <= 1'b0;
	    irq_1_inputsrc <= 1'b0;
	    irq_2_inputsrc <= 1'b0;

	    // GPIO Configuration, Data, and Control
	    // To-do:  Get user project pad defaults from external inputs
	    // to be configured by user or at project generation time.
	    // Pads 1 to 4 are the SPI and considered critical startup
	    // infrastructure, and should not be altered from the defaults
	    // below.  NOTE:  These are not startup values, but they should
	    // match the startup values applied to the GPIO, or else the
	    // GPIO should be always triggered to load at startup.

	    for (j = 0; j < `MPRJ_IO_PADS; j=j+1) begin
		if ((j < 2) || (j >= `MPRJ_IO_PADS - 2)) begin
		    gpio_configure[j] <= 'h1803;
                end else begin
		    if (j == 3) begin
			// j == 3 corresponds to CSB, which is a weak pull-up
	                gpio_configure[j] <= 'h0801;
		    end else begin
	                gpio_configure[j] <= 'h0403;
		    end
		end
	    end

	    mgmt_gpio_data <= 'd0;
	    mgmt_gpio_data_buf <= 'd0;
	    serial_bb_enable <= 1'b0;
	    serial_bb_load <= 1'b0;
	    serial_bb_data_1 <= 1'b0;
	    serial_bb_data_2 <= 1'b0;
	    serial_bb_clock <= 1'b0;
	    serial_bb_resetn <= 1'b0;
	    serial_xfer <= 1'b0;
	    hkspi_disable <= 1'b0;
	    pwr_ctrl_out <= 'd0;

        end else begin
	    if (cwstb == 1'b1) begin
                case (caddr)
	    	    /* Register 8'h00 is reserved for future use */
	    	    /* Registers 8'h01 to 8'h07 are read-only and cannot be written */
			///////////////////////////////////////////////////////////////////////
			// [Vic]: Remove PLL signals
            	    // 8'h08: begin
                	// pll_ena <= cdata[0];
                	// pll_dco_ena <= cdata[1];
            	    // end
            	    // 8'h09: begin
                	// pll_bypass <= cdata[0];
            	    // end
            	    8'h0a: begin
                	irq_spi <= cdata[0];
            	    end
            	    8'h0b: begin
                	reset_reg <= cdata[0];
            	    end

		    /* Register 0c (trap state) is read-only */

            	    // 8'h0d: begin
                	// pll_trim[7:0] <= cdata;
            	    // end
            	    // 8'h0e: begin
                	// pll_trim[15:8] <= cdata;
            	    // end
            	    // 8'h0f: begin
                	// pll_trim[23:16] <= cdata;
            	    // end
            	    // 8'h10: begin
                	// pll_trim[25:24] <= cdata[1:0];
            	    // end
            	    // 8'h11: begin
                	// pll90_sel <= cdata[5:3];
                	// pll_sel <= cdata[2:0];
            	    // end
            	    // 8'h12: begin
                	// pll_div <= cdata[4:0];
            	    // end
			///////////////////////////////////////////////////////////////////////
	    	    8'h13: begin
			serial_bb_data_2 <= cdata[6];
			serial_bb_data_1 <= cdata[5];
			serial_bb_clock  <= cdata[4];
			serial_bb_load   <= cdata[3];
			serial_bb_resetn <= cdata[2];
			serial_bb_enable <= cdata[1];
			serial_xfer <= cdata[0];
	    	    end
		    
		    /* Registers 16 to 19 (SRAM data) are read-only */

		    /* Register 1a (power monitor) is read-only */

            	    8'h1b: begin
			clk1_output_dest <= cdata[2];
			clk2_output_dest <= cdata[1];
			trap_output_dest <= cdata[0];
	    	    end
            	    8'h1c: begin
			irq_2_inputsrc <= cdata[1];
			irq_1_inputsrc <= cdata[0];
	    	    end
            	    8'h1d: begin
			gpio_configure[0][12:8] <= cdata[4:0];
	    	    end
            	    8'h1e: begin
			gpio_configure[0][7:0] <= cdata;
	    	    end
            	    8'h1f: begin
			gpio_configure[1][12:8] <= cdata[4:0];
	    	    end
            	    8'h20: begin
			gpio_configure[1][7:0] <= cdata;
	    	    end
            	    8'h21: begin
			gpio_configure[2][12:8] <= cdata[4:0];
	    	    end
            	    8'h22: begin
			gpio_configure[2][7:0] <= cdata;
	    	    end
            	    8'h23: begin
			gpio_configure[3][12:8] <= cdata[4:0];
	    	    end
            	    8'h24: begin
			gpio_configure[3][7:0] <= cdata;
	    	    end
            	    8'h25: begin
			gpio_configure[4][12:8] <= cdata[4:0];
	    	    end
            	    8'h26: begin
			gpio_configure[4][7:0] <= cdata;
	    	    end
            	    8'h27: begin
			gpio_configure[5][12:8] <= cdata[4:0];
	    	    end
            	    8'h28: begin
			gpio_configure[5][7:0] <= cdata;
	    	    end
            	    8'h29: begin
			gpio_configure[6][12:8] <= cdata[4:0];
	    	    end
            	    8'h2a: begin
			gpio_configure[6][7:0] <= cdata;
	    	    end
            	    8'h2b: begin
			gpio_configure[7][12:8] <= cdata[4:0];
	    	    end
            	    8'h2c: begin
			gpio_configure[7][7:0] <= cdata;
	    	    end
            	    8'h2d: begin
			gpio_configure[8][12:8] <= cdata[4:0];
	    	    end
            	    8'h2e: begin
			gpio_configure[8][7:0] <= cdata;
	    	    end
            	    8'h2f: begin
			gpio_configure[9][12:8] <= cdata[4:0];
	    	    end
            	    8'h30: begin
			gpio_configure[9][7:0] <= cdata;
	    	    end
            	    8'h31: begin
			gpio_configure[10][12:8] <= cdata[4:0];
	    	    end
            	    8'h32: begin
			gpio_configure[10][7:0] <= cdata;
	    	    end
            	    8'h33: begin
			gpio_configure[11][12:8] <= cdata[4:0];
	    	    end
            	    8'h34: begin
			gpio_configure[11][7:0] <= cdata;
	    	    end
            	    8'h35: begin
			gpio_configure[12][12:8] <= cdata[4:0];
	    	    end
            	    8'h36: begin
			gpio_configure[12][7:0] <= cdata;
	    	    end
            	    8'h37: begin
			gpio_configure[13][12:8] <= cdata[4:0];
	    	    end
            	    8'h38: begin
			gpio_configure[13][7:0] <= cdata;
	    	    end
            	    8'h39: begin
			gpio_configure[14][12:8] <= cdata[4:0];
	    	    end
            	    8'h3a: begin
			gpio_configure[14][7:0] <= cdata;
	    	    end
            	    8'h3b: begin
			gpio_configure[15][12:8] <= cdata[4:0];
	    	    end
            	    8'h3c: begin
			gpio_configure[15][7:0] <= cdata;
	    	    end
            	    8'h3d: begin
			gpio_configure[16][12:8] <= cdata[4:0];
	    	    end
            	    8'h3e: begin
			gpio_configure[16][7:0] <= cdata;
	    	    end
            	    8'h3f: begin
			gpio_configure[17][12:8] <= cdata[4:0];
	    	    end
            	    8'h40: begin
			gpio_configure[17][7:0] <= cdata;
	    	    end
            	    8'h41: begin
			gpio_configure[18][12:8] <= cdata[4:0];
	    	    end
            	    8'h42: begin
			gpio_configure[18][7:0] <= cdata;
	    	    end
            	    8'h43: begin
			gpio_configure[19][12:8] <= cdata[4:0];
	    	    end
            	    8'h44: begin
			gpio_configure[19][7:0] <= cdata;
	    	    end
            	    8'h45: begin
			gpio_configure[20][12:8] <= cdata[4:0];
	    	    end
            	    8'h46: begin
			gpio_configure[20][7:0] <= cdata;
	    	    end
            	    8'h47: begin
			gpio_configure[21][12:8] <= cdata[4:0];
	    	    end
            	    8'h48: begin
			gpio_configure[21][7:0] <= cdata;
	    	    end
            	    8'h49: begin
			gpio_configure[22][12:8] <= cdata[4:0];
	    	    end
            	    8'h4a: begin
			gpio_configure[22][7:0] <= cdata;
	    	    end
            	    8'h4b: begin
			gpio_configure[23][12:8] <= cdata[4:0];
	    	    end
            	    8'h4c: begin
			gpio_configure[23][7:0] <= cdata;
	    	    end
            	    8'h4d: begin
			gpio_configure[24][12:8] <= cdata[4:0];
	    	    end
            	    8'h4e: begin
			gpio_configure[24][7:0] <= cdata;
	    	    end
            	    8'h4f: begin
			gpio_configure[25][12:8] <= cdata[4:0];
	    	    end
            	    8'h50: begin
			gpio_configure[25][7:0] <= cdata;
	    	    end
            	    8'h51: begin
			gpio_configure[26][12:8] <= cdata[4:0];
	    	    end
            	    8'h52: begin
			gpio_configure[26][7:0] <= cdata;
	    	    end
            	    8'h53: begin
			gpio_configure[27][12:8] <= cdata[4:0];
	    	    end
            	    8'h54: begin
			gpio_configure[27][7:0] <= cdata;
	    	    end
            	    8'h55: begin
			gpio_configure[28][12:8] <= cdata[4:0];
	    	    end
            	    8'h56: begin
			gpio_configure[28][7:0] <= cdata;
	    	    end
            	    8'h57: begin
			gpio_configure[29][12:8] <= cdata[4:0];
	    	    end
            	    8'h58: begin
			gpio_configure[29][7:0] <= cdata;
	    	    end
            	    8'h59: begin
			gpio_configure[30][12:8] <= cdata[4:0];
	    	    end
            	    8'h5a: begin
			gpio_configure[30][7:0] <= cdata;
	    	    end
            	    8'h5b: begin
			gpio_configure[31][12:8] <= cdata[4:0];
	    	    end
            	    8'h5c: begin
			gpio_configure[31][7:0] <= cdata;
	    	    end
            	    8'h5d: begin
			gpio_configure[32][12:8] <= cdata[4:0];
	    	    end
            	    8'h5e: begin
			gpio_configure[32][7:0] <= cdata;
	    	    end
            	    8'h5f: begin
			gpio_configure[33][12:8] <= cdata[4:0];
	    	    end
            	    8'h60: begin
			gpio_configure[33][7:0] <= cdata;
	    	    end
            	    8'h61: begin
			gpio_configure[34][12:8] <= cdata[4:0];
	    	    end
            	    8'h62: begin
			gpio_configure[34][7:0] <= cdata;
	    	    end
            	    8'h63: begin
			gpio_configure[35][12:8] <= cdata[4:0];
	    	    end
            	    8'h64: begin
			gpio_configure[35][7:0] <= cdata;
	    	    end
            	    8'h65: begin
			gpio_configure[36][12:8] <= cdata[4:0];
	    	    end
            	    8'h66: begin
			gpio_configure[36][7:0] <= cdata;
	    	    end
            	    8'h67: begin
			gpio_configure[37][12:8] <= cdata[4:0];
	    	    end
            	    8'h68: begin
			gpio_configure[37][7:0] <= cdata;
	    	    end
	    	    8'h69: begin
			mgmt_gpio_data[37:32] <= cdata[5:0];
	    	    end
	    	    8'h6a: begin
			/* NOTE: mgmt_gpio_data updates only on the	*/
			/* upper byte write when writing through the	*/
			/* wishbone back-door.  This lets all bits	*/
			/* update at the same time.			*/
			if (spi_is_active) begin
			    mgmt_gpio_data[31:24] <= cdata;
			end else begin
			    mgmt_gpio_data[31:0] <= {cdata, mgmt_gpio_data_buf};
			end
	    	    end
	    	    8'h6b: begin
			if (spi_is_active) begin
			    mgmt_gpio_data[23:16] <= cdata;
			end else begin
			    mgmt_gpio_data_buf[23:16] <= cdata;
			end
	    	    end
	    	    8'h6c: begin
			if (spi_is_active) begin
			    mgmt_gpio_data[15:8] <= cdata;
			end else begin
			    mgmt_gpio_data_buf[15:8] <= cdata;
			end
	    	    end
	    	    8'h6d: begin
			if (spi_is_active) begin
			    mgmt_gpio_data[7:0] <= cdata;
			end else begin
			    mgmt_gpio_data_buf[7:0] <= cdata;
			end
	    	    end
	    	    8'h6e: begin
			pwr_ctrl_out <= cdata[3:0];
	    	    end
	    	    8'h6f: begin
			hkspi_disable <= cdata[0];
	    	    end
        	endcase	// (caddr)
    	    end else begin
	    	serial_xfer <= 1'b0;	// Serial transfer is self-resetting
		irq_spi <= 1'b0;	// IRQ is self-resetting
    	    end
    	end
    end
endmodule	// housekeeping


module vic_buff_inst (
        input A,
        output wire X );

//wire X;

assign X = A;
endmodule

module clkmux (
       input A,
       input B,
       input S0,
       output Y
       );

       assign Y = (S0)? B : A;

endmodule// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

//`default_nettype none

//-----------------------------------------------------------
// SPI controller for Caravel
//-----------------------------------------------------------
// housekeeping_spi.v
//------------------------------------------------------
// General purpose SPI module for the Caravel chip
//------------------------------------------------------
// Written by Tim Edwards
// efabless, inc., September 28, 2020
//------------------------------------------------
// This file is distributed free and open source
//------------------------------------------------

// SCK ---   Clock input
// SDI ---   Data  input
// SDO ---   Data  output
// CSB ---   Chip  select (sense negative)
// idata --- Data from chip to transmit out, in 8 bits
// odata --- Input data to chip, in 8 bits
// addr  --- Decoded address to upstream circuits
// rdstb --- Read strobe, tells upstream circuit that data will be latched.
// wrstb --- Write strobe, tells upstream circuit to latch odata.

// Data format (general purpose):
// 8 bit format
// 1st byte:   Command word (see below)
// 2nd byte:   Address word (register 0 to 255)
// 3rd byte:   Data word    (value 0 to 255)

// Command format:
// 00000000  No operation
// 10000000  Write until CSB raised
// 01000000  Read  until CSB raised
// 11000000  Simultaneous read/write until CSB raised
// 11000100  Pass-through read/write to management area flash SPI until CSB raised
// 11000010  Pass-through read/write to user area flash SPI until CSB raised
// wrnnn000  Read/write as above, for nnn = 1 to 7 bytes, then terminate

// Lower three bits are reserved for future use.
// All serial bytes are read and written msb first.

// Fixed control and status registers

// Address 0 is reserved and contains flags for SPI mode.  This is
// currently undefined and is always value 0.
// Address 1 is reserved and contains manufacturer ID low 8 bits.
// Address 2 is reserved and contains manufacturer ID high 4 bits.
// Address 3 is reserved and contains product ID (8 bits).
// Addresses 4 to 7 are reserved and contain the mask ID (32 bits).
// Addresses 8 to 255 are available for general purpose use.

`define COMMAND  3'b000
`define ADDRESS  3'b001
`define DATA     3'b010
`define USERPASS 3'b100
`define MGMTPASS 3'b101

module housekeeping_spi(reset, SCK, SDI, CSB, SDO,
	sdoenb, idata, odata, oaddr, rdstb, wrstb,
	pass_thru_mgmt, pass_thru_mgmt_delay,
	pass_thru_user, pass_thru_user_delay,
	pass_thru_mgmt_reset, pass_thru_user_reset);

    input reset;
    input SCK;
    input SDI;
    input CSB;
    output SDO;
    output sdoenb;
    input [7:0] idata;
    output [7:0] odata;
    output [7:0] oaddr;
    output rdstb;
    output wrstb; 
    output pass_thru_mgmt;
    output pass_thru_mgmt_delay;
    output pass_thru_user;
    output pass_thru_user_delay;
    output pass_thru_mgmt_reset;
    output pass_thru_user_reset;

    reg  [7:0]  addr;
    reg		wrstb;
    reg		rdstb;
    reg		sdoenb;
    reg  [2:0]  state;
    reg  [2:0]  count;
    reg		writemode;
    reg		readmode;
    reg  [2:0]	fixed;
    wire [7:0]  odata;
    reg  [6:0]  predata;
    wire [7:0]  oaddr;
    reg  [7:0]  ldata;
    reg		pass_thru_mgmt;
    reg		pass_thru_mgmt_delay;
    reg		pre_pass_thru_mgmt;
    reg		pass_thru_user;
    reg		pass_thru_user_delay;
    reg		pre_pass_thru_user;
    wire	csb_reset;

    assign odata = {predata, SDI};
    assign oaddr = (state == `ADDRESS) ? {addr[6:0], SDI} : addr;
    assign SDO = ldata[7];
    assign csb_reset = CSB | reset;
    assign pass_thru_mgmt_reset = pass_thru_mgmt_delay | pre_pass_thru_mgmt;
    assign pass_thru_user_reset = pass_thru_user_delay | pre_pass_thru_user;

    // Readback data is captured on the falling edge of SCK so that
    // it is guaranteed valid at the next rising edge.
    always @(negedge SCK or posedge csb_reset) begin
        if (csb_reset == 1'b1) begin
            wrstb <= 1'b0;
            ldata  <= 8'b00000000;
            sdoenb <= 1'b1;
        end else begin

            // After CSB low, 1st SCK starts command

            if (state == `DATA) begin
            	if (readmode == 1'b1) begin
                    sdoenb <= 1'b0;
                    if (count == 3'b000) begin
                	ldata <= idata;
                    end else begin
                	ldata <= {ldata[6:0], 1'b0};	// Shift out
                    end
                end else begin
                    sdoenb <= 1'b1;
                end

                // Apply write strobe on SCK negative edge on the next-to-last
                // data bit so that it updates data on the rising edge of SCK
                // on the last data bit.
 
                if (count == 3'b111) begin
                    if (writemode == 1'b1) begin
                        wrstb <= 1'b1;
                    end
                end else begin
                    wrstb <= 1'b0;
                end

	    end else if (state == `MGMTPASS || state == `USERPASS) begin
		wrstb <= 1'b0;
		sdoenb <= 1'b0;
            end else begin
                wrstb <= 1'b0;
                sdoenb <= 1'b1;
            end		// ! state `DATA
        end		// ! csb_reset
    end			// always @ ~SCK

    always @(posedge SCK or posedge csb_reset) begin
        if (csb_reset == 1'b1) begin
            // Default state on reset
            addr <= 8'h00;
	    rdstb <= 1'b0;
            predata <= 7'b0000000;
            state  <= `COMMAND;
            count  <= 3'b000;
            readmode <= 1'b0;
            writemode <= 1'b0;
            fixed <= 3'b000;
	    pass_thru_mgmt <= 1'b0;
	    pass_thru_mgmt_delay <= 1'b0;
	    pre_pass_thru_mgmt <= 1'b0;
	    pass_thru_user <= 1'b0;
	    pass_thru_user_delay <= 1'b0;
	    pre_pass_thru_user <= 1'b0;
        end else begin
            // After csb_reset low, 1st SCK starts command
            if (state == `COMMAND) begin
		rdstb <= 1'b0;
                count <= count + 1;
        	if (count == 3'b000) begin
	            writemode <= SDI;
	        end else if (count == 3'b001) begin
	            readmode <= SDI;
	        end else if (count < 3'b101) begin
	            fixed <= {fixed[1:0], SDI}; 
	        end else if (count == 3'b101) begin
		    pre_pass_thru_mgmt <= SDI;
	        end else if (count == 3'b110) begin
		    pre_pass_thru_user <= SDI;
		    pass_thru_mgmt_delay <= pre_pass_thru_mgmt;
	        end else if (count == 3'b111) begin
		    pass_thru_user_delay <= pre_pass_thru_user;
		    if (pre_pass_thru_mgmt == 1'b1) begin
			state <= `MGMTPASS;
			pre_pass_thru_mgmt <= 1'b0;
		    end else if (pre_pass_thru_user == 1'b1) begin
			state <= `USERPASS;
			pre_pass_thru_user <= 1'b0;
		    end else begin
	                state <= `ADDRESS;
		    end
	        end
            end else if (state == `ADDRESS) begin
	        count <= count + 1;
	        addr <= {addr[6:0], SDI};
	        if (count == 3'b111) begin
	            state <= `DATA;
		    if (readmode == 1'b1) begin
			rdstb <= 1'b1;
		    end
	        end else begin
		    rdstb <= 1'b0;
		end

            end else if (state == `DATA) begin
	        predata <= {predata[6:0], SDI};
	        count <= count + 1;
	        if (count == 3'b111) begin
	            if (fixed == 3'b001) begin
	                state <= `COMMAND;
	            end else if (fixed != 3'b000) begin
	                fixed <= fixed - 1;
	                addr <= addr + 1;	// Auto increment address (fixed)
	            end else begin	
	                addr <= addr + 1;	// Auto increment address (streaming)
	            end
		    if (readmode == 1'b1) begin
			rdstb <= 1'b1;
		    end
	        end else begin
		    rdstb <= 1'b0;
		end
	    end else if (state == `MGMTPASS) begin
		pass_thru_mgmt <= 1'b1;
	    end else if (state == `USERPASS) begin
		pass_thru_user <= 1'b1;
            end		// ! state `DATA | `MGMTPASS | `USERPASS
        end		// ! csb_reset 
    end			// always @ SCK

endmodule // housekeeping_spi
//`default_nettype wire
//--------------------------------------------------------------------------------
// Auto-generated by Migen (9a0be7a) & LiteX (470fc6f) on 2022-10-14 12:53:55
//--------------------------------------------------------------------------------
module mgmt_core(
	input wire core_clk,
	input wire core_rstn,
	output wire flash_cs_n,
	output reg flash_clk,
	output reg flash_io0_oeb,
	output wire flash_io1_oeb,
	output wire flash_io2_oeb,
	output wire flash_io3_oeb,
	output reg flash_io0_do,
	output wire flash_io1_do,
	output wire flash_io2_do,
	output wire flash_io3_do,
	input wire flash_io0_di,
	input wire flash_io1_di,
	input wire flash_io2_di,
	input wire flash_io3_di,
	output reg spi_clk,
	output reg spi_cs_n,
	output reg spi_mosi,
	input wire spi_miso,
	output wire spi_sdoenb,
	output wire mprj_wb_iena,
	output wire mprj_cyc_o,
	output wire mprj_stb_o,
	output wire mprj_we_o,
	output wire [3:0] mprj_sel_o,
	output reg [31:0] mprj_adr_o,
	output wire [31:0] mprj_dat_o,
	input wire [31:0] mprj_dat_i,
	input wire mprj_ack_i,
	input wire [31:0] hk_dat_i,
	output wire hk_stb_o,
	output wire hk_cyc_o,
	input wire hk_ack_i,
	output reg serial_tx,
	input wire serial_rx,
	input wire debug_in,
	output wire debug_out,
	output wire debug_oeb,
	output wire debug_mode,
	output wire uart_enabled,
	output wire gpio_out_pad,
	input wire gpio_in_pad,
	output wire gpio_outenb_pad,
	output wire gpio_inenb_pad,
	output wire gpio_mode0_pad,
	output wire gpio_mode1_pad,
	output reg [127:0] la_output,
	input wire [127:0] la_input,
	output reg [127:0] la_oenb,
	output reg [127:0] la_iena,
	output wire qspi_enabled,
	output wire spi_enabled,
	output wire trap,
	output wire [2:0] user_irq_ena,
	input wire [5:0] user_irq,

    input wire clk_in,
    output wire clk_out,
    input wire resetn_in,
    output wire resetn_out,
    input wire serial_load_in,
    output wire serial_load_out,
    input wire serial_data_2_in,
    output wire serial_data_2_out,
    input wire serial_resetn_in,
    output wire serial_resetn_out,
    input wire serial_clock_in,
    output wire serial_clock_out,
    input wire rstb_l_in,
    output wire rstb_l_out
	// [Vic]: POR here is useless
    //input wire por_l_in,
    //output wire por_l_out,
    //input wire porb_h_in,
    //output wire porb_h_out
);

wire core_rst;
wire sys_clk;
wire sys_rst;
wire por_clk;
reg int_rst;
reg mgmtsoc_soc_rst;
wire mgmtsoc_cpu_rst;
reg [1:0] mgmtsoc_reset_storage;
reg mgmtsoc_reset_re;
reg [31:0] mgmtsoc_scratch_storage;
reg mgmtsoc_scratch_re;
wire [31:0] mgmtsoc_bus_errors_status;
wire mgmtsoc_bus_errors_we;
reg mgmtsoc_bus_errors_re;
wire mgmtsoc_bus_error;
reg [31:0] mgmtsoc_bus_errors;
wire mgmtsoc_reset;
reg [31:0] mgmtsoc_interrupt;
wire [29:0] mgmtsoc_ibus_ibus_adr;
wire [31:0] mgmtsoc_ibus_ibus_dat_w;
wire [31:0] mgmtsoc_ibus_ibus_dat_r;
wire [3:0] mgmtsoc_ibus_ibus_sel;
wire mgmtsoc_ibus_ibus_cyc;
wire mgmtsoc_ibus_ibus_stb;
wire mgmtsoc_ibus_ibus_ack;
wire mgmtsoc_ibus_ibus_we;
wire [2:0] mgmtsoc_ibus_ibus_cti;
wire [1:0] mgmtsoc_ibus_ibus_bte;
wire mgmtsoc_ibus_ibus_err;
wire [29:0] mgmtsoc_dbus_dbus_adr;
wire [31:0] mgmtsoc_dbus_dbus_dat_w;
wire [31:0] mgmtsoc_dbus_dbus_dat_r;
wire [3:0] mgmtsoc_dbus_dbus_sel;
wire mgmtsoc_dbus_dbus_cyc;
wire mgmtsoc_dbus_dbus_stb;
wire mgmtsoc_dbus_dbus_ack;
wire mgmtsoc_dbus_dbus_we;
wire [2:0] mgmtsoc_dbus_dbus_cti;
wire [1:0] mgmtsoc_dbus_dbus_bte;
wire mgmtsoc_dbus_dbus_err;
reg mgmtsoc_vexriscv_debug_reset;
reg mgmtsoc_vexriscv_ibus_err;
reg mgmtsoc_vexriscv_dbus_err;
reg mgmtsoc_vexriscv_i_cmd_valid;
reg mgmtsoc_vexriscv_i_cmd_payload_wr;
reg [7:0] mgmtsoc_vexriscv_i_cmd_payload_address;
reg [31:0] mgmtsoc_vexriscv_i_cmd_payload_data;
wire mgmtsoc_vexriscv_o_cmd_ready;
wire [31:0] mgmtsoc_vexriscv_o_rsp_data;
wire mgmtsoc_vexriscv_o_resetOut;
reg mgmtsoc_vexriscv_reset_debug_logic;
reg mgmtsoc_vexriscv_transfer_complete;
reg mgmtsoc_vexriscv_transfer_in_progress;
reg mgmtsoc_vexriscv_transfer_wait_for_ack;
wire [29:0] mgmtsoc_vexriscv_debug_bus_adr;
wire [31:0] mgmtsoc_vexriscv_debug_bus_dat_w;
reg [31:0] mgmtsoc_vexriscv_debug_bus_dat_r;
wire [3:0] mgmtsoc_vexriscv_debug_bus_sel;
wire mgmtsoc_vexriscv_debug_bus_cyc;
wire mgmtsoc_vexriscv_debug_bus_stb;
reg mgmtsoc_vexriscv_debug_bus_ack;
wire mgmtsoc_vexriscv_debug_bus_we;
wire [2:0] mgmtsoc_vexriscv_debug_bus_cti;
wire [1:0] mgmtsoc_vexriscv_debug_bus_bte;
wire mgmtsoc_vexriscv_debug_bus_err = 1'd0;
wire [31:0] mgmtsoc_vexriscv = 32'd268435456;
reg [31:0] mgmtsoc_load_storage;
reg mgmtsoc_load_re;
reg [31:0] mgmtsoc_reload_storage;
reg mgmtsoc_reload_re;
reg mgmtsoc_en_storage;
reg mgmtsoc_en_re;
reg mgmtsoc_update_value_storage;
reg mgmtsoc_update_value_re;
reg [31:0] mgmtsoc_value_status;
wire mgmtsoc_value_we;
reg mgmtsoc_value_re;
wire mgmtsoc_irq;
wire mgmtsoc_zero_status;
reg mgmtsoc_zero_pending;
wire mgmtsoc_zero_trigger;
reg mgmtsoc_zero_clear;
reg mgmtsoc_zero_trigger_d;
wire mgmtsoc_zero0;
wire mgmtsoc_status_status;
wire mgmtsoc_status_we;
reg mgmtsoc_status_re;
wire mgmtsoc_zero1;
wire mgmtsoc_pending_status;
wire mgmtsoc_pending_we;
reg mgmtsoc_pending_re;
reg mgmtsoc_pending_r;
wire mgmtsoc_zero2;
reg mgmtsoc_enable_storage;
reg mgmtsoc_enable_re;
reg [31:0] mgmtsoc_value;
wire [29:0] dff_bus_adr;
wire [31:0] dff_bus_dat_w;
wire [31:0] dff_bus_dat_r;
wire [3:0] dff_bus_sel;
wire dff_bus_cyc;
wire dff_bus_stb;
reg dff_bus_ack;
wire dff_bus_we;
wire [2:0] dff_bus_cti;
wire [1:0] dff_bus_bte;
wire dff_bus_err = 1'd0;
wire [31:0] dff_di;
wire [31:0] dff_do;
reg [3:0] dff_we;
wire dff_en;
wire [29:0] dff2_bus_adr;
wire [31:0] dff2_bus_dat_w;
wire [31:0] dff2_bus_dat_r;
wire [3:0] dff2_bus_sel;
wire dff2_bus_cyc;
wire dff2_bus_stb;
reg dff2_bus_ack;
wire dff2_bus_we;
wire [2:0] dff2_bus_cti;
wire [1:0] dff2_bus_bte;
wire dff2_bus_err = 1'd0;
wire [31:0] dff2_di;
wire [31:0] dff2_do;
reg [3:0] dff2_we;
wire dff2_en;
reg mgmtsoc_litespisdrphycore_source_valid;
wire mgmtsoc_litespisdrphycore_source_ready;
wire mgmtsoc_litespisdrphycore_source_first = 1'd0;
reg mgmtsoc_litespisdrphycore_source_last;
wire [31:0] mgmtsoc_litespisdrphycore_source_payload_data;
wire mgmtsoc_litespisdrphycore_sink_valid;
reg mgmtsoc_litespisdrphycore_sink_ready;
wire mgmtsoc_litespisdrphycore_sink_first;
wire mgmtsoc_litespisdrphycore_sink_last;
wire [31:0] mgmtsoc_litespisdrphycore_sink_payload_data;
wire [5:0] mgmtsoc_litespisdrphycore_sink_payload_len;
wire [3:0] mgmtsoc_litespisdrphycore_sink_payload_width;
wire [7:0] mgmtsoc_litespisdrphycore_sink_payload_mask;
wire mgmtsoc_litespisdrphycore_cs;
wire [7:0] mgmtsoc_litespisdrphycore_spi_clk_divisor;
reg [7:0] mgmtsoc_litespisdrphycore_storage;
reg mgmtsoc_litespisdrphycore_re;
wire [7:0] mgmtsoc_litespisdrphycore_div;
wire [7:0] mgmtsoc_litespisdrphycore_sample_cnt;
wire [7:0] mgmtsoc_litespisdrphycore_update_cnt;
wire mgmtsoc_litespisdrphycore_posedge;
wire mgmtsoc_litespisdrphycore_negedge;
wire mgmtsoc_litespisdrphycore_sample;
wire mgmtsoc_litespisdrphycore_update;
reg mgmtsoc_litespisdrphycore_en;
reg [7:0] mgmtsoc_litespisdrphycore_cnt;
wire mgmtsoc_litespisdrphycore_en_int = 1'd0;
reg mgmtsoc_litespisdrphycore_clk;
reg mgmtsoc_litespisdrphycore_posedge_reg;
reg mgmtsoc_litespisdrphycore_posedge_reg2;
wire mgmtsoc_litespisdrphycore_wait;
wire mgmtsoc_litespisdrphycore_done;
reg [3:0] mgmtsoc_litespisdrphycore_count;
wire mgmtsoc_litespisdrphycore_cs_enable;
reg mgmtsoc_litespisdrphycore_dq_o;
reg [1:0] mgmtsoc_litespisdrphycore_dq_i;
wire mgmtsoc_litespisdrphycore_dq_oe;
reg [7:0] mgmtsoc_litespisdrphycore_sr_cnt;
reg mgmtsoc_litespisdrphycore_sr_out_load;
reg mgmtsoc_litespisdrphycore_sr_out_shift;
reg [31:0] mgmtsoc_litespisdrphycore_sr_out;
reg mgmtsoc_litespisdrphycore_sr_in_shift;
reg [31:0] mgmtsoc_litespisdrphycore_sr_in;
wire mgmtsoc_litespisdrphycore0 = 1'd0;
wire [1:0] mgmtsoc_litespisdrphycore1 = 2'd0;
wire [3:0] mgmtsoc_litespisdrphycore2 = 4'd0;
wire [7:0] mgmtsoc_litespisdrphycore3 = 8'd0;
wire mgmtsoc_crossbar_source_valid;
wire mgmtsoc_crossbar_source_ready;
wire mgmtsoc_crossbar_source_first;
wire mgmtsoc_crossbar_source_last;
wire [31:0] mgmtsoc_crossbar_source_payload_data;
wire [5:0] mgmtsoc_crossbar_source_payload_len;
wire [3:0] mgmtsoc_crossbar_source_payload_width;
wire [7:0] mgmtsoc_crossbar_source_payload_mask;
wire mgmtsoc_crossbar_sink_valid;
wire mgmtsoc_crossbar_sink_ready;
wire mgmtsoc_crossbar_sink_first;
wire mgmtsoc_crossbar_sink_last;
wire [31:0] mgmtsoc_crossbar_sink_payload_data;
reg mgmtsoc_crossbar_cs;
reg mgmtsoc_litespimmap_source_valid;
wire mgmtsoc_litespimmap_source_ready;
wire mgmtsoc_litespimmap_source_first = 1'd0;
reg mgmtsoc_litespimmap_source_last;
reg [31:0] mgmtsoc_litespimmap_source_payload_data;
reg [5:0] mgmtsoc_litespimmap_source_payload_len;
reg [3:0] mgmtsoc_litespimmap_source_payload_width;
reg [7:0] mgmtsoc_litespimmap_source_payload_mask;
wire mgmtsoc_litespimmap_sink_valid;
reg mgmtsoc_litespimmap_sink_ready;
wire mgmtsoc_litespimmap_sink_first;
wire mgmtsoc_litespimmap_sink_last;
wire [31:0] mgmtsoc_litespimmap_sink_payload_data;
wire [29:0] mgmtsoc_litespimmap_bus_adr;
wire [31:0] mgmtsoc_litespimmap_bus_dat_w;
reg [31:0] mgmtsoc_litespimmap_bus_dat_r;
wire [3:0] mgmtsoc_litespimmap_bus_sel;
wire mgmtsoc_litespimmap_bus_cyc;
wire mgmtsoc_litespimmap_bus_stb;
reg mgmtsoc_litespimmap_bus_ack;
wire mgmtsoc_litespimmap_bus_we;
wire [2:0] mgmtsoc_litespimmap_bus_cti;
wire [1:0] mgmtsoc_litespimmap_bus_bte;
wire mgmtsoc_litespimmap_bus_err = 1'd0;
reg mgmtsoc_litespimmap_cs;
reg mgmtsoc_litespimmap_burst_cs;
reg [29:0] mgmtsoc_litespimmap_burst_adr;
reg mgmtsoc_litespimmap_wait;
wire mgmtsoc_litespimmap_done;
reg [8:0] mgmtsoc_litespimmap_count;
reg [7:0] mgmtsoc_litespimmap_storage;
reg mgmtsoc_litespimmap_re;
wire [7:0] mgmtsoc_litespimmap_spi_dummy_bits;
wire [31:0] mgmtsoc_litespimmap_dummy = 32'd57005;
wire [1:0] mgmtsoc_litespimmap = 2'd0;
wire mgmtsoc_port_mmap_user_port_source_valid;
wire mgmtsoc_port_mmap_user_port_source_ready;
wire mgmtsoc_port_mmap_user_port_source_first;
wire mgmtsoc_port_mmap_user_port_source_last;
wire [31:0] mgmtsoc_port_mmap_user_port_source_payload_data;
wire mgmtsoc_port_mmap_user_port_sink_valid;
wire mgmtsoc_port_mmap_user_port_sink_ready;
wire mgmtsoc_port_mmap_user_port_sink_first;
wire mgmtsoc_port_mmap_user_port_sink_last;
wire [31:0] mgmtsoc_port_mmap_user_port_sink_payload_data;
wire [5:0] mgmtsoc_port_mmap_user_port_sink_payload_len;
wire [3:0] mgmtsoc_port_mmap_user_port_sink_payload_width;
wire [7:0] mgmtsoc_port_mmap_user_port_sink_payload_mask;
wire mgmtsoc_port_mmap_internal_port_source_valid;
wire mgmtsoc_port_mmap_internal_port_source_ready;
wire mgmtsoc_port_mmap_internal_port_source_first;
wire mgmtsoc_port_mmap_internal_port_source_last;
wire [31:0] mgmtsoc_port_mmap_internal_port_source_payload_data;
wire mgmtsoc_port_mmap_internal_port_sink_valid;
wire mgmtsoc_port_mmap_internal_port_sink_ready;
wire mgmtsoc_port_mmap_internal_port_sink_first;
wire mgmtsoc_port_mmap_internal_port_sink_last;
wire [31:0] mgmtsoc_port_mmap_internal_port_sink_payload_data;
wire [5:0] mgmtsoc_port_mmap_internal_port_sink_payload_len;
wire [3:0] mgmtsoc_port_mmap_internal_port_sink_payload_width;
wire [7:0] mgmtsoc_port_mmap_internal_port_sink_payload_mask;
wire mgmtsoc_port_mmap_request;
wire mgmtsoc_master_sink_sink_valid;
wire mgmtsoc_master_sink_sink_ready;
wire mgmtsoc_master_sink_sink_first;
wire mgmtsoc_master_sink_sink_last;
wire [31:0] mgmtsoc_master_sink_sink_payload_data;
wire mgmtsoc_master_source_source_valid;
wire mgmtsoc_master_source_source_ready;
wire mgmtsoc_master_source_source_first;
wire mgmtsoc_master_source_source_last;
wire [31:0] mgmtsoc_master_source_source_payload_data;
wire [5:0] mgmtsoc_master_source_source_payload_len;
wire [3:0] mgmtsoc_master_source_source_payload_width;
wire [7:0] mgmtsoc_master_source_source_payload_mask;
wire mgmtsoc_master_cs;
reg mgmtsoc_master_cs_storage;
reg mgmtsoc_master_cs_re;
wire [7:0] mgmtsoc_master_len;
wire [3:0] mgmtsoc_master_width;
wire [7:0] mgmtsoc_master_mask;
reg [23:0] mgmtsoc_master_phyconfig_storage;
reg mgmtsoc_master_phyconfig_re;
reg mgmtsoc_master_rxtx_re;
wire [31:0] mgmtsoc_master_rxtx_r;
reg mgmtsoc_master_rxtx_we;
wire [31:0] mgmtsoc_master_rxtx_w;
wire mgmtsoc_master_tx_ready;
wire mgmtsoc_master_rx_ready;
reg [1:0] mgmtsoc_master_status_status;
wire mgmtsoc_master_status_we;
reg mgmtsoc_master_status_re;
wire mgmtsoc_master_tx_fifo_sink_valid;
wire mgmtsoc_master_tx_fifo_sink_ready;
wire mgmtsoc_master_tx_fifo_sink_first = 1'd0;
wire mgmtsoc_master_tx_fifo_sink_last;
wire [31:0] mgmtsoc_master_tx_fifo_sink_payload_data;
wire [5:0] mgmtsoc_master_tx_fifo_sink_payload_len;
wire [3:0] mgmtsoc_master_tx_fifo_sink_payload_width;
wire [7:0] mgmtsoc_master_tx_fifo_sink_payload_mask;
reg mgmtsoc_master_tx_fifo_source_valid;
wire mgmtsoc_master_tx_fifo_source_ready;
reg mgmtsoc_master_tx_fifo_source_first;
reg mgmtsoc_master_tx_fifo_source_last;
reg [31:0] mgmtsoc_master_tx_fifo_source_payload_data;
reg [5:0] mgmtsoc_master_tx_fifo_source_payload_len;
reg [3:0] mgmtsoc_master_tx_fifo_source_payload_width;
reg [7:0] mgmtsoc_master_tx_fifo_source_payload_mask;
wire mgmtsoc_master_rx_fifo_sink_valid;
wire mgmtsoc_master_rx_fifo_sink_ready;
wire mgmtsoc_master_rx_fifo_sink_first;
wire mgmtsoc_master_rx_fifo_sink_last;
wire [31:0] mgmtsoc_master_rx_fifo_sink_payload_data;
reg mgmtsoc_master_rx_fifo_source_valid;
wire mgmtsoc_master_rx_fifo_source_ready;
reg mgmtsoc_master_rx_fifo_source_first;
reg mgmtsoc_master_rx_fifo_source_last;
reg [31:0] mgmtsoc_master_rx_fifo_source_payload_data;
wire mgmtsoc_port_master_user_port_source_valid;
wire mgmtsoc_port_master_user_port_source_ready;
wire mgmtsoc_port_master_user_port_source_first;
wire mgmtsoc_port_master_user_port_source_last;
wire [31:0] mgmtsoc_port_master_user_port_source_payload_data;
wire mgmtsoc_port_master_user_port_sink_valid;
wire mgmtsoc_port_master_user_port_sink_ready;
wire mgmtsoc_port_master_user_port_sink_first;
wire mgmtsoc_port_master_user_port_sink_last;
wire [31:0] mgmtsoc_port_master_user_port_sink_payload_data;
wire [5:0] mgmtsoc_port_master_user_port_sink_payload_len;
wire [3:0] mgmtsoc_port_master_user_port_sink_payload_width;
wire [7:0] mgmtsoc_port_master_user_port_sink_payload_mask;
wire mgmtsoc_port_master_internal_port_source_valid;
wire mgmtsoc_port_master_internal_port_source_ready;
wire mgmtsoc_port_master_internal_port_source_first;
wire mgmtsoc_port_master_internal_port_source_last;
wire [31:0] mgmtsoc_port_master_internal_port_source_payload_data;
wire mgmtsoc_port_master_internal_port_sink_valid;
wire mgmtsoc_port_master_internal_port_sink_ready;
wire mgmtsoc_port_master_internal_port_sink_first;
wire mgmtsoc_port_master_internal_port_sink_last;
wire [31:0] mgmtsoc_port_master_internal_port_sink_payload_data;
wire [5:0] mgmtsoc_port_master_internal_port_sink_payload_len;
wire [3:0] mgmtsoc_port_master_internal_port_sink_payload_width;
wire [7:0] mgmtsoc_port_master_internal_port_sink_payload_mask;
wire mgmtsoc_port_master_request;
wire spi_master_start0;
wire [7:0] spi_master_length0;
reg spi_master_done0;
reg spi_master_irq;
wire [7:0] spi_master_mosi;
reg [7:0] spi_master_miso;
wire spi_master_cs;
wire spi_master_cs_mode;
wire spi_master_loopback;
wire [15:0] spi_master_clk_divider0;
reg spi_master_start1;
wire [7:0] spi_master_length1;
reg [15:0] spi_master_control_storage;
reg spi_master_control_re;
wire spi_master_done1;
wire spi_master_status_status;
wire spi_master_status_we;
reg spi_master_status_re;
reg [7:0] spi_master_mosi_storage;
reg spi_master_mosi_re;
wire [7:0] spi_master_miso_status;
wire spi_master_miso_we;
reg spi_master_miso_re;
wire spi_master_sel;
wire spi_master_mode0;
reg [16:0] spi_master_cs_storage;
reg spi_master_cs_re;
wire spi_master_mode1;
reg spi_master_loopback_storage;
reg spi_master_loopback_re;
reg spi_master_clk_enable;
reg spi_master_xfer_enable;
reg [2:0] spi_master_count;
reg spi_master_mosi_latch;
reg spi_master_miso_latch;
reg [15:0] spi_master_clk_divider1;
wire spi_master_clk_rise;
wire spi_master_clk_fall;
reg [7:0] spi_master_mosi_data;
reg [2:0] spi_master_mosi_sel;
reg [7:0] spi_master_miso_data;
reg [15:0] spimaster_storage;
reg spimaster_re;
wire [29:0] mprj_adr;
wire [31:0] mprj_dat_w;
wire [31:0] mprj_dat_r;
wire [3:0] mprj_sel;
wire mprj_cyc;
wire mprj_stb;
wire mprj_ack;
wire mprj_we;
wire [2:0] mprj_cti;
wire [1:0] mprj_bte;
wire mprj_err = 1'd0;
reg mprj_wb_iena_storage;
reg mprj_wb_iena_re;
wire [29:0] hk_adr;
wire [31:0] hk_dat_w;
wire [31:0] hk_dat_r;
wire [3:0] hk_sel;
wire hk_cyc;
wire hk_stb;
wire hk_ack;
wire hk_we;
wire [2:0] hk_cti;
wire [1:0] hk_bte;
wire hk_err = 1'd0;
reg sys_uart_rx;
reg sys_uart_tx;
wire uart_phy_tx_sink_valid;
reg uart_phy_tx_sink_ready;
wire uart_phy_tx_sink_first;
wire uart_phy_tx_sink_last;
wire [7:0] uart_phy_tx_sink_payload_data;
reg [7:0] uart_phy_tx_data;
reg [3:0] uart_phy_tx_count;
reg uart_phy_tx_enable;
reg uart_phy_tx_tick;
reg [31:0] uart_phy_tx_phase;
reg uart_phy_rx_source_valid;
wire uart_phy_rx_source_ready;
wire uart_phy_rx_source_first = 1'd0;
wire uart_phy_rx_source_last = 1'd0;
reg [7:0] uart_phy_rx_source_payload_data;
reg [7:0] uart_phy_rx_data;
reg [3:0] uart_phy_rx_count;
reg uart_phy_rx_enable;
reg uart_phy_rx_tick;
reg [31:0] uart_phy_rx_phase;
wire uart_phy_rx_rx;
reg uart_phy_rx_rx_d;
reg uart_rxtx_re;
wire [7:0] uart_rxtx_r;
reg uart_rxtx_we;
wire [7:0] uart_rxtx_w;
wire uart_txfull_status;
wire uart_txfull_we;
reg uart_txfull_re;
wire uart_rxempty_status;
wire uart_rxempty_we;
reg uart_rxempty_re;
wire uart_irq;
wire uart_tx_status;
reg uart_tx_pending;
wire uart_tx_trigger;
reg uart_tx_clear;
reg uart_tx_trigger_d;
wire uart_rx_status;
reg uart_rx_pending;
wire uart_rx_trigger;
reg uart_rx_clear;
reg uart_rx_trigger_d;
wire uart_tx0;
wire uart_rx0;
reg [1:0] uart_status_status;
wire uart_status_we;
reg uart_status_re;
wire uart_tx1;
wire uart_rx1;
reg [1:0] uart_pending_status;
wire uart_pending_we;
reg uart_pending_re;
reg [1:0] uart_pending_r;
wire uart_tx2;
wire uart_rx2;
reg [1:0] uart_enable_storage;
reg uart_enable_re;
wire uart_txempty_status;
wire uart_txempty_we;
reg uart_txempty_re;
wire uart_rxfull_status;
wire uart_rxfull_we;
reg uart_rxfull_re;
wire uart_uart_sink_valid;
wire uart_uart_sink_ready;
wire uart_uart_sink_first;
wire uart_uart_sink_last;
wire [7:0] uart_uart_sink_payload_data;
wire uart_uart_source_valid;
wire uart_uart_source_ready;
wire uart_uart_source_first;
wire uart_uart_source_last;
wire [7:0] uart_uart_source_payload_data;
wire uart_tx_fifo_sink_valid;
wire uart_tx_fifo_sink_ready;
wire uart_tx_fifo_sink_first = 1'd0;
wire uart_tx_fifo_sink_last = 1'd0;
wire [7:0] uart_tx_fifo_sink_payload_data;
wire uart_tx_fifo_source_valid;
wire uart_tx_fifo_source_ready;
wire uart_tx_fifo_source_first;
wire uart_tx_fifo_source_last;
wire [7:0] uart_tx_fifo_source_payload_data;
wire uart_tx_fifo_re;
reg uart_tx_fifo_readable;
wire uart_tx_fifo_syncfifo_we;
wire uart_tx_fifo_syncfifo_writable;
wire uart_tx_fifo_syncfifo_re;
wire uart_tx_fifo_syncfifo_readable;
wire [9:0] uart_tx_fifo_syncfifo_din;
wire [9:0] uart_tx_fifo_syncfifo_dout;
reg [4:0] uart_tx_fifo_level0;
wire uart_tx_fifo_replace = 1'd0;
reg [3:0] uart_tx_fifo_produce;
reg [3:0] uart_tx_fifo_consume;
reg [3:0] uart_tx_fifo_wrport_adr;
wire [9:0] uart_tx_fifo_wrport_dat_r;
wire uart_tx_fifo_wrport_we;
wire [9:0] uart_tx_fifo_wrport_dat_w;
wire uart_tx_fifo_do_read;
wire [3:0] uart_tx_fifo_rdport_adr;
wire [9:0] uart_tx_fifo_rdport_dat_r;
wire uart_tx_fifo_rdport_re;
wire [4:0] uart_tx_fifo_level1;
wire [7:0] uart_tx_fifo_fifo_in_payload_data;
wire uart_tx_fifo_fifo_in_first;
wire uart_tx_fifo_fifo_in_last;
wire [7:0] uart_tx_fifo_fifo_out_payload_data;
wire uart_tx_fifo_fifo_out_first;
wire uart_tx_fifo_fifo_out_last;
wire uart_rx_fifo_sink_valid;
wire uart_rx_fifo_sink_ready;
wire uart_rx_fifo_sink_first;
wire uart_rx_fifo_sink_last;
wire [7:0] uart_rx_fifo_sink_payload_data;
wire uart_rx_fifo_source_valid;
wire uart_rx_fifo_source_ready;
wire uart_rx_fifo_source_first;
wire uart_rx_fifo_source_last;
wire [7:0] uart_rx_fifo_source_payload_data;
wire uart_rx_fifo_re;
reg uart_rx_fifo_readable;
wire uart_rx_fifo_syncfifo_we;
wire uart_rx_fifo_syncfifo_writable;
wire uart_rx_fifo_syncfifo_re;
wire uart_rx_fifo_syncfifo_readable;
wire [9:0] uart_rx_fifo_syncfifo_din;
wire [9:0] uart_rx_fifo_syncfifo_dout;
reg [4:0] uart_rx_fifo_level0;
wire uart_rx_fifo_replace = 1'd0;
reg [3:0] uart_rx_fifo_produce;
reg [3:0] uart_rx_fifo_consume;
reg [3:0] uart_rx_fifo_wrport_adr;
wire [9:0] uart_rx_fifo_wrport_dat_r;
wire uart_rx_fifo_wrport_we;
wire [9:0] uart_rx_fifo_wrport_dat_w;
wire uart_rx_fifo_do_read;
wire [3:0] uart_rx_fifo_rdport_adr;
wire [9:0] uart_rx_fifo_rdport_dat_r;
wire uart_rx_fifo_rdport_re;
wire [4:0] uart_rx_fifo_level1;
wire [7:0] uart_rx_fifo_fifo_in_payload_data;
wire uart_rx_fifo_fifo_in_first;
wire uart_rx_fifo_fifo_in_last;
wire [7:0] uart_rx_fifo_fifo_out_payload_data;
wire uart_rx_fifo_fifo_out_first;
wire uart_rx_fifo_fifo_out_last;
reg dbg_uart_dbg_uart_rx;
reg dbg_uart_dbg_uart_tx;
reg dbg_uart_tx_sink_valid;
reg dbg_uart_tx_sink_ready;
wire dbg_uart_tx_sink_last;
reg [7:0] dbg_uart_tx_sink_payload_data;
reg [7:0] dbg_uart_tx_data;
reg [3:0] dbg_uart_tx_count;
reg dbg_uart_tx_enable;
reg dbg_uart_tx_tick;
reg [31:0] dbg_uart_tx_phase;
reg dbg_uart_rx_source_valid;
reg dbg_uart_rx_source_ready;
reg [7:0] dbg_uart_rx_source_payload_data;
reg [7:0] dbg_uart_rx_data;
reg [3:0] dbg_uart_rx_count;
reg dbg_uart_rx_enable;
reg dbg_uart_rx_tick;
reg [31:0] dbg_uart_rx_phase;
wire dbg_uart_rx_rx;
reg dbg_uart_rx_rx_d;
wire [29:0] dbg_uart_wishbone_adr;
wire [31:0] dbg_uart_wishbone_dat_w;
wire [31:0] dbg_uart_wishbone_dat_r;
wire [3:0] dbg_uart_wishbone_sel;
reg dbg_uart_wishbone_cyc;
reg dbg_uart_wishbone_stb;
wire dbg_uart_wishbone_ack;
reg dbg_uart_wishbone_we;
wire [2:0] dbg_uart_wishbone_cti = 3'd0;
wire [1:0] dbg_uart_wishbone_bte = 2'd0;
wire dbg_uart_wishbone_err;
reg [7:0] dbg_uart_cmd;
reg dbg_uart_incr;
reg [7:0] dbg_uart_length;
reg [31:0] dbg_uart_address;
reg [31:0] dbg_uart_data;
reg [1:0] dbg_uart_bytes_count;
reg [7:0] dbg_uart_words_count;
wire dbg_uart_reset;
wire dbg_uart_wait;
wire dbg_uart_done;
reg [19:0] dbg_uart_count;
reg dbg_uart_is_ongoing;
reg debug_oeb_storage;
reg debug_oeb_re;
reg debug_mode_storage;
reg debug_mode_re;
wire uart_enabled_o;
reg uart_enabled_storage;
reg uart_enabled_re;
reg gpio_mode1_storage;
reg gpio_mode1_re;
reg gpio_mode0_storage;
reg gpio_mode0_re;
reg gpio_ien_storage;
reg gpio_ien_re;
reg gpio_oe_storage;
reg gpio_oe_re;
wire gpio_in_status;
wire gpio_in_we;
reg gpio_in_re;
reg gpio_out_storage;
reg gpio_out_re;
reg [127:0] la_ien_storage;
reg la_ien_re;
reg [127:0] la_oe_storage;
reg la_oe_re;
reg [127:0] la_in_status;
wire la_in_we;
reg la_in_re;
reg [127:0] la_out_storage;
reg la_out_re;
reg spi_enabled_storage;
reg spi_enabled_re;
reg [2:0] user_irq_ena_storage;
reg user_irq_ena_re;
wire gpioin0_in_status;
wire gpioin0_in_we;
reg gpioin0_in_re;
reg gpioin0_gpioin0_mode_storage;
reg gpioin0_gpioin0_mode_re;
reg gpioin0_gpioin0_edge_storage;
reg gpioin0_gpioin0_edge_re;
wire gpioin0_gpioin0_irq;
reg gpioin0_gpioin0_in_pads_n_d;
wire gpioin0_gpioin0_status;
reg gpioin0_gpioin0_pending;
reg gpioin0_gpioin0_trigger;
reg gpioin0_gpioin0_clear;
reg gpioin0_gpioin0_trigger_d;
wire gpioin1_in_status;
wire gpioin1_in_we;
reg gpioin1_in_re;
reg gpioin1_gpioin1_mode_storage;
reg gpioin1_gpioin1_mode_re;
reg gpioin1_gpioin1_edge_storage;
reg gpioin1_gpioin1_edge_re;
wire gpioin1_gpioin1_irq;
reg gpioin1_gpioin1_in_pads_n_d;
wire gpioin1_gpioin1_status;
reg gpioin1_gpioin1_pending;
reg gpioin1_gpioin1_trigger;
reg gpioin1_gpioin1_clear;
reg gpioin1_gpioin1_trigger_d;
wire gpioin2_in_status;
wire gpioin2_in_we;
reg gpioin2_in_re;
reg gpioin2_gpioin2_mode_storage;
reg gpioin2_gpioin2_mode_re;
reg gpioin2_gpioin2_edge_storage;
reg gpioin2_gpioin2_edge_re;
wire gpioin2_gpioin2_irq;
reg gpioin2_gpioin2_in_pads_n_d;
wire gpioin2_gpioin2_status;
reg gpioin2_gpioin2_pending;
reg gpioin2_gpioin2_trigger;
reg gpioin2_gpioin2_clear;
reg gpioin2_gpioin2_trigger_d;
wire gpioin3_in_status;
wire gpioin3_in_we;
reg gpioin3_in_re;
reg gpioin3_gpioin3_mode_storage;
reg gpioin3_gpioin3_mode_re;
reg gpioin3_gpioin3_edge_storage;
reg gpioin3_gpioin3_edge_re;
wire gpioin3_gpioin3_irq;
reg gpioin3_gpioin3_in_pads_n_d;
wire gpioin3_gpioin3_status;
reg gpioin3_gpioin3_pending;
reg gpioin3_gpioin3_trigger;
reg gpioin3_gpioin3_clear;
reg gpioin3_gpioin3_trigger_d;
wire gpioin4_in_status;
wire gpioin4_in_we;
reg gpioin4_in_re;
reg gpioin4_gpioin4_mode_storage;
reg gpioin4_gpioin4_mode_re;
reg gpioin4_gpioin4_edge_storage;
reg gpioin4_gpioin4_edge_re;
wire gpioin4_gpioin4_irq;
reg gpioin4_gpioin4_in_pads_n_d;
wire gpioin4_gpioin4_status;
reg gpioin4_gpioin4_pending;
reg gpioin4_gpioin4_trigger;
reg gpioin4_gpioin4_clear;
reg gpioin4_gpioin4_trigger_d;
wire gpioin5_in_status;
wire gpioin5_in_we;
reg gpioin5_in_re;
reg gpioin5_gpioin5_mode_storage;
reg gpioin5_gpioin5_mode_re;
reg gpioin5_gpioin5_edge_storage;
reg gpioin5_gpioin5_edge_re;
wire gpioin5_gpioin5_irq;
reg gpioin5_gpioin5_in_pads_n_d;
wire gpioin5_gpioin5_status;
reg gpioin5_gpioin5_pending;
reg gpioin5_gpioin5_trigger;
reg gpioin5_gpioin5_clear;
reg gpioin5_gpioin5_trigger_d;
reg [1:0] litespiphy_state;
reg [1:0] litespiphy_next_state;
reg [7:0] mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value;
reg mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value_ce;
wire [1:0] litespi_request;
reg litespi_grant;
reg litespi_tx_mux_source_valid;
wire litespi_tx_mux_source_ready;
reg litespi_tx_mux_source_first;
reg litespi_tx_mux_source_last;
reg [31:0] litespi_tx_mux_source_payload_data;
reg [5:0] litespi_tx_mux_source_payload_len;
reg [3:0] litespi_tx_mux_source_payload_width;
reg [7:0] litespi_tx_mux_source_payload_mask;
wire litespi_tx_mux_endpoint0_sink_valid;
reg litespi_tx_mux_endpoint0_sink_ready;
wire litespi_tx_mux_endpoint0_sink_first;
wire litespi_tx_mux_endpoint0_sink_last;
wire [31:0] litespi_tx_mux_endpoint0_sink_payload_data;
wire [5:0] litespi_tx_mux_endpoint0_sink_payload_len;
wire [3:0] litespi_tx_mux_endpoint0_sink_payload_width;
wire [7:0] litespi_tx_mux_endpoint0_sink_payload_mask;
wire litespi_tx_mux_endpoint1_sink_valid;
reg litespi_tx_mux_endpoint1_sink_ready;
wire litespi_tx_mux_endpoint1_sink_first;
wire litespi_tx_mux_endpoint1_sink_last;
wire [31:0] litespi_tx_mux_endpoint1_sink_payload_data;
wire [5:0] litespi_tx_mux_endpoint1_sink_payload_len;
wire [3:0] litespi_tx_mux_endpoint1_sink_payload_width;
wire [7:0] litespi_tx_mux_endpoint1_sink_payload_mask;
wire litespi_tx_mux_sel;
wire litespi_rx_demux_sink_valid;
reg litespi_rx_demux_sink_ready;
wire litespi_rx_demux_sink_first;
wire litespi_rx_demux_sink_last;
wire [31:0] litespi_rx_demux_sink_payload_data;
reg litespi_rx_demux_endpoint0_source_valid;
wire litespi_rx_demux_endpoint0_source_ready;
reg litespi_rx_demux_endpoint0_source_first;
reg litespi_rx_demux_endpoint0_source_last;
reg [31:0] litespi_rx_demux_endpoint0_source_payload_data;
reg litespi_rx_demux_endpoint1_source_valid;
wire litespi_rx_demux_endpoint1_source_ready;
reg litespi_rx_demux_endpoint1_source_first;
reg litespi_rx_demux_endpoint1_source_last;
reg [31:0] litespi_rx_demux_endpoint1_source_payload_data;
wire litespi_rx_demux_sel;
reg [3:0] litespi_state;
reg [3:0] litespi_next_state;
reg mgmtsoc_litespimmap_burst_cs_litespi_next_value0;
reg mgmtsoc_litespimmap_burst_cs_litespi_next_value_ce0;
reg [29:0] mgmtsoc_litespimmap_burst_adr_litespi_next_value1;
reg mgmtsoc_litespimmap_burst_adr_litespi_next_value_ce1;
reg [1:0] spimaster_state;
reg [1:0] spimaster_next_state;
reg [2:0] spi_master_count_spimaster_next_value;
reg spi_master_count_spimaster_next_value_ce;
reg rs232phy_rs232phytx_state;
reg rs232phy_rs232phytx_next_state;
reg [3:0] uart_phy_tx_count_rs232phy_rs232phytx_next_value0;
reg uart_phy_tx_count_rs232phy_rs232phytx_next_value_ce0;
reg sys_uart_tx_rs232phy_rs232phytx_next_value1;
reg sys_uart_tx_rs232phy_rs232phytx_next_value_ce1;
reg [7:0] uart_phy_tx_data_rs232phy_rs232phytx_next_value2;
reg uart_phy_tx_data_rs232phy_rs232phytx_next_value_ce2;
reg rs232phy_rs232phyrx_state;
reg rs232phy_rs232phyrx_next_state;
reg [3:0] uart_phy_rx_count_rs232phy_rs232phyrx_next_value0;
reg uart_phy_rx_count_rs232phy_rs232phyrx_next_value_ce0;
reg [7:0] uart_phy_rx_data_rs232phy_rs232phyrx_next_value1;
reg uart_phy_rx_data_rs232phy_rs232phyrx_next_value_ce1;
reg uartwishbonebridge_rs232phytx_state;
reg uartwishbonebridge_rs232phytx_next_state;
reg [3:0] dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value0;
reg dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value_ce0;
reg dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value1;
reg dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value_ce1;
reg [7:0] dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value2;
reg dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value_ce2;
reg uartwishbonebridge_rs232phyrx_state;
reg uartwishbonebridge_rs232phyrx_next_state;
reg [3:0] dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value0;
reg dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value_ce0;
reg [7:0] dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value1;
reg dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value_ce1;
reg [2:0] uartwishbonebridge_state;
reg [2:0] uartwishbonebridge_next_state;
reg [1:0] dbg_uart_bytes_count_uartwishbonebridge_next_value0;
reg dbg_uart_bytes_count_uartwishbonebridge_next_value_ce0;
reg [7:0] dbg_uart_words_count_uartwishbonebridge_next_value1;
reg dbg_uart_words_count_uartwishbonebridge_next_value_ce1;
reg [7:0] dbg_uart_cmd_uartwishbonebridge_next_value2;
reg dbg_uart_cmd_uartwishbonebridge_next_value_ce2;
reg [7:0] dbg_uart_length_uartwishbonebridge_next_value3;
reg dbg_uart_length_uartwishbonebridge_next_value_ce3;
reg [31:0] dbg_uart_address_uartwishbonebridge_next_value4;
reg dbg_uart_address_uartwishbonebridge_next_value_ce4;
reg dbg_uart_incr_uartwishbonebridge_next_value5;
reg dbg_uart_incr_uartwishbonebridge_next_value_ce5;
reg [31:0] dbg_uart_data_uartwishbonebridge_next_value6;
reg dbg_uart_data_uartwishbonebridge_next_value_ce6;
wire gpioin0_i00;
wire gpioin0_status_status;
wire gpioin0_status_we;
reg gpioin0_status_re;
wire gpioin0_i01;
wire gpioin0_pending_status;
wire gpioin0_pending_we;
reg gpioin0_pending_re;
reg gpioin0_pending_r;
wire gpioin0_i02;
reg gpioin0_enable_storage;
reg gpioin0_enable_re;
wire gpioin1_i00;
wire gpioin1_status_status;
wire gpioin1_status_we;
reg gpioin1_status_re;
wire gpioin1_i01;
wire gpioin1_pending_status;
wire gpioin1_pending_we;
reg gpioin1_pending_re;
reg gpioin1_pending_r;
wire gpioin1_i02;
reg gpioin1_enable_storage;
reg gpioin1_enable_re;
wire gpioin2_i00;
wire gpioin2_status_status;
wire gpioin2_status_we;
reg gpioin2_status_re;
wire gpioin2_i01;
wire gpioin2_pending_status;
wire gpioin2_pending_we;
reg gpioin2_pending_re;
reg gpioin2_pending_r;
wire gpioin2_i02;
reg gpioin2_enable_storage;
reg gpioin2_enable_re;
wire gpioin3_i00;
wire gpioin3_status_status;
wire gpioin3_status_we;
reg gpioin3_status_re;
wire gpioin3_i01;
wire gpioin3_pending_status;
wire gpioin3_pending_we;
reg gpioin3_pending_re;
reg gpioin3_pending_r;
wire gpioin3_i02;
reg gpioin3_enable_storage;
reg gpioin3_enable_re;
wire gpioin4_i00;
wire gpioin4_status_status;
wire gpioin4_status_we;
reg gpioin4_status_re;
wire gpioin4_i01;
wire gpioin4_pending_status;
wire gpioin4_pending_we;
reg gpioin4_pending_re;
reg gpioin4_pending_r;
wire gpioin4_i02;
reg gpioin4_enable_storage;
reg gpioin4_enable_re;
wire gpioin5_i00;
wire gpioin5_status_status;
wire gpioin5_status_we;
reg gpioin5_status_re;
wire gpioin5_i01;
wire gpioin5_pending_status;
wire gpioin5_pending_we;
reg gpioin5_pending_re;
reg gpioin5_pending_r;
wire gpioin5_i02;
reg gpioin5_enable_storage;
reg gpioin5_enable_re;
reg [13:0] mgmtsoc_adr;
reg mgmtsoc_we;
reg [31:0] mgmtsoc_dat_w;
wire [31:0] mgmtsoc_dat_r;
wire [29:0] mgmtsoc_wishbone_adr;
wire [31:0] mgmtsoc_wishbone_dat_w;
reg [31:0] mgmtsoc_wishbone_dat_r;
wire [3:0] mgmtsoc_wishbone_sel;
wire mgmtsoc_wishbone_cyc;
wire mgmtsoc_wishbone_stb;
reg mgmtsoc_wishbone_ack;
wire mgmtsoc_wishbone_we;
wire [2:0] mgmtsoc_wishbone_cti;
wire [1:0] mgmtsoc_wishbone_bte;
wire mgmtsoc_wishbone_err = 1'd0;
wire [29:0] shared_adr;
wire [31:0] shared_dat_w;
reg [31:0] shared_dat_r;
wire [3:0] shared_sel;
wire shared_cyc;
wire shared_stb;
reg shared_ack;
wire shared_we;
wire [2:0] shared_cti;
wire [1:0] shared_bte;
wire shared_err;
wire [2:0] request;
reg [1:0] grant;
reg [6:0] slave_sel;
reg [6:0] slave_sel_r;
reg error;
wire wait_1;
wire done;
reg [19:0] count;
wire [13:0] interface0_bank_bus_adr;
wire interface0_bank_bus_we;
wire [31:0] interface0_bank_bus_dat_w;
reg [31:0] interface0_bank_bus_dat_r;
reg csrbank0_reset0_re;
wire [1:0] csrbank0_reset0_r;
reg csrbank0_reset0_we;
wire [1:0] csrbank0_reset0_w;
reg csrbank0_scratch0_re;
wire [31:0] csrbank0_scratch0_r;
reg csrbank0_scratch0_we;
wire [31:0] csrbank0_scratch0_w;
reg csrbank0_bus_errors_re;
wire [31:0] csrbank0_bus_errors_r;
reg csrbank0_bus_errors_we;
wire [31:0] csrbank0_bus_errors_w;
wire csrbank0_sel;
wire [13:0] interface1_bank_bus_adr;
wire interface1_bank_bus_we;
wire [31:0] interface1_bank_bus_dat_w;
reg [31:0] interface1_bank_bus_dat_r;
reg csrbank1_out0_re;
wire csrbank1_out0_r;
reg csrbank1_out0_we;
wire csrbank1_out0_w;
wire csrbank1_sel;
wire [13:0] interface2_bank_bus_adr;
wire interface2_bank_bus_we;
wire [31:0] interface2_bank_bus_dat_w;
reg [31:0] interface2_bank_bus_dat_r;
reg csrbank2_out0_re;
wire csrbank2_out0_r;
reg csrbank2_out0_we;
wire csrbank2_out0_w;
wire csrbank2_sel;
wire [13:0] interface3_bank_bus_adr;
wire interface3_bank_bus_we;
wire [31:0] interface3_bank_bus_dat_w;
reg [31:0] interface3_bank_bus_dat_r;
reg csrbank3_mmap_dummy_bits0_re;
wire [7:0] csrbank3_mmap_dummy_bits0_r;
reg csrbank3_mmap_dummy_bits0_we;
wire [7:0] csrbank3_mmap_dummy_bits0_w;
reg csrbank3_master_cs0_re;
wire csrbank3_master_cs0_r;
reg csrbank3_master_cs0_we;
wire csrbank3_master_cs0_w;
reg csrbank3_master_phyconfig0_re;
wire [23:0] csrbank3_master_phyconfig0_r;
reg csrbank3_master_phyconfig0_we;
wire [23:0] csrbank3_master_phyconfig0_w;
reg csrbank3_master_status_re;
wire [1:0] csrbank3_master_status_r;
reg csrbank3_master_status_we;
wire [1:0] csrbank3_master_status_w;
wire csrbank3_sel;
wire [13:0] interface4_bank_bus_adr;
wire interface4_bank_bus_we;
wire [31:0] interface4_bank_bus_dat_w;
reg [31:0] interface4_bank_bus_dat_r;
reg csrbank4_clk_divisor0_re;
wire [7:0] csrbank4_clk_divisor0_r;
reg csrbank4_clk_divisor0_we;
wire [7:0] csrbank4_clk_divisor0_w;
wire csrbank4_sel;
wire [13:0] interface5_bank_bus_adr;
wire interface5_bank_bus_we;
wire [31:0] interface5_bank_bus_dat_w;
reg [31:0] interface5_bank_bus_dat_r;
reg csrbank5_mode10_re;
wire csrbank5_mode10_r;
reg csrbank5_mode10_we;
wire csrbank5_mode10_w;
reg csrbank5_mode00_re;
wire csrbank5_mode00_r;
reg csrbank5_mode00_we;
wire csrbank5_mode00_w;
reg csrbank5_ien0_re;
wire csrbank5_ien0_r;
reg csrbank5_ien0_we;
wire csrbank5_ien0_w;
reg csrbank5_oe0_re;
wire csrbank5_oe0_r;
reg csrbank5_oe0_we;
wire csrbank5_oe0_w;
reg csrbank5_in_re;
wire csrbank5_in_r;
reg csrbank5_in_we;
wire csrbank5_in_w;
reg csrbank5_out0_re;
wire csrbank5_out0_r;
reg csrbank5_out0_we;
wire csrbank5_out0_w;
wire csrbank5_sel;
wire [13:0] interface6_bank_bus_adr;
wire interface6_bank_bus_we;
wire [31:0] interface6_bank_bus_dat_w;
reg [31:0] interface6_bank_bus_dat_r;
reg csrbank6_ien3_re;
wire [31:0] csrbank6_ien3_r;
reg csrbank6_ien3_we;
wire [31:0] csrbank6_ien3_w;
reg csrbank6_ien2_re;
wire [31:0] csrbank6_ien2_r;
reg csrbank6_ien2_we;
wire [31:0] csrbank6_ien2_w;
reg csrbank6_ien1_re;
wire [31:0] csrbank6_ien1_r;
reg csrbank6_ien1_we;
wire [31:0] csrbank6_ien1_w;
reg csrbank6_ien0_re;
wire [31:0] csrbank6_ien0_r;
reg csrbank6_ien0_we;
wire [31:0] csrbank6_ien0_w;
reg csrbank6_oe3_re;
wire [31:0] csrbank6_oe3_r;
reg csrbank6_oe3_we;
wire [31:0] csrbank6_oe3_w;
reg csrbank6_oe2_re;
wire [31:0] csrbank6_oe2_r;
reg csrbank6_oe2_we;
wire [31:0] csrbank6_oe2_w;
reg csrbank6_oe1_re;
wire [31:0] csrbank6_oe1_r;
reg csrbank6_oe1_we;
wire [31:0] csrbank6_oe1_w;
reg csrbank6_oe0_re;
wire [31:0] csrbank6_oe0_r;
reg csrbank6_oe0_we;
wire [31:0] csrbank6_oe0_w;
reg csrbank6_in3_re;
wire [31:0] csrbank6_in3_r;
reg csrbank6_in3_we;
wire [31:0] csrbank6_in3_w;
reg csrbank6_in2_re;
wire [31:0] csrbank6_in2_r;
reg csrbank6_in2_we;
wire [31:0] csrbank6_in2_w;
reg csrbank6_in1_re;
wire [31:0] csrbank6_in1_r;
reg csrbank6_in1_we;
wire [31:0] csrbank6_in1_w;
reg csrbank6_in0_re;
wire [31:0] csrbank6_in0_r;
reg csrbank6_in0_we;
wire [31:0] csrbank6_in0_w;
reg csrbank6_out3_re;
wire [31:0] csrbank6_out3_r;
reg csrbank6_out3_we;
wire [31:0] csrbank6_out3_w;
reg csrbank6_out2_re;
wire [31:0] csrbank6_out2_r;
reg csrbank6_out2_we;
wire [31:0] csrbank6_out2_w;
reg csrbank6_out1_re;
wire [31:0] csrbank6_out1_r;
reg csrbank6_out1_we;
wire [31:0] csrbank6_out1_w;
reg csrbank6_out0_re;
wire [31:0] csrbank6_out0_r;
reg csrbank6_out0_we;
wire [31:0] csrbank6_out0_w;
wire csrbank6_sel;
wire [13:0] interface7_bank_bus_adr;
wire interface7_bank_bus_we;
wire [31:0] interface7_bank_bus_dat_w;
reg [31:0] interface7_bank_bus_dat_r;
reg csrbank7_out0_re;
wire csrbank7_out0_r;
reg csrbank7_out0_we;
wire csrbank7_out0_w;
wire csrbank7_sel;
wire [13:0] interface8_bank_bus_adr;
wire interface8_bank_bus_we;
wire [31:0] interface8_bank_bus_dat_w;
reg [31:0] interface8_bank_bus_dat_r;
reg csrbank8_out0_re;
wire csrbank8_out0_r;
reg csrbank8_out0_we;
wire csrbank8_out0_w;
wire csrbank8_sel;
wire [13:0] interface9_bank_bus_adr;
wire interface9_bank_bus_we;
wire [31:0] interface9_bank_bus_dat_w;
reg [31:0] interface9_bank_bus_dat_r;
reg csrbank9_control0_re;
wire [15:0] csrbank9_control0_r;
reg csrbank9_control0_we;
wire [15:0] csrbank9_control0_w;
reg csrbank9_status_re;
wire csrbank9_status_r;
reg csrbank9_status_we;
wire csrbank9_status_w;
reg csrbank9_mosi0_re;
wire [7:0] csrbank9_mosi0_r;
reg csrbank9_mosi0_we;
wire [7:0] csrbank9_mosi0_w;
reg csrbank9_miso_re;
wire [7:0] csrbank9_miso_r;
reg csrbank9_miso_we;
wire [7:0] csrbank9_miso_w;
reg csrbank9_cs0_re;
wire [16:0] csrbank9_cs0_r;
reg csrbank9_cs0_we;
wire [16:0] csrbank9_cs0_w;
reg csrbank9_loopback0_re;
wire csrbank9_loopback0_r;
reg csrbank9_loopback0_we;
wire csrbank9_loopback0_w;
reg csrbank9_clk_divider0_re;
wire [15:0] csrbank9_clk_divider0_r;
reg csrbank9_clk_divider0_we;
wire [15:0] csrbank9_clk_divider0_w;
wire csrbank9_sel;
wire [13:0] interface10_bank_bus_adr;
wire interface10_bank_bus_we;
wire [31:0] interface10_bank_bus_dat_w;
reg [31:0] interface10_bank_bus_dat_r;
reg csrbank10_load0_re;
wire [31:0] csrbank10_load0_r;
reg csrbank10_load0_we;
wire [31:0] csrbank10_load0_w;
reg csrbank10_reload0_re;
wire [31:0] csrbank10_reload0_r;
reg csrbank10_reload0_we;
wire [31:0] csrbank10_reload0_w;
reg csrbank10_en0_re;
wire csrbank10_en0_r;
reg csrbank10_en0_we;
wire csrbank10_en0_w;
reg csrbank10_update_value0_re;
wire csrbank10_update_value0_r;
reg csrbank10_update_value0_we;
wire csrbank10_update_value0_w;
reg csrbank10_value_re;
wire [31:0] csrbank10_value_r;
reg csrbank10_value_we;
wire [31:0] csrbank10_value_w;
reg csrbank10_ev_status_re;
wire csrbank10_ev_status_r;
reg csrbank10_ev_status_we;
wire csrbank10_ev_status_w;
reg csrbank10_ev_pending_re;
wire csrbank10_ev_pending_r;
reg csrbank10_ev_pending_we;
wire csrbank10_ev_pending_w;
reg csrbank10_ev_enable0_re;
wire csrbank10_ev_enable0_r;
reg csrbank10_ev_enable0_we;
wire csrbank10_ev_enable0_w;
wire csrbank10_sel;
wire [13:0] interface11_bank_bus_adr;
wire interface11_bank_bus_we;
wire [31:0] interface11_bank_bus_dat_w;
reg [31:0] interface11_bank_bus_dat_r;
reg csrbank11_txfull_re;
wire csrbank11_txfull_r;
reg csrbank11_txfull_we;
wire csrbank11_txfull_w;
reg csrbank11_rxempty_re;
wire csrbank11_rxempty_r;
reg csrbank11_rxempty_we;
wire csrbank11_rxempty_w;
reg csrbank11_ev_status_re;
wire [1:0] csrbank11_ev_status_r;
reg csrbank11_ev_status_we;
wire [1:0] csrbank11_ev_status_w;
reg csrbank11_ev_pending_re;
wire [1:0] csrbank11_ev_pending_r;
reg csrbank11_ev_pending_we;
wire [1:0] csrbank11_ev_pending_w;
reg csrbank11_ev_enable0_re;
wire [1:0] csrbank11_ev_enable0_r;
reg csrbank11_ev_enable0_we;
wire [1:0] csrbank11_ev_enable0_w;
reg csrbank11_txempty_re;
wire csrbank11_txempty_r;
reg csrbank11_txempty_we;
wire csrbank11_txempty_w;
reg csrbank11_rxfull_re;
wire csrbank11_rxfull_r;
reg csrbank11_rxfull_we;
wire csrbank11_rxfull_w;
wire csrbank11_sel;
wire [13:0] interface12_bank_bus_adr;
wire interface12_bank_bus_we;
wire [31:0] interface12_bank_bus_dat_w;
reg [31:0] interface12_bank_bus_dat_r;
reg csrbank12_out0_re;
wire csrbank12_out0_r;
reg csrbank12_out0_we;
wire csrbank12_out0_w;
wire csrbank12_sel;
wire [13:0] interface13_bank_bus_adr;
wire interface13_bank_bus_we;
wire [31:0] interface13_bank_bus_dat_w;
reg [31:0] interface13_bank_bus_dat_r;
reg csrbank13_in_re;
wire csrbank13_in_r;
reg csrbank13_in_we;
wire csrbank13_in_w;
reg csrbank13_mode0_re;
wire csrbank13_mode0_r;
reg csrbank13_mode0_we;
wire csrbank13_mode0_w;
reg csrbank13_edge0_re;
wire csrbank13_edge0_r;
reg csrbank13_edge0_we;
wire csrbank13_edge0_w;
reg csrbank13_ev_status_re;
wire csrbank13_ev_status_r;
reg csrbank13_ev_status_we;
wire csrbank13_ev_status_w;
reg csrbank13_ev_pending_re;
wire csrbank13_ev_pending_r;
reg csrbank13_ev_pending_we;
wire csrbank13_ev_pending_w;
reg csrbank13_ev_enable0_re;
wire csrbank13_ev_enable0_r;
reg csrbank13_ev_enable0_we;
wire csrbank13_ev_enable0_w;
wire csrbank13_sel;
wire [13:0] interface14_bank_bus_adr;
wire interface14_bank_bus_we;
wire [31:0] interface14_bank_bus_dat_w;
reg [31:0] interface14_bank_bus_dat_r;
reg csrbank14_in_re;
wire csrbank14_in_r;
reg csrbank14_in_we;
wire csrbank14_in_w;
reg csrbank14_mode0_re;
wire csrbank14_mode0_r;
reg csrbank14_mode0_we;
wire csrbank14_mode0_w;
reg csrbank14_edge0_re;
wire csrbank14_edge0_r;
reg csrbank14_edge0_we;
wire csrbank14_edge0_w;
reg csrbank14_ev_status_re;
wire csrbank14_ev_status_r;
reg csrbank14_ev_status_we;
wire csrbank14_ev_status_w;
reg csrbank14_ev_pending_re;
wire csrbank14_ev_pending_r;
reg csrbank14_ev_pending_we;
wire csrbank14_ev_pending_w;
reg csrbank14_ev_enable0_re;
wire csrbank14_ev_enable0_r;
reg csrbank14_ev_enable0_we;
wire csrbank14_ev_enable0_w;
wire csrbank14_sel;
wire [13:0] interface15_bank_bus_adr;
wire interface15_bank_bus_we;
wire [31:0] interface15_bank_bus_dat_w;
reg [31:0] interface15_bank_bus_dat_r;
reg csrbank15_in_re;
wire csrbank15_in_r;
reg csrbank15_in_we;
wire csrbank15_in_w;
reg csrbank15_mode0_re;
wire csrbank15_mode0_r;
reg csrbank15_mode0_we;
wire csrbank15_mode0_w;
reg csrbank15_edge0_re;
wire csrbank15_edge0_r;
reg csrbank15_edge0_we;
wire csrbank15_edge0_w;
reg csrbank15_ev_status_re;
wire csrbank15_ev_status_r;
reg csrbank15_ev_status_we;
wire csrbank15_ev_status_w;
reg csrbank15_ev_pending_re;
wire csrbank15_ev_pending_r;
reg csrbank15_ev_pending_we;
wire csrbank15_ev_pending_w;
reg csrbank15_ev_enable0_re;
wire csrbank15_ev_enable0_r;
reg csrbank15_ev_enable0_we;
wire csrbank15_ev_enable0_w;
wire csrbank15_sel;
wire [13:0] interface16_bank_bus_adr;
wire interface16_bank_bus_we;
wire [31:0] interface16_bank_bus_dat_w;
reg [31:0] interface16_bank_bus_dat_r;
reg csrbank16_in_re;
wire csrbank16_in_r;
reg csrbank16_in_we;
wire csrbank16_in_w;
reg csrbank16_mode0_re;
wire csrbank16_mode0_r;
reg csrbank16_mode0_we;
wire csrbank16_mode0_w;
reg csrbank16_edge0_re;
wire csrbank16_edge0_r;
reg csrbank16_edge0_we;
wire csrbank16_edge0_w;
reg csrbank16_ev_status_re;
wire csrbank16_ev_status_r;
reg csrbank16_ev_status_we;
wire csrbank16_ev_status_w;
reg csrbank16_ev_pending_re;
wire csrbank16_ev_pending_r;
reg csrbank16_ev_pending_we;
wire csrbank16_ev_pending_w;
reg csrbank16_ev_enable0_re;
wire csrbank16_ev_enable0_r;
reg csrbank16_ev_enable0_we;
wire csrbank16_ev_enable0_w;
wire csrbank16_sel;
wire [13:0] interface17_bank_bus_adr;
wire interface17_bank_bus_we;
wire [31:0] interface17_bank_bus_dat_w;
reg [31:0] interface17_bank_bus_dat_r;
reg csrbank17_in_re;
wire csrbank17_in_r;
reg csrbank17_in_we;
wire csrbank17_in_w;
reg csrbank17_mode0_re;
wire csrbank17_mode0_r;
reg csrbank17_mode0_we;
wire csrbank17_mode0_w;
reg csrbank17_edge0_re;
wire csrbank17_edge0_r;
reg csrbank17_edge0_we;
wire csrbank17_edge0_w;
reg csrbank17_ev_status_re;
wire csrbank17_ev_status_r;
reg csrbank17_ev_status_we;
wire csrbank17_ev_status_w;
reg csrbank17_ev_pending_re;
wire csrbank17_ev_pending_r;
reg csrbank17_ev_pending_we;
wire csrbank17_ev_pending_w;
reg csrbank17_ev_enable0_re;
wire csrbank17_ev_enable0_r;
reg csrbank17_ev_enable0_we;
wire csrbank17_ev_enable0_w;
wire csrbank17_sel;
wire [13:0] interface18_bank_bus_adr;
wire interface18_bank_bus_we;
wire [31:0] interface18_bank_bus_dat_w;
reg [31:0] interface18_bank_bus_dat_r;
reg csrbank18_in_re;
wire csrbank18_in_r;
reg csrbank18_in_we;
wire csrbank18_in_w;
reg csrbank18_mode0_re;
wire csrbank18_mode0_r;
reg csrbank18_mode0_we;
wire csrbank18_mode0_w;
reg csrbank18_edge0_re;
wire csrbank18_edge0_r;
reg csrbank18_edge0_we;
wire csrbank18_edge0_w;
reg csrbank18_ev_status_re;
wire csrbank18_ev_status_r;
reg csrbank18_ev_status_we;
wire csrbank18_ev_status_w;
reg csrbank18_ev_pending_re;
wire csrbank18_ev_pending_r;
reg csrbank18_ev_pending_we;
wire csrbank18_ev_pending_w;
reg csrbank18_ev_enable0_re;
wire csrbank18_ev_enable0_r;
reg csrbank18_ev_enable0_we;
wire csrbank18_ev_enable0_w;
wire csrbank18_sel;
wire [13:0] interface19_bank_bus_adr;
wire interface19_bank_bus_we;
wire [31:0] interface19_bank_bus_dat_w;
reg [31:0] interface19_bank_bus_dat_r;
reg csrbank19_out0_re;
wire [2:0] csrbank19_out0_r;
reg csrbank19_out0_we;
wire [2:0] csrbank19_out0_w;
wire csrbank19_sel;
wire [13:0] csr_interconnect_adr;
wire csr_interconnect_we;
wire [31:0] csr_interconnect_dat_w;
wire [31:0] csr_interconnect_dat_r;
reg state;
reg next_state;
reg [29:0] comb_array_muxed0;
reg [31:0] comb_array_muxed1;
reg [3:0] comb_array_muxed2;
reg comb_array_muxed3;
reg comb_array_muxed4;
reg comb_array_muxed5;
reg [2:0] comb_array_muxed6;
reg [1:0] comb_array_muxed7;
reg sync_array_muxed;
wire sdrio_clk;
wire sdrio_clk_1;
wire sdrio_clk_2;
wire sdrio_clk_3;
reg multiregimpl0_regs0;
reg multiregimpl0_regs1;
reg multiregimpl1_regs0;
reg multiregimpl1_regs1;
reg multiregimpl2_regs0;
reg multiregimpl2_regs1;
reg multiregimpl3_regs0;
reg multiregimpl3_regs1;
reg multiregimpl4_regs0;
reg multiregimpl4_regs1;
reg multiregimpl5_regs0;
reg multiregimpl5_regs1;
reg multiregimpl6_regs0;
reg multiregimpl6_regs1;
reg multiregimpl7_regs0;
reg multiregimpl7_regs1;
reg multiregimpl8_regs0;
reg multiregimpl8_regs1;
reg multiregimpl9_regs0;
reg multiregimpl9_regs1;
reg multiregimpl10_regs0;
reg multiregimpl10_regs1;
reg multiregimpl11_regs0;
reg multiregimpl11_regs1;
reg multiregimpl12_regs0;
reg multiregimpl12_regs1;
reg multiregimpl13_regs0;
reg multiregimpl13_regs1;
reg multiregimpl14_regs0;
reg multiregimpl14_regs1;
reg multiregimpl15_regs0;
reg multiregimpl15_regs1;
reg multiregimpl16_regs0;
reg multiregimpl16_regs1;
reg multiregimpl17_regs0;
reg multiregimpl17_regs1;
reg multiregimpl18_regs0;
reg multiregimpl18_regs1;
reg multiregimpl19_regs0;
reg multiregimpl19_regs1;
reg multiregimpl20_regs0;
reg multiregimpl20_regs1;
reg multiregimpl21_regs0;
reg multiregimpl21_regs1;
reg multiregimpl22_regs0;
reg multiregimpl22_regs1;
reg multiregimpl23_regs0;
reg multiregimpl23_regs1;
reg multiregimpl24_regs0;
reg multiregimpl24_regs1;
reg multiregimpl25_regs0;
reg multiregimpl25_regs1;
reg multiregimpl26_regs0;
reg multiregimpl26_regs1;
reg multiregimpl27_regs0;
reg multiregimpl27_regs1;
reg multiregimpl28_regs0;
reg multiregimpl28_regs1;
reg multiregimpl29_regs0;
reg multiregimpl29_regs1;
reg multiregimpl30_regs0;
reg multiregimpl30_regs1;
reg multiregimpl31_regs0;
reg multiregimpl31_regs1;
reg multiregimpl32_regs0;
reg multiregimpl32_regs1;
reg multiregimpl33_regs0;
reg multiregimpl33_regs1;
reg multiregimpl34_regs0;
reg multiregimpl34_regs1;
reg multiregimpl35_regs0;
reg multiregimpl35_regs1;
reg multiregimpl36_regs0;
reg multiregimpl36_regs1;
reg multiregimpl37_regs0;
reg multiregimpl37_regs1;
reg multiregimpl38_regs0;
reg multiregimpl38_regs1;
reg multiregimpl39_regs0;
reg multiregimpl39_regs1;
reg multiregimpl40_regs0;
reg multiregimpl40_regs1;
reg multiregimpl41_regs0;
reg multiregimpl41_regs1;
reg multiregimpl42_regs0;
reg multiregimpl42_regs1;
reg multiregimpl43_regs0;
reg multiregimpl43_regs1;
reg multiregimpl44_regs0;
reg multiregimpl44_regs1;
reg multiregimpl45_regs0;
reg multiregimpl45_regs1;
reg multiregimpl46_regs0;
reg multiregimpl46_regs1;
reg multiregimpl47_regs0;
reg multiregimpl47_regs1;
reg multiregimpl48_regs0;
reg multiregimpl48_regs1;
reg multiregimpl49_regs0;
reg multiregimpl49_regs1;
reg multiregimpl50_regs0;
reg multiregimpl50_regs1;
reg multiregimpl51_regs0;
reg multiregimpl51_regs1;
reg multiregimpl52_regs0;
reg multiregimpl52_regs1;
reg multiregimpl53_regs0;
reg multiregimpl53_regs1;
reg multiregimpl54_regs0;
reg multiregimpl54_regs1;
reg multiregimpl55_regs0;
reg multiregimpl55_regs1;
reg multiregimpl56_regs0;
reg multiregimpl56_regs1;
reg multiregimpl57_regs0;
reg multiregimpl57_regs1;
reg multiregimpl58_regs0;
reg multiregimpl58_regs1;
reg multiregimpl59_regs0;
reg multiregimpl59_regs1;
reg multiregimpl60_regs0;
reg multiregimpl60_regs1;
reg multiregimpl61_regs0;
reg multiregimpl61_regs1;
reg multiregimpl62_regs0;
reg multiregimpl62_regs1;
reg multiregimpl63_regs0;
reg multiregimpl63_regs1;
reg multiregimpl64_regs0;
reg multiregimpl64_regs1;
reg multiregimpl65_regs0;
reg multiregimpl65_regs1;
reg multiregimpl66_regs0;
reg multiregimpl66_regs1;
reg multiregimpl67_regs0;
reg multiregimpl67_regs1;
reg multiregimpl68_regs0;
reg multiregimpl68_regs1;
reg multiregimpl69_regs0;
reg multiregimpl69_regs1;
reg multiregimpl70_regs0;
reg multiregimpl70_regs1;
reg multiregimpl71_regs0;
reg multiregimpl71_regs1;
reg multiregimpl72_regs0;
reg multiregimpl72_regs1;
reg multiregimpl73_regs0;
reg multiregimpl73_regs1;
reg multiregimpl74_regs0;
reg multiregimpl74_regs1;
reg multiregimpl75_regs0;
reg multiregimpl75_regs1;
reg multiregimpl76_regs0;
reg multiregimpl76_regs1;
reg multiregimpl77_regs0;
reg multiregimpl77_regs1;
reg multiregimpl78_regs0;
reg multiregimpl78_regs1;
reg multiregimpl79_regs0;
reg multiregimpl79_regs1;
reg multiregimpl80_regs0;
reg multiregimpl80_regs1;
reg multiregimpl81_regs0;
reg multiregimpl81_regs1;
reg multiregimpl82_regs0;
reg multiregimpl82_regs1;
reg multiregimpl83_regs0;
reg multiregimpl83_regs1;
reg multiregimpl84_regs0;
reg multiregimpl84_regs1;
reg multiregimpl85_regs0;
reg multiregimpl85_regs1;
reg multiregimpl86_regs0;
reg multiregimpl86_regs1;
reg multiregimpl87_regs0;
reg multiregimpl87_regs1;
reg multiregimpl88_regs0;
reg multiregimpl88_regs1;
reg multiregimpl89_regs0;
reg multiregimpl89_regs1;
reg multiregimpl90_regs0;
reg multiregimpl90_regs1;
reg multiregimpl91_regs0;
reg multiregimpl91_regs1;
reg multiregimpl92_regs0;
reg multiregimpl92_regs1;
reg multiregimpl93_regs0;
reg multiregimpl93_regs1;
reg multiregimpl94_regs0;
reg multiregimpl94_regs1;
reg multiregimpl95_regs0;
reg multiregimpl95_regs1;
reg multiregimpl96_regs0;
reg multiregimpl96_regs1;
reg multiregimpl97_regs0;
reg multiregimpl97_regs1;
reg multiregimpl98_regs0;
reg multiregimpl98_regs1;
reg multiregimpl99_regs0;
reg multiregimpl99_regs1;
reg multiregimpl100_regs0;
reg multiregimpl100_regs1;
reg multiregimpl101_regs0;
reg multiregimpl101_regs1;
reg multiregimpl102_regs0;
reg multiregimpl102_regs1;
reg multiregimpl103_regs0;
reg multiregimpl103_regs1;
reg multiregimpl104_regs0;
reg multiregimpl104_regs1;
reg multiregimpl105_regs0;
reg multiregimpl105_regs1;
reg multiregimpl106_regs0;
reg multiregimpl106_regs1;
reg multiregimpl107_regs0;
reg multiregimpl107_regs1;
reg multiregimpl108_regs0;
reg multiregimpl108_regs1;
reg multiregimpl109_regs0;
reg multiregimpl109_regs1;
reg multiregimpl110_regs0;
reg multiregimpl110_regs1;
reg multiregimpl111_regs0;
reg multiregimpl111_regs1;
reg multiregimpl112_regs0;
reg multiregimpl112_regs1;
reg multiregimpl113_regs0;
reg multiregimpl113_regs1;
reg multiregimpl114_regs0;
reg multiregimpl114_regs1;
reg multiregimpl115_regs0;
reg multiregimpl115_regs1;
reg multiregimpl116_regs0;
reg multiregimpl116_regs1;
reg multiregimpl117_regs0;
reg multiregimpl117_regs1;
reg multiregimpl118_regs0;
reg multiregimpl118_regs1;
reg multiregimpl119_regs0;
reg multiregimpl119_regs1;
reg multiregimpl120_regs0;
reg multiregimpl120_regs1;
reg multiregimpl121_regs0;
reg multiregimpl121_regs1;
reg multiregimpl122_regs0;
reg multiregimpl122_regs1;
reg multiregimpl123_regs0;
reg multiregimpl123_regs1;
reg multiregimpl124_regs0;
reg multiregimpl124_regs1;
reg multiregimpl125_regs0;
reg multiregimpl125_regs1;
reg multiregimpl126_regs0;
reg multiregimpl126_regs1;
reg multiregimpl127_regs0;
reg multiregimpl127_regs1;
reg multiregimpl128_regs0;
reg multiregimpl128_regs1;
reg multiregimpl129_regs0;
reg multiregimpl129_regs1;
reg multiregimpl130_regs0;
reg multiregimpl130_regs1;
reg multiregimpl131_regs0;
reg multiregimpl131_regs1;
reg multiregimpl132_regs0;
reg multiregimpl132_regs1;
reg multiregimpl133_regs0;
reg multiregimpl133_regs1;
reg multiregimpl134_regs0;
reg multiregimpl134_regs1;
reg multiregimpl135_regs0;
reg multiregimpl135_regs1;
reg multiregimpl136_regs0;
reg multiregimpl136_regs1;

assign core_rst = (~core_rstn);
assign mgmtsoc_reset = (mgmtsoc_soc_rst | mgmtsoc_cpu_rst);
assign spi_sdoenb = (~spi_cs_n);
assign mprj_cyc_o = mprj_cyc;
assign mprj_stb_o = mprj_stb;
assign mprj_we_o = mprj_we;
assign mprj_sel_o = mprj_sel;
always @(*) begin
	mprj_adr_o = 32'd0;
	mprj_adr_o[31:2] = mprj_adr;
	mprj_adr_o[1:0] = 1'd0;
end
assign mprj_dat_r = mprj_dat_i;
assign mprj_dat_o = mprj_dat_w;
assign mprj_ack = mprj_ack_i;
assign hk_stb_o = hk_stb;
assign hk_cyc_o = hk_cyc;
assign hk_dat_r = hk_dat_i;
assign hk_ack = hk_ack_i;
assign debug_out = 1'd0;
always @(*) begin
	sys_uart_rx = 1'd0;
	if ((debug_in == 1'd1)) begin
	end else begin
		sys_uart_rx = serial_rx;
	end
end
always @(*) begin
	dbg_uart_dbg_uart_rx = 1'd0;
	if ((debug_in == 1'd1)) begin
		dbg_uart_dbg_uart_rx = serial_rx;
	end else begin
	end
end
always @(*) begin
	serial_tx = 1'd0;
	if ((debug_in == 1'd1)) begin
		serial_tx = dbg_uart_dbg_uart_tx;
	end else begin
		serial_tx = sys_uart_tx;
	end
end
assign uart_enabled = (uart_enabled_o | debug_in);
assign qspi_enabled = 1'd0;
assign trap = 1'd0;

assign clk_out = clk_in;
assign resetn_out = resetn_in;
assign serial_load_out = serial_load_in;
assign serial_data_2_out = serial_data_2_in;
assign serial_resetn_out = serial_resetn_in;
assign serial_clock_out = serial_clock_in;
assign rstb_l_out = rstb_l_in;

// [Vic]: POR is useless here
//assign por_l_out = por_l_in;
//assign porb_h_out = porb_h_in;

assign mgmtsoc_bus_error = error;
always @(*) begin
	mgmtsoc_interrupt = 32'd0;
	mgmtsoc_interrupt[0] = mgmtsoc_irq;
	mgmtsoc_interrupt[1] = uart_irq;
	mgmtsoc_interrupt[2] = gpioin0_gpioin0_irq;
	mgmtsoc_interrupt[3] = gpioin1_gpioin1_irq;
	mgmtsoc_interrupt[4] = gpioin2_gpioin2_irq;
	mgmtsoc_interrupt[5] = gpioin3_gpioin3_irq;
	mgmtsoc_interrupt[6] = gpioin4_gpioin4_irq;
	mgmtsoc_interrupt[7] = gpioin5_gpioin5_irq;
end
assign sys_clk = core_clk;
assign por_clk = core_clk;
assign sys_rst = int_rst;
assign mgmtsoc_bus_errors_status = mgmtsoc_bus_errors;
assign mgmtsoc_zero_trigger = (mgmtsoc_value == 1'd0);
assign mgmtsoc_zero0 = mgmtsoc_zero_status;
assign mgmtsoc_zero1 = mgmtsoc_zero_pending;
always @(*) begin
	mgmtsoc_zero_clear = 1'd0;
	if ((mgmtsoc_pending_re & mgmtsoc_pending_r)) begin
		mgmtsoc_zero_clear = 1'd1;
	end
end
assign mgmtsoc_irq = (mgmtsoc_pending_status & mgmtsoc_enable_storage);
assign mgmtsoc_zero_status = mgmtsoc_zero_trigger;
assign dff_di = dff_bus_dat_w[31:0];
always @(*) begin
	dff_we = 4'd0;
	dff_we[0] = (((dff_bus_sel[0] & dff_bus_we) & dff_bus_stb) & dff_bus_cyc);
	dff_we[1] = (((dff_bus_sel[1] & dff_bus_we) & dff_bus_stb) & dff_bus_cyc);
	dff_we[2] = (((dff_bus_sel[2] & dff_bus_we) & dff_bus_stb) & dff_bus_cyc);
	dff_we[3] = (((dff_bus_sel[3] & dff_bus_we) & dff_bus_stb) & dff_bus_cyc);
end
assign dff_bus_dat_r[31:0] = dff_do;
assign dff_en = (dff_bus_stb & dff_bus_cyc);
assign dff2_di = dff2_bus_dat_w[31:0];
always @(*) begin
	dff2_we = 4'd0;
	dff2_we[0] = (((dff2_bus_sel[0] & dff2_bus_we) & dff2_bus_stb) & dff2_bus_cyc);
	dff2_we[1] = (((dff2_bus_sel[1] & dff2_bus_we) & dff2_bus_stb) & dff2_bus_cyc);
	dff2_we[2] = (((dff2_bus_sel[2] & dff2_bus_we) & dff2_bus_stb) & dff2_bus_cyc);
	dff2_we[3] = (((dff2_bus_sel[3] & dff2_bus_we) & dff2_bus_stb) & dff2_bus_cyc);
end
assign dff2_bus_dat_r[31:0] = dff2_do;
assign dff2_en = (dff2_bus_stb & dff2_bus_cyc);
assign mgmtsoc_litespisdrphycore_div = mgmtsoc_litespisdrphycore_spi_clk_divisor;
assign mgmtsoc_litespisdrphycore_sample_cnt = 1'd1;
assign mgmtsoc_litespisdrphycore_update_cnt = 1'd1;
assign mgmtsoc_litespisdrphycore_wait = mgmtsoc_litespisdrphycore_cs;
assign mgmtsoc_litespisdrphycore_cs_enable = mgmtsoc_litespisdrphycore_done;
assign flash_cs_n = (~mgmtsoc_litespisdrphycore_cs_enable);
assign flash_io1_oeb = 1'd1;
assign flash_io1_do = 1'd0;
assign flash_io2_do = 1'd0;
assign flash_io3_do = 1'd0;
assign flash_io2_oeb = 1'd1;
assign flash_io3_oeb = 1'd1;
assign mgmtsoc_litespisdrphycore_dq_oe = mgmtsoc_litespisdrphycore_sink_payload_mask;
always @(*) begin
	mgmtsoc_litespisdrphycore_dq_o = 1'd0;
	case (mgmtsoc_litespisdrphycore_sink_payload_width)
		1'd1: begin
			mgmtsoc_litespisdrphycore_dq_o = mgmtsoc_litespisdrphycore_sr_out[31];
		end
		2'd2: begin
			mgmtsoc_litespisdrphycore_dq_o = mgmtsoc_litespisdrphycore_sr_out[31:30];
		end
		3'd4: begin
			mgmtsoc_litespisdrphycore_dq_o = mgmtsoc_litespisdrphycore_sr_out[31:28];
		end
		4'd8: begin
			mgmtsoc_litespisdrphycore_dq_o = mgmtsoc_litespisdrphycore_sr_out[31:24];
		end
	endcase
end
assign mgmtsoc_litespisdrphycore_source_payload_data = mgmtsoc_litespisdrphycore_sr_in;
assign mgmtsoc_litespisdrphycore_spi_clk_divisor = mgmtsoc_litespisdrphycore_storage;
assign mgmtsoc_litespisdrphycore_posedge = ((mgmtsoc_litespisdrphycore_en & (~mgmtsoc_litespisdrphycore_clk)) & (mgmtsoc_litespisdrphycore_cnt == mgmtsoc_litespisdrphycore_div));
assign mgmtsoc_litespisdrphycore_negedge = ((mgmtsoc_litespisdrphycore_en & mgmtsoc_litespisdrphycore_clk) & (mgmtsoc_litespisdrphycore_cnt == mgmtsoc_litespisdrphycore_div));
assign mgmtsoc_litespisdrphycore_sample = (mgmtsoc_litespisdrphycore_cnt == mgmtsoc_litespisdrphycore_sample_cnt);
assign mgmtsoc_litespisdrphycore_update = (mgmtsoc_litespisdrphycore_cnt == mgmtsoc_litespisdrphycore_update_cnt);
assign mgmtsoc_litespisdrphycore_done = (mgmtsoc_litespisdrphycore_count == 1'd0);
always @(*) begin
	litespiphy_next_state = 2'd0;
	litespiphy_next_state = litespiphy_state;
	case (litespiphy_state)
		1'd1: begin
			if (mgmtsoc_litespisdrphycore_negedge) begin
				if ((mgmtsoc_litespisdrphycore_sr_cnt == 1'd0)) begin
					litespiphy_next_state = 2'd2;
				end
			end
		end
		2'd2: begin
			if (((mgmtsoc_litespisdrphycore_spi_clk_divisor > 1'd0) | mgmtsoc_litespisdrphycore_posedge_reg2)) begin
				litespiphy_next_state = 2'd3;
			end
		end
		2'd3: begin
			if (mgmtsoc_litespisdrphycore_source_ready) begin
				litespiphy_next_state = 1'd0;
			end
		end
		default: begin
			if ((mgmtsoc_litespisdrphycore_cs_enable & mgmtsoc_litespisdrphycore_sink_valid)) begin
				litespiphy_next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_sink_ready = 1'd0;
	case (litespiphy_state)
		1'd1: begin
		end
		2'd2: begin
			if (((mgmtsoc_litespisdrphycore_spi_clk_divisor > 1'd0) | mgmtsoc_litespisdrphycore_posedge_reg2)) begin
				mgmtsoc_litespisdrphycore_sink_ready = 1'd1;
			end
		end
		2'd3: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_en = 1'd0;
	case (litespiphy_state)
		1'd1: begin
			mgmtsoc_litespisdrphycore_en = 1'd1;
		end
		2'd2: begin
		end
		2'd3: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value = 8'd0;
	case (litespiphy_state)
		1'd1: begin
			if (mgmtsoc_litespisdrphycore_negedge) begin
				mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value = (mgmtsoc_litespisdrphycore_sr_cnt - mgmtsoc_litespisdrphycore_sink_payload_width);
			end
		end
		2'd2: begin
		end
		2'd3: begin
		end
		default: begin
			if ((mgmtsoc_litespisdrphycore_cs_enable & mgmtsoc_litespisdrphycore_sink_valid)) begin
				mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value = (mgmtsoc_litespisdrphycore_sink_payload_len - mgmtsoc_litespisdrphycore_sink_payload_width);
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_sr_out_load = 1'd0;
	case (litespiphy_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		default: begin
			if ((mgmtsoc_litespisdrphycore_cs_enable & mgmtsoc_litespisdrphycore_sink_valid)) begin
				mgmtsoc_litespisdrphycore_sr_out_load = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value_ce = 1'd0;
	case (litespiphy_state)
		1'd1: begin
			if (mgmtsoc_litespisdrphycore_negedge) begin
				mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value_ce = 1'd1;
			end
		end
		2'd2: begin
		end
		2'd3: begin
		end
		default: begin
			if ((mgmtsoc_litespisdrphycore_cs_enable & mgmtsoc_litespisdrphycore_sink_valid)) begin
				mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value_ce = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_sr_out_shift = 1'd0;
	case (litespiphy_state)
		1'd1: begin
			if (mgmtsoc_litespisdrphycore_negedge) begin
				mgmtsoc_litespisdrphycore_sr_out_shift = 1'd1;
			end
		end
		2'd2: begin
		end
		2'd3: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_sr_in_shift = 1'd0;
	case (litespiphy_state)
		1'd1: begin
			if (mgmtsoc_litespisdrphycore_posedge_reg2) begin
				mgmtsoc_litespisdrphycore_sr_in_shift = 1'd1;
			end
		end
		2'd2: begin
			if (((mgmtsoc_litespisdrphycore_spi_clk_divisor > 1'd0) | mgmtsoc_litespisdrphycore_posedge_reg2)) begin
				mgmtsoc_litespisdrphycore_sr_in_shift = (mgmtsoc_litespisdrphycore_spi_clk_divisor == 1'd0);
			end
		end
		2'd3: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_source_valid = 1'd0;
	case (litespiphy_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespisdrphycore_source_valid = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_source_last = 1'd0;
	case (litespiphy_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespisdrphycore_source_last = 1'd1;
		end
		default: begin
		end
	endcase
end
assign mgmtsoc_litespisdrphycore_cs = mgmtsoc_crossbar_cs;
assign mgmtsoc_litespimmap_sink_valid = mgmtsoc_port_mmap_user_port_source_valid;
assign mgmtsoc_port_mmap_user_port_source_ready = mgmtsoc_litespimmap_sink_ready;
assign mgmtsoc_litespimmap_sink_first = mgmtsoc_port_mmap_user_port_source_first;
assign mgmtsoc_litespimmap_sink_last = mgmtsoc_port_mmap_user_port_source_last;
assign mgmtsoc_litespimmap_sink_payload_data = mgmtsoc_port_mmap_user_port_source_payload_data;
assign mgmtsoc_port_mmap_user_port_sink_valid = mgmtsoc_litespimmap_source_valid;
assign mgmtsoc_litespimmap_source_ready = mgmtsoc_port_mmap_user_port_sink_ready;
assign mgmtsoc_port_mmap_user_port_sink_first = mgmtsoc_litespimmap_source_first;
assign mgmtsoc_port_mmap_user_port_sink_last = mgmtsoc_litespimmap_source_last;
assign mgmtsoc_port_mmap_user_port_sink_payload_data = mgmtsoc_litespimmap_source_payload_data;
assign mgmtsoc_port_mmap_user_port_sink_payload_len = mgmtsoc_litespimmap_source_payload_len;
assign mgmtsoc_port_mmap_user_port_sink_payload_width = mgmtsoc_litespimmap_source_payload_width;
assign mgmtsoc_port_mmap_user_port_sink_payload_mask = mgmtsoc_litespimmap_source_payload_mask;
assign mgmtsoc_master_sink_sink_valid = mgmtsoc_port_master_user_port_source_valid;
assign mgmtsoc_port_master_user_port_source_ready = mgmtsoc_master_sink_sink_ready;
assign mgmtsoc_master_sink_sink_first = mgmtsoc_port_master_user_port_source_first;
assign mgmtsoc_master_sink_sink_last = mgmtsoc_port_master_user_port_source_last;
assign mgmtsoc_master_sink_sink_payload_data = mgmtsoc_port_master_user_port_source_payload_data;
assign mgmtsoc_port_master_user_port_sink_valid = mgmtsoc_master_source_source_valid;
assign mgmtsoc_master_source_source_ready = mgmtsoc_port_master_user_port_sink_ready;
assign mgmtsoc_port_master_user_port_sink_first = mgmtsoc_master_source_source_first;
assign mgmtsoc_port_master_user_port_sink_last = mgmtsoc_master_source_source_last;
assign mgmtsoc_port_master_user_port_sink_payload_data = mgmtsoc_master_source_source_payload_data;
assign mgmtsoc_port_master_user_port_sink_payload_len = mgmtsoc_master_source_source_payload_len;
assign mgmtsoc_port_master_user_port_sink_payload_width = mgmtsoc_master_source_source_payload_width;
assign mgmtsoc_port_master_user_port_sink_payload_mask = mgmtsoc_master_source_source_payload_mask;
assign mgmtsoc_litespisdrphycore_sink_valid = mgmtsoc_crossbar_source_valid;
assign mgmtsoc_crossbar_source_ready = mgmtsoc_litespisdrphycore_sink_ready;
assign mgmtsoc_litespisdrphycore_sink_first = mgmtsoc_crossbar_source_first;
assign mgmtsoc_litespisdrphycore_sink_last = mgmtsoc_crossbar_source_last;
assign mgmtsoc_litespisdrphycore_sink_payload_data = mgmtsoc_crossbar_source_payload_data;
assign mgmtsoc_litespisdrphycore_sink_payload_len = mgmtsoc_crossbar_source_payload_len;
assign mgmtsoc_litespisdrphycore_sink_payload_width = mgmtsoc_crossbar_source_payload_width;
assign mgmtsoc_litespisdrphycore_sink_payload_mask = mgmtsoc_crossbar_source_payload_mask;
assign mgmtsoc_crossbar_sink_valid = mgmtsoc_litespisdrphycore_source_valid;
assign mgmtsoc_litespisdrphycore_source_ready = mgmtsoc_crossbar_sink_ready;
assign mgmtsoc_crossbar_sink_first = mgmtsoc_litespisdrphycore_source_first;
assign mgmtsoc_crossbar_sink_last = mgmtsoc_litespisdrphycore_source_last;
assign mgmtsoc_crossbar_sink_payload_data = mgmtsoc_litespisdrphycore_source_payload_data;
assign mgmtsoc_port_mmap_internal_port_sink_valid = mgmtsoc_port_mmap_user_port_sink_valid;
assign mgmtsoc_port_mmap_user_port_sink_ready = mgmtsoc_port_mmap_internal_port_sink_ready;
assign mgmtsoc_port_mmap_internal_port_sink_first = mgmtsoc_port_mmap_user_port_sink_first;
assign mgmtsoc_port_mmap_internal_port_sink_last = mgmtsoc_port_mmap_user_port_sink_last;
assign mgmtsoc_port_mmap_internal_port_sink_payload_data = mgmtsoc_port_mmap_user_port_sink_payload_data;
assign mgmtsoc_port_mmap_internal_port_sink_payload_len = mgmtsoc_port_mmap_user_port_sink_payload_len;
assign mgmtsoc_port_mmap_internal_port_sink_payload_width = mgmtsoc_port_mmap_user_port_sink_payload_width;
assign mgmtsoc_port_mmap_internal_port_sink_payload_mask = mgmtsoc_port_mmap_user_port_sink_payload_mask;
assign mgmtsoc_port_mmap_user_port_source_valid = mgmtsoc_port_mmap_internal_port_source_valid;
assign mgmtsoc_port_mmap_internal_port_source_ready = mgmtsoc_port_mmap_user_port_source_ready;
assign mgmtsoc_port_mmap_user_port_source_first = mgmtsoc_port_mmap_internal_port_source_first;
assign mgmtsoc_port_mmap_user_port_source_last = mgmtsoc_port_mmap_internal_port_source_last;
assign mgmtsoc_port_mmap_user_port_source_payload_data = mgmtsoc_port_mmap_internal_port_source_payload_data;
assign mgmtsoc_port_mmap_request = mgmtsoc_litespimmap_cs;
assign mgmtsoc_port_master_internal_port_sink_valid = mgmtsoc_port_master_user_port_sink_valid;
assign mgmtsoc_port_master_user_port_sink_ready = mgmtsoc_port_master_internal_port_sink_ready;
assign mgmtsoc_port_master_internal_port_sink_first = mgmtsoc_port_master_user_port_sink_first;
assign mgmtsoc_port_master_internal_port_sink_last = mgmtsoc_port_master_user_port_sink_last;
assign mgmtsoc_port_master_internal_port_sink_payload_data = mgmtsoc_port_master_user_port_sink_payload_data;
assign mgmtsoc_port_master_internal_port_sink_payload_len = mgmtsoc_port_master_user_port_sink_payload_len;
assign mgmtsoc_port_master_internal_port_sink_payload_width = mgmtsoc_port_master_user_port_sink_payload_width;
assign mgmtsoc_port_master_internal_port_sink_payload_mask = mgmtsoc_port_master_user_port_sink_payload_mask;
assign mgmtsoc_port_master_user_port_source_valid = mgmtsoc_port_master_internal_port_source_valid;
assign mgmtsoc_port_master_internal_port_source_ready = mgmtsoc_port_master_user_port_source_ready;
assign mgmtsoc_port_master_user_port_source_first = mgmtsoc_port_master_internal_port_source_first;
assign mgmtsoc_port_master_user_port_source_last = mgmtsoc_port_master_internal_port_source_last;
assign mgmtsoc_port_master_user_port_source_payload_data = mgmtsoc_port_master_internal_port_source_payload_data;
assign mgmtsoc_port_master_request = mgmtsoc_master_cs;
assign litespi_tx_mux_endpoint0_sink_valid = mgmtsoc_port_mmap_internal_port_sink_valid;
assign mgmtsoc_port_mmap_internal_port_sink_ready = litespi_tx_mux_endpoint0_sink_ready;
assign litespi_tx_mux_endpoint0_sink_first = mgmtsoc_port_mmap_internal_port_sink_first;
assign litespi_tx_mux_endpoint0_sink_last = mgmtsoc_port_mmap_internal_port_sink_last;
assign litespi_tx_mux_endpoint0_sink_payload_data = mgmtsoc_port_mmap_internal_port_sink_payload_data;
assign litespi_tx_mux_endpoint0_sink_payload_len = mgmtsoc_port_mmap_internal_port_sink_payload_len;
assign litespi_tx_mux_endpoint0_sink_payload_width = mgmtsoc_port_mmap_internal_port_sink_payload_width;
assign litespi_tx_mux_endpoint0_sink_payload_mask = mgmtsoc_port_mmap_internal_port_sink_payload_mask;
assign mgmtsoc_port_mmap_internal_port_source_valid = litespi_rx_demux_endpoint0_source_valid;
assign litespi_rx_demux_endpoint0_source_ready = mgmtsoc_port_mmap_internal_port_source_ready;
assign mgmtsoc_port_mmap_internal_port_source_first = litespi_rx_demux_endpoint0_source_first;
assign mgmtsoc_port_mmap_internal_port_source_last = litespi_rx_demux_endpoint0_source_last;
assign mgmtsoc_port_mmap_internal_port_source_payload_data = litespi_rx_demux_endpoint0_source_payload_data;
assign litespi_tx_mux_endpoint1_sink_valid = mgmtsoc_port_master_internal_port_sink_valid;
assign mgmtsoc_port_master_internal_port_sink_ready = litespi_tx_mux_endpoint1_sink_ready;
assign litespi_tx_mux_endpoint1_sink_first = mgmtsoc_port_master_internal_port_sink_first;
assign litespi_tx_mux_endpoint1_sink_last = mgmtsoc_port_master_internal_port_sink_last;
assign litespi_tx_mux_endpoint1_sink_payload_data = mgmtsoc_port_master_internal_port_sink_payload_data;
assign litespi_tx_mux_endpoint1_sink_payload_len = mgmtsoc_port_master_internal_port_sink_payload_len;
assign litespi_tx_mux_endpoint1_sink_payload_width = mgmtsoc_port_master_internal_port_sink_payload_width;
assign litespi_tx_mux_endpoint1_sink_payload_mask = mgmtsoc_port_master_internal_port_sink_payload_mask;
assign mgmtsoc_port_master_internal_port_source_valid = litespi_rx_demux_endpoint1_source_valid;
assign litespi_rx_demux_endpoint1_source_ready = mgmtsoc_port_master_internal_port_source_ready;
assign mgmtsoc_port_master_internal_port_source_first = litespi_rx_demux_endpoint1_source_first;
assign mgmtsoc_port_master_internal_port_source_last = litespi_rx_demux_endpoint1_source_last;
assign mgmtsoc_port_master_internal_port_source_payload_data = litespi_rx_demux_endpoint1_source_payload_data;
assign litespi_request = {mgmtsoc_port_master_request, mgmtsoc_port_mmap_request};
assign mgmtsoc_crossbar_source_valid = litespi_tx_mux_source_valid;
assign litespi_tx_mux_source_ready = mgmtsoc_crossbar_source_ready;
assign mgmtsoc_crossbar_source_first = litespi_tx_mux_source_first;
assign mgmtsoc_crossbar_source_last = litespi_tx_mux_source_last;
assign mgmtsoc_crossbar_source_payload_data = litespi_tx_mux_source_payload_data;
assign mgmtsoc_crossbar_source_payload_len = litespi_tx_mux_source_payload_len;
assign mgmtsoc_crossbar_source_payload_width = litespi_tx_mux_source_payload_width;
assign mgmtsoc_crossbar_source_payload_mask = litespi_tx_mux_source_payload_mask;
assign litespi_tx_mux_sel = litespi_grant;
assign litespi_rx_demux_sink_valid = mgmtsoc_crossbar_sink_valid;
assign mgmtsoc_crossbar_sink_ready = litespi_rx_demux_sink_ready;
assign litespi_rx_demux_sink_first = mgmtsoc_crossbar_sink_first;
assign litespi_rx_demux_sink_last = mgmtsoc_crossbar_sink_last;
assign litespi_rx_demux_sink_payload_data = mgmtsoc_crossbar_sink_payload_data;
assign litespi_rx_demux_sel = litespi_grant;
always @(*) begin
	mgmtsoc_crossbar_cs = 1'd0;
	case (litespi_grant)
		1'd0: begin
			mgmtsoc_crossbar_cs = mgmtsoc_litespimmap_cs;
		end
		1'd1: begin
			mgmtsoc_crossbar_cs = mgmtsoc_master_cs;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_source_valid = 1'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_source_valid = litespi_tx_mux_endpoint0_sink_valid;
		end
		1'd1: begin
			litespi_tx_mux_source_valid = litespi_tx_mux_endpoint1_sink_valid;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_endpoint1_sink_ready = 1'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
		end
		1'd1: begin
			litespi_tx_mux_endpoint1_sink_ready = litespi_tx_mux_source_ready;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_source_first = 1'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_source_first = litespi_tx_mux_endpoint0_sink_first;
		end
		1'd1: begin
			litespi_tx_mux_source_first = litespi_tx_mux_endpoint1_sink_first;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_source_last = 1'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_source_last = litespi_tx_mux_endpoint0_sink_last;
		end
		1'd1: begin
			litespi_tx_mux_source_last = litespi_tx_mux_endpoint1_sink_last;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_source_payload_data = 32'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_source_payload_data = litespi_tx_mux_endpoint0_sink_payload_data;
		end
		1'd1: begin
			litespi_tx_mux_source_payload_data = litespi_tx_mux_endpoint1_sink_payload_data;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_source_payload_len = 6'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_source_payload_len = litespi_tx_mux_endpoint0_sink_payload_len;
		end
		1'd1: begin
			litespi_tx_mux_source_payload_len = litespi_tx_mux_endpoint1_sink_payload_len;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_source_payload_width = 4'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_source_payload_width = litespi_tx_mux_endpoint0_sink_payload_width;
		end
		1'd1: begin
			litespi_tx_mux_source_payload_width = litespi_tx_mux_endpoint1_sink_payload_width;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_source_payload_mask = 8'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_source_payload_mask = litespi_tx_mux_endpoint0_sink_payload_mask;
		end
		1'd1: begin
			litespi_tx_mux_source_payload_mask = litespi_tx_mux_endpoint1_sink_payload_mask;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_endpoint0_sink_ready = 1'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_endpoint0_sink_ready = litespi_tx_mux_source_ready;
		end
		1'd1: begin
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_sink_ready = 1'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
			litespi_rx_demux_sink_ready = litespi_rx_demux_endpoint0_source_ready;
		end
		1'd1: begin
			litespi_rx_demux_sink_ready = litespi_rx_demux_endpoint1_source_ready;
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint0_source_valid = 1'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
			litespi_rx_demux_endpoint0_source_valid = litespi_rx_demux_sink_valid;
		end
		1'd1: begin
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint0_source_first = 1'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
			litespi_rx_demux_endpoint0_source_first = litespi_rx_demux_sink_first;
		end
		1'd1: begin
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint0_source_last = 1'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
			litespi_rx_demux_endpoint0_source_last = litespi_rx_demux_sink_last;
		end
		1'd1: begin
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint0_source_payload_data = 32'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
			litespi_rx_demux_endpoint0_source_payload_data = litespi_rx_demux_sink_payload_data;
		end
		1'd1: begin
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint1_source_valid = 1'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
		end
		1'd1: begin
			litespi_rx_demux_endpoint1_source_valid = litespi_rx_demux_sink_valid;
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint1_source_first = 1'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
		end
		1'd1: begin
			litespi_rx_demux_endpoint1_source_first = litespi_rx_demux_sink_first;
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint1_source_last = 1'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
		end
		1'd1: begin
			litespi_rx_demux_endpoint1_source_last = litespi_rx_demux_sink_last;
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint1_source_payload_data = 32'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
		end
		1'd1: begin
			litespi_rx_demux_endpoint1_source_payload_data = litespi_rx_demux_sink_payload_data;
		end
	endcase
end
assign mgmtsoc_litespimmap_spi_dummy_bits = mgmtsoc_litespimmap_storage;
assign mgmtsoc_litespimmap_done = (mgmtsoc_litespimmap_count == 1'd0);
always @(*) begin
	litespi_next_state = 4'd0;
	litespi_next_state = litespi_state;
	case (litespi_state)
		1'd1: begin
			if (mgmtsoc_litespimmap_source_ready) begin
				litespi_next_state = 2'd2;
			end
		end
		2'd2: begin
			if (mgmtsoc_litespimmap_sink_valid) begin
				litespi_next_state = 2'd3;
			end
		end
		2'd3: begin
			if (mgmtsoc_litespimmap_source_ready) begin
				litespi_next_state = 3'd4;
			end
		end
		3'd4: begin
			if (mgmtsoc_litespimmap_sink_valid) begin
				if ((mgmtsoc_litespimmap_spi_dummy_bits == 1'd0)) begin
					litespi_next_state = 3'd7;
				end else begin
					litespi_next_state = 3'd5;
				end
			end
		end
		3'd5: begin
			if (mgmtsoc_litespimmap_source_ready) begin
				litespi_next_state = 3'd6;
			end
		end
		3'd6: begin
			if (mgmtsoc_litespimmap_sink_valid) begin
				litespi_next_state = 3'd7;
			end
		end
		3'd7: begin
			if (mgmtsoc_litespimmap_source_ready) begin
				litespi_next_state = 4'd8;
			end
		end
		4'd8: begin
			if (mgmtsoc_litespimmap_sink_valid) begin
				litespi_next_state = 1'd0;
			end
		end
		default: begin
			if (((mgmtsoc_litespimmap_bus_cyc & mgmtsoc_litespimmap_bus_stb) & (~mgmtsoc_litespimmap_bus_we))) begin
				if ((mgmtsoc_litespimmap_burst_cs & (mgmtsoc_litespimmap_bus_adr == mgmtsoc_litespimmap_burst_adr))) begin
					litespi_next_state = 3'd7;
				end else begin
					litespi_next_state = 1'd1;
				end
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_bus_dat_r = 32'd0;
	case (litespi_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
			mgmtsoc_litespimmap_bus_dat_r = {mgmtsoc_litespimmap_sink_payload_data[7:0], mgmtsoc_litespimmap_sink_payload_data[15:8], mgmtsoc_litespimmap_sink_payload_data[23:16], mgmtsoc_litespimmap_sink_payload_data[31:24]};
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_source_valid = 1'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_source_valid = 1'd1;
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_source_valid = 1'd1;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_source_valid = 1'd1;
		end
		3'd6: begin
		end
		3'd7: begin
			mgmtsoc_litespimmap_source_valid = 1'd1;
		end
		4'd8: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_burst_cs_litespi_next_value0 = 1'd0;
	case (litespi_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_burst_cs_litespi_next_value0 = 1'd1;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_burst_cs_litespi_next_value0 = 1'd1;
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
		end
		default: begin
			mgmtsoc_litespimmap_burst_cs_litespi_next_value0 = (mgmtsoc_litespimmap_burst_cs & (~mgmtsoc_litespimmap_done));
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_burst_cs_litespi_next_value_ce0 = 1'd0;
	case (litespi_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_burst_cs_litespi_next_value_ce0 = 1'd1;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_burst_cs_litespi_next_value_ce0 = 1'd1;
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
		end
		default: begin
			mgmtsoc_litespimmap_burst_cs_litespi_next_value_ce0 = 1'd1;
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_source_last = 1'd0;
	case (litespi_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		3'd7: begin
			mgmtsoc_litespimmap_source_last = 1'd1;
		end
		4'd8: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_bus_ack = 1'd0;
	case (litespi_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
			if (mgmtsoc_litespimmap_sink_valid) begin
				mgmtsoc_litespimmap_bus_ack = 1'd1;
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_source_payload_data = 32'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_source_payload_data = 2'd3;
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_source_payload_data = {mgmtsoc_litespimmap_bus_adr, mgmtsoc_litespimmap};
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_source_payload_data = mgmtsoc_litespimmap_dummy;
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_source_payload_len = 6'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_source_payload_len = 4'd8;
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_source_payload_len = 5'd24;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_source_payload_len = mgmtsoc_litespimmap_spi_dummy_bits;
		end
		3'd6: begin
		end
		3'd7: begin
			mgmtsoc_litespimmap_source_payload_len = 6'd32;
		end
		4'd8: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_source_payload_width = 4'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_source_payload_width = 1'd1;
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_source_payload_width = 1'd1;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_source_payload_width = 1'd1;
		end
		3'd6: begin
		end
		3'd7: begin
			mgmtsoc_litespimmap_source_payload_width = 1'd1;
		end
		4'd8: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_source_payload_mask = 8'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_source_payload_mask = 1'd1;
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_source_payload_mask = 1'd1;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_source_payload_mask = 1'd1;
		end
		3'd6: begin
		end
		3'd7: begin
			mgmtsoc_litespimmap_source_payload_mask = 1'd0;
		end
		4'd8: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_burst_adr_litespi_next_value1 = 30'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_burst_adr_litespi_next_value1 = mgmtsoc_litespimmap_bus_adr;
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_burst_adr_litespi_next_value1 = mgmtsoc_litespimmap_bus_adr;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_burst_adr_litespi_next_value1 = mgmtsoc_litespimmap_bus_adr;
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
			if (mgmtsoc_litespimmap_sink_valid) begin
				mgmtsoc_litespimmap_burst_adr_litespi_next_value1 = (mgmtsoc_litespimmap_burst_adr + 1'd1);
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_cs = 1'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		2'd2: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		2'd3: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		3'd4: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		3'd5: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		3'd6: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		3'd7: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		4'd8: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		default: begin
			mgmtsoc_litespimmap_cs = mgmtsoc_litespimmap_burst_cs;
			if (((mgmtsoc_litespimmap_bus_cyc & mgmtsoc_litespimmap_bus_stb) & (~mgmtsoc_litespimmap_bus_we))) begin
				if ((mgmtsoc_litespimmap_burst_cs & (mgmtsoc_litespimmap_bus_adr == mgmtsoc_litespimmap_burst_adr))) begin
				end else begin
					mgmtsoc_litespimmap_cs = 1'd0;
				end
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_burst_adr_litespi_next_value_ce1 = 1'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_burst_adr_litespi_next_value_ce1 = 1'd1;
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_burst_adr_litespi_next_value_ce1 = 1'd1;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_burst_adr_litespi_next_value_ce1 = 1'd1;
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
			if (mgmtsoc_litespimmap_sink_valid) begin
				mgmtsoc_litespimmap_burst_adr_litespi_next_value_ce1 = 1'd1;
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_sink_ready = 1'd0;
	case (litespi_state)
		1'd1: begin
		end
		2'd2: begin
			mgmtsoc_litespimmap_sink_ready = 1'd1;
		end
		2'd3: begin
		end
		3'd4: begin
			mgmtsoc_litespimmap_sink_ready = 1'd1;
		end
		3'd5: begin
		end
		3'd6: begin
			mgmtsoc_litespimmap_sink_ready = 1'd1;
		end
		3'd7: begin
		end
		4'd8: begin
			mgmtsoc_litespimmap_sink_ready = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_wait = 1'd0;
	case (litespi_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
		end
		default: begin
			mgmtsoc_litespimmap_wait = 1'd1;
		end
	endcase
end
assign mgmtsoc_master_rx_fifo_sink_valid = mgmtsoc_master_sink_sink_valid;
assign mgmtsoc_master_sink_sink_ready = mgmtsoc_master_rx_fifo_sink_ready;
assign mgmtsoc_master_rx_fifo_sink_first = mgmtsoc_master_sink_sink_first;
assign mgmtsoc_master_rx_fifo_sink_last = mgmtsoc_master_sink_sink_last;
assign mgmtsoc_master_rx_fifo_sink_payload_data = mgmtsoc_master_sink_sink_payload_data;
assign mgmtsoc_master_source_source_valid = mgmtsoc_master_tx_fifo_source_valid;
assign mgmtsoc_master_tx_fifo_source_ready = mgmtsoc_master_source_source_ready;
assign mgmtsoc_master_source_source_first = mgmtsoc_master_tx_fifo_source_first;
assign mgmtsoc_master_source_source_last = mgmtsoc_master_tx_fifo_source_last;
assign mgmtsoc_master_source_source_payload_data = mgmtsoc_master_tx_fifo_source_payload_data;
assign mgmtsoc_master_source_source_payload_len = mgmtsoc_master_tx_fifo_source_payload_len;
assign mgmtsoc_master_source_source_payload_width = mgmtsoc_master_tx_fifo_source_payload_width;
assign mgmtsoc_master_source_source_payload_mask = mgmtsoc_master_tx_fifo_source_payload_mask;
assign mgmtsoc_master_cs = mgmtsoc_master_cs_storage;
assign mgmtsoc_master_tx_fifo_sink_valid = mgmtsoc_master_rxtx_re;
assign mgmtsoc_master_tx_ready = mgmtsoc_master_tx_fifo_sink_ready;
assign mgmtsoc_master_tx_fifo_sink_payload_data = mgmtsoc_master_rxtx_r;
assign mgmtsoc_master_tx_fifo_sink_payload_len = mgmtsoc_master_len;
assign mgmtsoc_master_tx_fifo_sink_payload_width = mgmtsoc_master_width;
assign mgmtsoc_master_tx_fifo_sink_payload_mask = mgmtsoc_master_mask;
assign mgmtsoc_master_tx_fifo_sink_last = 1'd1;
assign mgmtsoc_master_rx_fifo_source_ready = mgmtsoc_master_rxtx_we;
assign mgmtsoc_master_rx_ready = mgmtsoc_master_rx_fifo_source_valid;
assign mgmtsoc_master_rxtx_w = mgmtsoc_master_rx_fifo_source_payload_data;
assign mgmtsoc_master_tx_fifo_sink_ready = ((~mgmtsoc_master_tx_fifo_source_valid) | mgmtsoc_master_tx_fifo_source_ready);
assign mgmtsoc_master_rx_fifo_sink_ready = ((~mgmtsoc_master_rx_fifo_source_valid) | mgmtsoc_master_rx_fifo_source_ready);
assign spi_master_start0 = spi_master_start1;
assign spi_master_length0 = spi_master_length1;
assign spi_master_done1 = spi_master_done0;
assign spi_master_mosi = spi_master_mosi_storage;
assign spi_master_miso_status = spi_master_miso;
assign spi_master_cs = spi_master_sel;
assign spi_master_cs_mode = spi_master_mode0;
assign spi_master_loopback = spi_master_mode1;
assign spi_master_clk_rise = (spi_master_clk_divider1 == (spi_master_clk_divider0[15:1] - 1'd1));
assign spi_master_clk_fall = (spi_master_clk_divider1 == (spi_master_clk_divider0 - 1'd1));
assign spi_master_clk_divider0 = spimaster_storage;
always @(*) begin
	spimaster_next_state = 2'd0;
	spimaster_next_state = spimaster_state;
	case (spimaster_state)
		1'd1: begin
			if (spi_master_clk_fall) begin
				spimaster_next_state = 2'd2;
			end
		end
		2'd2: begin
			if (spi_master_clk_fall) begin
				if ((spi_master_count == (spi_master_length0 - 1'd1))) begin
					spimaster_next_state = 2'd3;
				end
			end
		end
		2'd3: begin
			if (spi_master_clk_rise) begin
				spimaster_next_state = 1'd0;
			end
		end
		default: begin
			if (spi_master_start0) begin
				spimaster_next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	spi_master_count_spimaster_next_value = 3'd0;
	case (spimaster_state)
		1'd1: begin
			spi_master_count_spimaster_next_value = 1'd0;
		end
		2'd2: begin
			if (spi_master_clk_fall) begin
				spi_master_count_spimaster_next_value = (spi_master_count + 1'd1);
			end
		end
		2'd3: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	spi_master_done0 = 1'd0;
	case (spimaster_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		default: begin
			spi_master_done0 = 1'd1;
			if (spi_master_start0) begin
				spi_master_done0 = 1'd0;
			end
		end
	endcase
end
always @(*) begin
	spi_master_count_spimaster_next_value_ce = 1'd0;
	case (spimaster_state)
		1'd1: begin
			spi_master_count_spimaster_next_value_ce = 1'd1;
		end
		2'd2: begin
			if (spi_master_clk_fall) begin
				spi_master_count_spimaster_next_value_ce = 1'd1;
			end
		end
		2'd3: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	spi_master_irq = 1'd0;
	case (spimaster_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			if (spi_master_clk_rise) begin
				spi_master_irq = 1'd1;
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	spi_master_clk_enable = 1'd0;
	case (spimaster_state)
		1'd1: begin
		end
		2'd2: begin
			spi_master_clk_enable = 1'd1;
		end
		2'd3: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	spi_master_xfer_enable = 1'd0;
	case (spimaster_state)
		1'd1: begin
			if (spi_master_clk_fall) begin
				spi_master_xfer_enable = 1'd1;
			end
		end
		2'd2: begin
			spi_master_xfer_enable = 1'd1;
		end
		2'd3: begin
			spi_master_xfer_enable = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	spi_master_mosi_latch = 1'd0;
	case (spimaster_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		default: begin
			if (spi_master_start0) begin
				spi_master_mosi_latch = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	spi_master_miso_latch = 1'd0;
	case (spimaster_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			if (spi_master_clk_rise) begin
				spi_master_miso_latch = 1'd1;
			end
		end
		default: begin
		end
	endcase
end
assign mprj_wb_iena = mprj_wb_iena_storage;
always @(*) begin
	rs232phy_rs232phytx_next_state = 1'd0;
	rs232phy_rs232phytx_next_state = rs232phy_rs232phytx_state;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				if ((uart_phy_tx_count == 4'd9)) begin
					rs232phy_rs232phytx_next_state = 1'd0;
				end
			end
		end
		default: begin
			if (uart_phy_tx_sink_valid) begin
				rs232phy_rs232phytx_next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	sys_uart_tx_rs232phy_rs232phytx_next_value_ce1 = 1'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				sys_uart_tx_rs232phy_rs232phytx_next_value_ce1 = 1'd1;
			end
		end
		default: begin
			sys_uart_tx_rs232phy_rs232phytx_next_value_ce1 = 1'd1;
			if (uart_phy_tx_sink_valid) begin
				sys_uart_tx_rs232phy_rs232phytx_next_value_ce1 = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	uart_phy_tx_data_rs232phy_rs232phytx_next_value2 = 8'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				uart_phy_tx_data_rs232phy_rs232phytx_next_value2 = {1'd1, uart_phy_tx_data[7:1]};
			end
		end
		default: begin
			if (uart_phy_tx_sink_valid) begin
				uart_phy_tx_data_rs232phy_rs232phytx_next_value2 = uart_phy_tx_sink_payload_data;
			end
		end
	endcase
end
always @(*) begin
	uart_phy_tx_sink_ready = 1'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				if ((uart_phy_tx_count == 4'd9)) begin
					uart_phy_tx_sink_ready = 1'd1;
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	uart_phy_tx_data_rs232phy_rs232phytx_next_value_ce2 = 1'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				uart_phy_tx_data_rs232phy_rs232phytx_next_value_ce2 = 1'd1;
			end
		end
		default: begin
			if (uart_phy_tx_sink_valid) begin
				uart_phy_tx_data_rs232phy_rs232phytx_next_value_ce2 = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	uart_phy_tx_enable = 1'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			uart_phy_tx_enable = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	uart_phy_tx_count_rs232phy_rs232phytx_next_value0 = 4'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				uart_phy_tx_count_rs232phy_rs232phytx_next_value0 = (uart_phy_tx_count + 1'd1);
			end
		end
		default: begin
			uart_phy_tx_count_rs232phy_rs232phytx_next_value0 = 1'd0;
		end
	endcase
end
always @(*) begin
	uart_phy_tx_count_rs232phy_rs232phytx_next_value_ce0 = 1'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				uart_phy_tx_count_rs232phy_rs232phytx_next_value_ce0 = 1'd1;
			end
		end
		default: begin
			uart_phy_tx_count_rs232phy_rs232phytx_next_value_ce0 = 1'd1;
		end
	endcase
end
always @(*) begin
	sys_uart_tx_rs232phy_rs232phytx_next_value1 = 1'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				sys_uart_tx_rs232phy_rs232phytx_next_value1 = uart_phy_tx_data;
			end
		end
		default: begin
			sys_uart_tx_rs232phy_rs232phytx_next_value1 = 1'd1;
			if (uart_phy_tx_sink_valid) begin
				sys_uart_tx_rs232phy_rs232phytx_next_value1 = 1'd0;
			end
		end
	endcase
end
always @(*) begin
	rs232phy_rs232phyrx_next_state = 1'd0;
	rs232phy_rs232phyrx_next_state = rs232phy_rs232phyrx_state;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			if (uart_phy_rx_tick) begin
				if ((uart_phy_rx_count == 4'd9)) begin
					rs232phy_rs232phyrx_next_state = 1'd0;
				end
			end
		end
		default: begin
			if (((uart_phy_rx_rx == 1'd0) & (uart_phy_rx_rx_d == 1'd1))) begin
				rs232phy_rs232phyrx_next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	uart_phy_rx_data_rs232phy_rs232phyrx_next_value1 = 8'd0;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			if (uart_phy_rx_tick) begin
				uart_phy_rx_data_rs232phy_rs232phyrx_next_value1 = {uart_phy_rx_rx, uart_phy_rx_data[7:1]};
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	uart_phy_rx_data_rs232phy_rs232phyrx_next_value_ce1 = 1'd0;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			if (uart_phy_rx_tick) begin
				uart_phy_rx_data_rs232phy_rs232phyrx_next_value_ce1 = 1'd1;
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	uart_phy_rx_source_valid = 1'd0;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			if (uart_phy_rx_tick) begin
				if ((uart_phy_rx_count == 4'd9)) begin
					uart_phy_rx_source_valid = (uart_phy_rx_rx == 1'd1);
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	uart_phy_rx_source_payload_data = 8'd0;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			if (uart_phy_rx_tick) begin
				if ((uart_phy_rx_count == 4'd9)) begin
					uart_phy_rx_source_payload_data = uart_phy_rx_data;
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	uart_phy_rx_enable = 1'd0;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			uart_phy_rx_enable = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	uart_phy_rx_count_rs232phy_rs232phyrx_next_value0 = 4'd0;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			if (uart_phy_rx_tick) begin
				uart_phy_rx_count_rs232phy_rs232phyrx_next_value0 = (uart_phy_rx_count + 1'd1);
			end
		end
		default: begin
			uart_phy_rx_count_rs232phy_rs232phyrx_next_value0 = 1'd0;
		end
	endcase
end
always @(*) begin
	uart_phy_rx_count_rs232phy_rs232phyrx_next_value_ce0 = 1'd0;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			if (uart_phy_rx_tick) begin
				uart_phy_rx_count_rs232phy_rs232phyrx_next_value_ce0 = 1'd1;
			end
		end
		default: begin
			uart_phy_rx_count_rs232phy_rs232phyrx_next_value_ce0 = 1'd1;
		end
	endcase
end
assign uart_uart_sink_valid = uart_phy_rx_source_valid;
assign uart_phy_rx_source_ready = uart_uart_sink_ready;
assign uart_uart_sink_first = uart_phy_rx_source_first;
assign uart_uart_sink_last = uart_phy_rx_source_last;
assign uart_uart_sink_payload_data = uart_phy_rx_source_payload_data;
assign uart_phy_tx_sink_valid = uart_uart_source_valid;
assign uart_uart_source_ready = uart_phy_tx_sink_ready;
assign uart_phy_tx_sink_first = uart_uart_source_first;
assign uart_phy_tx_sink_last = uart_uart_source_last;
assign uart_phy_tx_sink_payload_data = uart_uart_source_payload_data;
assign uart_tx_fifo_sink_valid = uart_rxtx_re;
assign uart_tx_fifo_sink_payload_data = uart_rxtx_r;
assign uart_uart_source_valid = uart_tx_fifo_source_valid;
assign uart_tx_fifo_source_ready = uart_uart_source_ready;
assign uart_uart_source_first = uart_tx_fifo_source_first;
assign uart_uart_source_last = uart_tx_fifo_source_last;
assign uart_uart_source_payload_data = uart_tx_fifo_source_payload_data;
assign uart_txfull_status = (~uart_tx_fifo_sink_ready);
assign uart_txempty_status = (~uart_tx_fifo_source_valid);
assign uart_tx_trigger = uart_tx_fifo_sink_ready;
assign uart_rx_fifo_sink_valid = uart_uart_sink_valid;
assign uart_uart_sink_ready = uart_rx_fifo_sink_ready;
assign uart_rx_fifo_sink_first = uart_uart_sink_first;
assign uart_rx_fifo_sink_last = uart_uart_sink_last;
assign uart_rx_fifo_sink_payload_data = uart_uart_sink_payload_data;
assign uart_rxtx_w = uart_rx_fifo_source_payload_data;
assign uart_rx_fifo_source_ready = (uart_rx_clear | (1'd0 & uart_rxtx_we));
assign uart_rxempty_status = (~uart_rx_fifo_source_valid);
assign uart_rxfull_status = (~uart_rx_fifo_sink_ready);
assign uart_rx_trigger = uart_rx_fifo_source_valid;
assign uart_tx0 = uart_tx_status;
assign uart_tx1 = uart_tx_pending;
always @(*) begin
	uart_tx_clear = 1'd0;
	if ((uart_pending_re & uart_pending_r[0])) begin
		uart_tx_clear = 1'd1;
	end
end
assign uart_rx0 = uart_rx_status;
assign uart_rx1 = uart_rx_pending;
always @(*) begin
	uart_rx_clear = 1'd0;
	if ((uart_pending_re & uart_pending_r[1])) begin
		uart_rx_clear = 1'd1;
	end
end
assign uart_irq = ((uart_pending_status[0] & uart_enable_storage[0]) | (uart_pending_status[1] & uart_enable_storage[1]));
assign uart_tx_status = uart_tx_trigger;
assign uart_rx_status = uart_rx_trigger;
assign uart_tx_fifo_syncfifo_din = {uart_tx_fifo_fifo_in_last, uart_tx_fifo_fifo_in_first, uart_tx_fifo_fifo_in_payload_data};
assign {uart_tx_fifo_fifo_out_last, uart_tx_fifo_fifo_out_first, uart_tx_fifo_fifo_out_payload_data} = uart_tx_fifo_syncfifo_dout;
assign uart_tx_fifo_sink_ready = uart_tx_fifo_syncfifo_writable;
assign uart_tx_fifo_syncfifo_we = uart_tx_fifo_sink_valid;
assign uart_tx_fifo_fifo_in_first = uart_tx_fifo_sink_first;
assign uart_tx_fifo_fifo_in_last = uart_tx_fifo_sink_last;
assign uart_tx_fifo_fifo_in_payload_data = uart_tx_fifo_sink_payload_data;
assign uart_tx_fifo_source_valid = uart_tx_fifo_readable;
assign uart_tx_fifo_source_first = uart_tx_fifo_fifo_out_first;
assign uart_tx_fifo_source_last = uart_tx_fifo_fifo_out_last;
assign uart_tx_fifo_source_payload_data = uart_tx_fifo_fifo_out_payload_data;
assign uart_tx_fifo_re = uart_tx_fifo_source_ready;
assign uart_tx_fifo_syncfifo_re = (uart_tx_fifo_syncfifo_readable & ((~uart_tx_fifo_readable) | uart_tx_fifo_re));
assign uart_tx_fifo_level1 = (uart_tx_fifo_level0 + uart_tx_fifo_readable);
always @(*) begin
	uart_tx_fifo_wrport_adr = 4'd0;
	if (uart_tx_fifo_replace) begin
		uart_tx_fifo_wrport_adr = (uart_tx_fifo_produce - 1'd1);
	end else begin
		uart_tx_fifo_wrport_adr = uart_tx_fifo_produce;
	end
end
assign uart_tx_fifo_wrport_dat_w = uart_tx_fifo_syncfifo_din;
assign uart_tx_fifo_wrport_we = (uart_tx_fifo_syncfifo_we & (uart_tx_fifo_syncfifo_writable | uart_tx_fifo_replace));
assign uart_tx_fifo_do_read = (uart_tx_fifo_syncfifo_readable & uart_tx_fifo_syncfifo_re);
assign uart_tx_fifo_rdport_adr = uart_tx_fifo_consume;
assign uart_tx_fifo_syncfifo_dout = uart_tx_fifo_rdport_dat_r;
assign uart_tx_fifo_rdport_re = uart_tx_fifo_do_read;
assign uart_tx_fifo_syncfifo_writable = (uart_tx_fifo_level0 != 5'd16);
assign uart_tx_fifo_syncfifo_readable = (uart_tx_fifo_level0 != 1'd0);
assign uart_rx_fifo_syncfifo_din = {uart_rx_fifo_fifo_in_last, uart_rx_fifo_fifo_in_first, uart_rx_fifo_fifo_in_payload_data};
assign {uart_rx_fifo_fifo_out_last, uart_rx_fifo_fifo_out_first, uart_rx_fifo_fifo_out_payload_data} = uart_rx_fifo_syncfifo_dout;
assign uart_rx_fifo_sink_ready = uart_rx_fifo_syncfifo_writable;
assign uart_rx_fifo_syncfifo_we = uart_rx_fifo_sink_valid;
assign uart_rx_fifo_fifo_in_first = uart_rx_fifo_sink_first;
assign uart_rx_fifo_fifo_in_last = uart_rx_fifo_sink_last;
assign uart_rx_fifo_fifo_in_payload_data = uart_rx_fifo_sink_payload_data;
assign uart_rx_fifo_source_valid = uart_rx_fifo_readable;
assign uart_rx_fifo_source_first = uart_rx_fifo_fifo_out_first;
assign uart_rx_fifo_source_last = uart_rx_fifo_fifo_out_last;
assign uart_rx_fifo_source_payload_data = uart_rx_fifo_fifo_out_payload_data;
assign uart_rx_fifo_re = uart_rx_fifo_source_ready;
assign uart_rx_fifo_syncfifo_re = (uart_rx_fifo_syncfifo_readable & ((~uart_rx_fifo_readable) | uart_rx_fifo_re));
assign uart_rx_fifo_level1 = (uart_rx_fifo_level0 + uart_rx_fifo_readable);
always @(*) begin
	uart_rx_fifo_wrport_adr = 4'd0;
	if (uart_rx_fifo_replace) begin
		uart_rx_fifo_wrport_adr = (uart_rx_fifo_produce - 1'd1);
	end else begin
		uart_rx_fifo_wrport_adr = uart_rx_fifo_produce;
	end
end
assign uart_rx_fifo_wrport_dat_w = uart_rx_fifo_syncfifo_din;
assign uart_rx_fifo_wrport_we = (uart_rx_fifo_syncfifo_we & (uart_rx_fifo_syncfifo_writable | uart_rx_fifo_replace));
assign uart_rx_fifo_do_read = (uart_rx_fifo_syncfifo_readable & uart_rx_fifo_syncfifo_re);
assign uart_rx_fifo_rdport_adr = uart_rx_fifo_consume;
assign uart_rx_fifo_syncfifo_dout = uart_rx_fifo_rdport_dat_r;
assign uart_rx_fifo_rdport_re = uart_rx_fifo_do_read;
assign uart_rx_fifo_syncfifo_writable = (uart_rx_fifo_level0 != 5'd16);
assign uart_rx_fifo_syncfifo_readable = (uart_rx_fifo_level0 != 1'd0);
assign dbg_uart_wait = (~dbg_uart_is_ongoing);
assign dbg_uart_reset = dbg_uart_done;
assign dbg_uart_wishbone_adr = dbg_uart_address;
assign dbg_uart_wishbone_dat_w = dbg_uart_data;
assign dbg_uart_wishbone_sel = 4'd15;
always @(*) begin
	dbg_uart_tx_sink_payload_data = 8'd0;
	case (dbg_uart_bytes_count)
		1'd0: begin
			dbg_uart_tx_sink_payload_data = dbg_uart_data[31:24];
		end
		1'd1: begin
			dbg_uart_tx_sink_payload_data = dbg_uart_data[31:16];
		end
		2'd2: begin
			dbg_uart_tx_sink_payload_data = dbg_uart_data[31:8];
		end
		2'd3: begin
			dbg_uart_tx_sink_payload_data = dbg_uart_data[31:0];
		end
	endcase
end
assign dbg_uart_tx_sink_last = ((dbg_uart_bytes_count == 2'd3) & (dbg_uart_words_count == (dbg_uart_length - 1'd1)));
always @(*) begin
	uartwishbonebridge_rs232phytx_next_state = 1'd0;
	uartwishbonebridge_rs232phytx_next_state = uartwishbonebridge_rs232phytx_state;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				if ((dbg_uart_tx_count == 4'd9)) begin
					uartwishbonebridge_rs232phytx_next_state = 1'd0;
				end
			end
		end
		default: begin
			if (dbg_uart_tx_sink_valid) begin
				uartwishbonebridge_rs232phytx_next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_tx_sink_ready = 1'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				if ((dbg_uart_tx_count == 4'd9)) begin
					dbg_uart_tx_sink_ready = 1'd1;
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value2 = 8'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value2 = {1'd1, dbg_uart_tx_data[7:1]};
			end
		end
		default: begin
			if (dbg_uart_tx_sink_valid) begin
				dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value2 = dbg_uart_tx_sink_payload_data;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value_ce2 = 1'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value_ce2 = 1'd1;
			end
		end
		default: begin
			if (dbg_uart_tx_sink_valid) begin
				dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value_ce2 = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_tx_enable = 1'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			dbg_uart_tx_enable = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value0 = 4'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value0 = (dbg_uart_tx_count + 1'd1);
			end
		end
		default: begin
			dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value0 = 1'd0;
		end
	endcase
end
always @(*) begin
	dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value_ce0 = 1'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value_ce0 = 1'd1;
			end
		end
		default: begin
			dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value_ce0 = 1'd1;
		end
	endcase
end
always @(*) begin
	dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value1 = 1'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value1 = dbg_uart_tx_data;
			end
		end
		default: begin
			dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value1 = 1'd1;
			if (dbg_uart_tx_sink_valid) begin
				dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value1 = 1'd0;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value_ce1 = 1'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value_ce1 = 1'd1;
			end
		end
		default: begin
			dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value_ce1 = 1'd1;
			if (dbg_uart_tx_sink_valid) begin
				dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value_ce1 = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	uartwishbonebridge_rs232phyrx_next_state = 1'd0;
	uartwishbonebridge_rs232phyrx_next_state = uartwishbonebridge_rs232phyrx_state;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			if (dbg_uart_rx_tick) begin
				if ((dbg_uart_rx_count == 4'd9)) begin
					uartwishbonebridge_rs232phyrx_next_state = 1'd0;
				end
			end
		end
		default: begin
			if (((dbg_uart_rx_rx == 1'd0) & (dbg_uart_rx_rx_d == 1'd1))) begin
				uartwishbonebridge_rs232phyrx_next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_source_valid = 1'd0;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			if (dbg_uart_rx_tick) begin
				if ((dbg_uart_rx_count == 4'd9)) begin
					dbg_uart_rx_source_valid = (dbg_uart_rx_rx == 1'd1);
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value1 = 8'd0;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			if (dbg_uart_rx_tick) begin
				dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value1 = {dbg_uart_rx_rx, dbg_uart_rx_data[7:1]};
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value_ce1 = 1'd0;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			if (dbg_uart_rx_tick) begin
				dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value_ce1 = 1'd1;
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_source_payload_data = 8'd0;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			if (dbg_uart_rx_tick) begin
				if ((dbg_uart_rx_count == 4'd9)) begin
					dbg_uart_rx_source_payload_data = dbg_uart_rx_data;
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_enable = 1'd0;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			dbg_uart_rx_enable = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value0 = 4'd0;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			if (dbg_uart_rx_tick) begin
				dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value0 = (dbg_uart_rx_count + 1'd1);
			end
		end
		default: begin
			dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value0 = 1'd0;
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value_ce0 = 1'd0;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			if (dbg_uart_rx_tick) begin
				dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value_ce0 = 1'd1;
			end
		end
		default: begin
			dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value_ce0 = 1'd1;
		end
	endcase
end
always @(*) begin
	uartwishbonebridge_next_state = 3'd0;
	uartwishbonebridge_next_state = uartwishbonebridge_state;
	case (uartwishbonebridge_state)
		1'd1: begin
			if (dbg_uart_rx_source_valid) begin
				uartwishbonebridge_next_state = 2'd2;
			end
		end
		2'd2: begin
			if (dbg_uart_rx_source_valid) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					if (((dbg_uart_cmd == 1'd1) | (dbg_uart_cmd == 2'd3))) begin
						uartwishbonebridge_next_state = 2'd3;
					end else begin
						if (((dbg_uart_cmd == 2'd2) | (dbg_uart_cmd == 3'd4))) begin
							uartwishbonebridge_next_state = 3'd5;
						end else begin
							uartwishbonebridge_next_state = 1'd0;
						end
					end
				end
			end
		end
		2'd3: begin
			if (dbg_uart_rx_source_valid) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					uartwishbonebridge_next_state = 3'd4;
				end
			end
		end
		3'd4: begin
			if (dbg_uart_wishbone_ack) begin
				if ((dbg_uart_words_count == (dbg_uart_length - 1'd1))) begin
					uartwishbonebridge_next_state = 1'd0;
				end else begin
					uartwishbonebridge_next_state = 2'd3;
				end
			end
		end
		3'd5: begin
			if (dbg_uart_wishbone_ack) begin
				uartwishbonebridge_next_state = 3'd6;
			end
		end
		3'd6: begin
			if (dbg_uart_tx_sink_ready) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					if ((dbg_uart_words_count == (dbg_uart_length - 1'd1))) begin
						uartwishbonebridge_next_state = 1'd0;
					end else begin
						uartwishbonebridge_next_state = 3'd5;
					end
				end
			end
		end
		default: begin
			if (dbg_uart_rx_source_valid) begin
				uartwishbonebridge_next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_bytes_count_uartwishbonebridge_next_value0 = 2'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_bytes_count_uartwishbonebridge_next_value0 = (dbg_uart_bytes_count + 1'd1);
			end
		end
		2'd3: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_bytes_count_uartwishbonebridge_next_value0 = (dbg_uart_bytes_count + 1'd1);
			end
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
			if (dbg_uart_tx_sink_ready) begin
				dbg_uart_bytes_count_uartwishbonebridge_next_value0 = (dbg_uart_bytes_count + 1'd1);
			end
		end
		default: begin
			dbg_uart_bytes_count_uartwishbonebridge_next_value0 = 1'd0;
		end
	endcase
end
always @(*) begin
	dbg_uart_bytes_count_uartwishbonebridge_next_value_ce0 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_bytes_count_uartwishbonebridge_next_value_ce0 = 1'd1;
			end
		end
		2'd3: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_bytes_count_uartwishbonebridge_next_value_ce0 = 1'd1;
			end
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
			if (dbg_uart_tx_sink_ready) begin
				dbg_uart_bytes_count_uartwishbonebridge_next_value_ce0 = 1'd1;
			end
		end
		default: begin
			dbg_uart_bytes_count_uartwishbonebridge_next_value_ce0 = 1'd1;
		end
	endcase
end
always @(*) begin
	dbg_uart_wishbone_cyc = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
			dbg_uart_wishbone_cyc = 1'd1;
		end
		3'd5: begin
			dbg_uart_wishbone_cyc = 1'd1;
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_wishbone_stb = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
			dbg_uart_wishbone_stb = 1'd1;
		end
		3'd5: begin
			dbg_uart_wishbone_stb = 1'd1;
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_words_count_uartwishbonebridge_next_value1 = 8'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
			if (dbg_uart_wishbone_ack) begin
				dbg_uart_words_count_uartwishbonebridge_next_value1 = (dbg_uart_words_count + 1'd1);
			end
		end
		3'd5: begin
		end
		3'd6: begin
			if (dbg_uart_tx_sink_ready) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					dbg_uart_words_count_uartwishbonebridge_next_value1 = (dbg_uart_words_count + 1'd1);
				end
			end
		end
		default: begin
			dbg_uart_words_count_uartwishbonebridge_next_value1 = 1'd0;
		end
	endcase
end
always @(*) begin
	dbg_uart_wishbone_we = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
			dbg_uart_wishbone_we = 1'd1;
		end
		3'd5: begin
			dbg_uart_wishbone_we = 1'd0;
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_words_count_uartwishbonebridge_next_value_ce1 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
			if (dbg_uart_wishbone_ack) begin
				dbg_uart_words_count_uartwishbonebridge_next_value_ce1 = 1'd1;
			end
		end
		3'd5: begin
		end
		3'd6: begin
			if (dbg_uart_tx_sink_ready) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					dbg_uart_words_count_uartwishbonebridge_next_value_ce1 = 1'd1;
				end
			end
		end
		default: begin
			dbg_uart_words_count_uartwishbonebridge_next_value_ce1 = 1'd1;
		end
	endcase
end
always @(*) begin
	dbg_uart_cmd_uartwishbonebridge_next_value2 = 8'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		default: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_cmd_uartwishbonebridge_next_value2 = dbg_uart_rx_source_payload_data;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_cmd_uartwishbonebridge_next_value_ce2 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		default: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_cmd_uartwishbonebridge_next_value_ce2 = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_length_uartwishbonebridge_next_value3 = 8'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_length_uartwishbonebridge_next_value3 = dbg_uart_rx_source_payload_data;
			end
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_length_uartwishbonebridge_next_value_ce3 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_length_uartwishbonebridge_next_value_ce3 = 1'd1;
			end
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_address_uartwishbonebridge_next_value4 = 32'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_address_uartwishbonebridge_next_value4 = {dbg_uart_address, dbg_uart_rx_source_payload_data};
			end
		end
		2'd3: begin
		end
		3'd4: begin
			if (dbg_uart_wishbone_ack) begin
				dbg_uart_address_uartwishbonebridge_next_value4 = (dbg_uart_address + dbg_uart_incr);
			end
		end
		3'd5: begin
		end
		3'd6: begin
			if (dbg_uart_tx_sink_ready) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					dbg_uart_address_uartwishbonebridge_next_value4 = (dbg_uart_address + dbg_uart_incr);
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_address_uartwishbonebridge_next_value_ce4 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_address_uartwishbonebridge_next_value_ce4 = 1'd1;
			end
		end
		2'd3: begin
		end
		3'd4: begin
			if (dbg_uart_wishbone_ack) begin
				dbg_uart_address_uartwishbonebridge_next_value_ce4 = 1'd1;
			end
		end
		3'd5: begin
		end
		3'd6: begin
			if (dbg_uart_tx_sink_ready) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					dbg_uart_address_uartwishbonebridge_next_value_ce4 = 1'd1;
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_incr_uartwishbonebridge_next_value5 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
			if (dbg_uart_rx_source_valid) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					if (((dbg_uart_cmd == 1'd1) | (dbg_uart_cmd == 2'd3))) begin
						dbg_uart_incr_uartwishbonebridge_next_value5 = (dbg_uart_cmd == 1'd1);
					end else begin
						if (((dbg_uart_cmd == 2'd2) | (dbg_uart_cmd == 3'd4))) begin
							dbg_uart_incr_uartwishbonebridge_next_value5 = (dbg_uart_cmd == 2'd2);
						end else begin
						end
					end
				end
			end
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_incr_uartwishbonebridge_next_value_ce5 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
			if (dbg_uart_rx_source_valid) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					if (((dbg_uart_cmd == 1'd1) | (dbg_uart_cmd == 2'd3))) begin
						dbg_uart_incr_uartwishbonebridge_next_value_ce5 = 1'd1;
					end else begin
						if (((dbg_uart_cmd == 2'd2) | (dbg_uart_cmd == 3'd4))) begin
							dbg_uart_incr_uartwishbonebridge_next_value_ce5 = 1'd1;
						end else begin
						end
					end
				end
			end
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_tx_sink_valid = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
			dbg_uart_tx_sink_valid = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_data_uartwishbonebridge_next_value6 = 32'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_data_uartwishbonebridge_next_value6 = {dbg_uart_data, dbg_uart_rx_source_payload_data};
			end
		end
		3'd4: begin
		end
		3'd5: begin
			if (dbg_uart_wishbone_ack) begin
				dbg_uart_data_uartwishbonebridge_next_value6 = dbg_uart_wishbone_dat_r;
			end
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_is_ongoing = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		default: begin
			dbg_uart_is_ongoing = 1'd1;
		end
	endcase
end
always @(*) begin
	dbg_uart_data_uartwishbonebridge_next_value_ce6 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_data_uartwishbonebridge_next_value_ce6 = 1'd1;
			end
		end
		3'd4: begin
		end
		3'd5: begin
			if (dbg_uart_wishbone_ack) begin
				dbg_uart_data_uartwishbonebridge_next_value_ce6 = 1'd1;
			end
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_source_ready = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
			dbg_uart_rx_source_ready = 1'd1;
		end
		2'd2: begin
			dbg_uart_rx_source_ready = 1'd1;
		end
		2'd3: begin
			dbg_uart_rx_source_ready = 1'd1;
		end
		3'd4: begin
			dbg_uart_rx_source_ready = 1'd0;
		end
		3'd5: begin
			dbg_uart_rx_source_ready = 1'd0;
		end
		3'd6: begin
			dbg_uart_rx_source_ready = 1'd0;
		end
		default: begin
			dbg_uart_rx_source_ready = 1'd1;
		end
	endcase
end
assign dbg_uart_done = (dbg_uart_count == 1'd0);
assign debug_oeb = debug_oeb_storage;
assign debug_mode = debug_mode_storage;
assign uart_enabled_o = uart_enabled_storage;
assign gpio_mode0_pad = gpio_mode0_storage;
assign gpio_mode1_pad = gpio_mode1_storage;
assign gpio_inenb_pad = (~gpio_ien_storage);
assign gpio_outenb_pad = (~gpio_oe_storage);
assign gpio_out_pad = gpio_out_storage;
always @(*) begin
	la_iena = 128'd0;
	la_iena[0] = (~la_ien_storage[0]);
	la_iena[1] = (~la_ien_storage[1]);
	la_iena[2] = (~la_ien_storage[2]);
	la_iena[3] = (~la_ien_storage[3]);
	la_iena[4] = (~la_ien_storage[4]);
	la_iena[5] = (~la_ien_storage[5]);
	la_iena[6] = (~la_ien_storage[6]);
	la_iena[7] = (~la_ien_storage[7]);
	la_iena[8] = (~la_ien_storage[8]);
	la_iena[9] = (~la_ien_storage[9]);
	la_iena[10] = (~la_ien_storage[10]);
	la_iena[11] = (~la_ien_storage[11]);
	la_iena[12] = (~la_ien_storage[12]);
	la_iena[13] = (~la_ien_storage[13]);
	la_iena[14] = (~la_ien_storage[14]);
	la_iena[15] = (~la_ien_storage[15]);
	la_iena[16] = (~la_ien_storage[16]);
	la_iena[17] = (~la_ien_storage[17]);
	la_iena[18] = (~la_ien_storage[18]);
	la_iena[19] = (~la_ien_storage[19]);
	la_iena[20] = (~la_ien_storage[20]);
	la_iena[21] = (~la_ien_storage[21]);
	la_iena[22] = (~la_ien_storage[22]);
	la_iena[23] = (~la_ien_storage[23]);
	la_iena[24] = (~la_ien_storage[24]);
	la_iena[25] = (~la_ien_storage[25]);
	la_iena[26] = (~la_ien_storage[26]);
	la_iena[27] = (~la_ien_storage[27]);
	la_iena[28] = (~la_ien_storage[28]);
	la_iena[29] = (~la_ien_storage[29]);
	la_iena[30] = (~la_ien_storage[30]);
	la_iena[31] = (~la_ien_storage[31]);
	la_iena[32] = (~la_ien_storage[32]);
	la_iena[33] = (~la_ien_storage[33]);
	la_iena[34] = (~la_ien_storage[34]);
	la_iena[35] = (~la_ien_storage[35]);
	la_iena[36] = (~la_ien_storage[36]);
	la_iena[37] = (~la_ien_storage[37]);
	la_iena[38] = (~la_ien_storage[38]);
	la_iena[39] = (~la_ien_storage[39]);
	la_iena[40] = (~la_ien_storage[40]);
	la_iena[41] = (~la_ien_storage[41]);
	la_iena[42] = (~la_ien_storage[42]);
	la_iena[43] = (~la_ien_storage[43]);
	la_iena[44] = (~la_ien_storage[44]);
	la_iena[45] = (~la_ien_storage[45]);
	la_iena[46] = (~la_ien_storage[46]);
	la_iena[47] = (~la_ien_storage[47]);
	la_iena[48] = (~la_ien_storage[48]);
	la_iena[49] = (~la_ien_storage[49]);
	la_iena[50] = (~la_ien_storage[50]);
	la_iena[51] = (~la_ien_storage[51]);
	la_iena[52] = (~la_ien_storage[52]);
	la_iena[53] = (~la_ien_storage[53]);
	la_iena[54] = (~la_ien_storage[54]);
	la_iena[55] = (~la_ien_storage[55]);
	la_iena[56] = (~la_ien_storage[56]);
	la_iena[57] = (~la_ien_storage[57]);
	la_iena[58] = (~la_ien_storage[58]);
	la_iena[59] = (~la_ien_storage[59]);
	la_iena[60] = (~la_ien_storage[60]);
	la_iena[61] = (~la_ien_storage[61]);
	la_iena[62] = (~la_ien_storage[62]);
	la_iena[63] = (~la_ien_storage[63]);
	la_iena[64] = (~la_ien_storage[64]);
	la_iena[65] = (~la_ien_storage[65]);
	la_iena[66] = (~la_ien_storage[66]);
	la_iena[67] = (~la_ien_storage[67]);
	la_iena[68] = (~la_ien_storage[68]);
	la_iena[69] = (~la_ien_storage[69]);
	la_iena[70] = (~la_ien_storage[70]);
	la_iena[71] = (~la_ien_storage[71]);
	la_iena[72] = (~la_ien_storage[72]);
	la_iena[73] = (~la_ien_storage[73]);
	la_iena[74] = (~la_ien_storage[74]);
	la_iena[75] = (~la_ien_storage[75]);
	la_iena[76] = (~la_ien_storage[76]);
	la_iena[77] = (~la_ien_storage[77]);
	la_iena[78] = (~la_ien_storage[78]);
	la_iena[79] = (~la_ien_storage[79]);
	la_iena[80] = (~la_ien_storage[80]);
	la_iena[81] = (~la_ien_storage[81]);
	la_iena[82] = (~la_ien_storage[82]);
	la_iena[83] = (~la_ien_storage[83]);
	la_iena[84] = (~la_ien_storage[84]);
	la_iena[85] = (~la_ien_storage[85]);
	la_iena[86] = (~la_ien_storage[86]);
	la_iena[87] = (~la_ien_storage[87]);
	la_iena[88] = (~la_ien_storage[88]);
	la_iena[89] = (~la_ien_storage[89]);
	la_iena[90] = (~la_ien_storage[90]);
	la_iena[91] = (~la_ien_storage[91]);
	la_iena[92] = (~la_ien_storage[92]);
	la_iena[93] = (~la_ien_storage[93]);
	la_iena[94] = (~la_ien_storage[94]);
	la_iena[95] = (~la_ien_storage[95]);
	la_iena[96] = (~la_ien_storage[96]);
	la_iena[97] = (~la_ien_storage[97]);
	la_iena[98] = (~la_ien_storage[98]);
	la_iena[99] = (~la_ien_storage[99]);
	la_iena[100] = (~la_ien_storage[100]);
	la_iena[101] = (~la_ien_storage[101]);
	la_iena[102] = (~la_ien_storage[102]);
	la_iena[103] = (~la_ien_storage[103]);
	la_iena[104] = (~la_ien_storage[104]);
	la_iena[105] = (~la_ien_storage[105]);
	la_iena[106] = (~la_ien_storage[106]);
	la_iena[107] = (~la_ien_storage[107]);
	la_iena[108] = (~la_ien_storage[108]);
	la_iena[109] = (~la_ien_storage[109]);
	la_iena[110] = (~la_ien_storage[110]);
	la_iena[111] = (~la_ien_storage[111]);
	la_iena[112] = (~la_ien_storage[112]);
	la_iena[113] = (~la_ien_storage[113]);
	la_iena[114] = (~la_ien_storage[114]);
	la_iena[115] = (~la_ien_storage[115]);
	la_iena[116] = (~la_ien_storage[116]);
	la_iena[117] = (~la_ien_storage[117]);
	la_iena[118] = (~la_ien_storage[118]);
	la_iena[119] = (~la_ien_storage[119]);
	la_iena[120] = (~la_ien_storage[120]);
	la_iena[121] = (~la_ien_storage[121]);
	la_iena[122] = (~la_ien_storage[122]);
	la_iena[123] = (~la_ien_storage[123]);
	la_iena[124] = (~la_ien_storage[124]);
	la_iena[125] = (~la_ien_storage[125]);
	la_iena[126] = (~la_ien_storage[126]);
	la_iena[127] = (~la_ien_storage[127]);
end
always @(*) begin
	la_oenb = 128'd0;
	la_oenb[0] = (~la_oe_storage[0]);
	la_oenb[1] = (~la_oe_storage[1]);
	la_oenb[2] = (~la_oe_storage[2]);
	la_oenb[3] = (~la_oe_storage[3]);
	la_oenb[4] = (~la_oe_storage[4]);
	la_oenb[5] = (~la_oe_storage[5]);
	la_oenb[6] = (~la_oe_storage[6]);
	la_oenb[7] = (~la_oe_storage[7]);
	la_oenb[8] = (~la_oe_storage[8]);
	la_oenb[9] = (~la_oe_storage[9]);
	la_oenb[10] = (~la_oe_storage[10]);
	la_oenb[11] = (~la_oe_storage[11]);
	la_oenb[12] = (~la_oe_storage[12]);
	la_oenb[13] = (~la_oe_storage[13]);
	la_oenb[14] = (~la_oe_storage[14]);
	la_oenb[15] = (~la_oe_storage[15]);
	la_oenb[16] = (~la_oe_storage[16]);
	la_oenb[17] = (~la_oe_storage[17]);
	la_oenb[18] = (~la_oe_storage[18]);
	la_oenb[19] = (~la_oe_storage[19]);
	la_oenb[20] = (~la_oe_storage[20]);
	la_oenb[21] = (~la_oe_storage[21]);
	la_oenb[22] = (~la_oe_storage[22]);
	la_oenb[23] = (~la_oe_storage[23]);
	la_oenb[24] = (~la_oe_storage[24]);
	la_oenb[25] = (~la_oe_storage[25]);
	la_oenb[26] = (~la_oe_storage[26]);
	la_oenb[27] = (~la_oe_storage[27]);
	la_oenb[28] = (~la_oe_storage[28]);
	la_oenb[29] = (~la_oe_storage[29]);
	la_oenb[30] = (~la_oe_storage[30]);
	la_oenb[31] = (~la_oe_storage[31]);
	la_oenb[32] = (~la_oe_storage[32]);
	la_oenb[33] = (~la_oe_storage[33]);
	la_oenb[34] = (~la_oe_storage[34]);
	la_oenb[35] = (~la_oe_storage[35]);
	la_oenb[36] = (~la_oe_storage[36]);
	la_oenb[37] = (~la_oe_storage[37]);
	la_oenb[38] = (~la_oe_storage[38]);
	la_oenb[39] = (~la_oe_storage[39]);
	la_oenb[40] = (~la_oe_storage[40]);
	la_oenb[41] = (~la_oe_storage[41]);
	la_oenb[42] = (~la_oe_storage[42]);
	la_oenb[43] = (~la_oe_storage[43]);
	la_oenb[44] = (~la_oe_storage[44]);
	la_oenb[45] = (~la_oe_storage[45]);
	la_oenb[46] = (~la_oe_storage[46]);
	la_oenb[47] = (~la_oe_storage[47]);
	la_oenb[48] = (~la_oe_storage[48]);
	la_oenb[49] = (~la_oe_storage[49]);
	la_oenb[50] = (~la_oe_storage[50]);
	la_oenb[51] = (~la_oe_storage[51]);
	la_oenb[52] = (~la_oe_storage[52]);
	la_oenb[53] = (~la_oe_storage[53]);
	la_oenb[54] = (~la_oe_storage[54]);
	la_oenb[55] = (~la_oe_storage[55]);
	la_oenb[56] = (~la_oe_storage[56]);
	la_oenb[57] = (~la_oe_storage[57]);
	la_oenb[58] = (~la_oe_storage[58]);
	la_oenb[59] = (~la_oe_storage[59]);
	la_oenb[60] = (~la_oe_storage[60]);
	la_oenb[61] = (~la_oe_storage[61]);
	la_oenb[62] = (~la_oe_storage[62]);
	la_oenb[63] = (~la_oe_storage[63]);
	la_oenb[64] = (~la_oe_storage[64]);
	la_oenb[65] = (~la_oe_storage[65]);
	la_oenb[66] = (~la_oe_storage[66]);
	la_oenb[67] = (~la_oe_storage[67]);
	la_oenb[68] = (~la_oe_storage[68]);
	la_oenb[69] = (~la_oe_storage[69]);
	la_oenb[70] = (~la_oe_storage[70]);
	la_oenb[71] = (~la_oe_storage[71]);
	la_oenb[72] = (~la_oe_storage[72]);
	la_oenb[73] = (~la_oe_storage[73]);
	la_oenb[74] = (~la_oe_storage[74]);
	la_oenb[75] = (~la_oe_storage[75]);
	la_oenb[76] = (~la_oe_storage[76]);
	la_oenb[77] = (~la_oe_storage[77]);
	la_oenb[78] = (~la_oe_storage[78]);
	la_oenb[79] = (~la_oe_storage[79]);
	la_oenb[80] = (~la_oe_storage[80]);
	la_oenb[81] = (~la_oe_storage[81]);
	la_oenb[82] = (~la_oe_storage[82]);
	la_oenb[83] = (~la_oe_storage[83]);
	la_oenb[84] = (~la_oe_storage[84]);
	la_oenb[85] = (~la_oe_storage[85]);
	la_oenb[86] = (~la_oe_storage[86]);
	la_oenb[87] = (~la_oe_storage[87]);
	la_oenb[88] = (~la_oe_storage[88]);
	la_oenb[89] = (~la_oe_storage[89]);
	la_oenb[90] = (~la_oe_storage[90]);
	la_oenb[91] = (~la_oe_storage[91]);
	la_oenb[92] = (~la_oe_storage[92]);
	la_oenb[93] = (~la_oe_storage[93]);
	la_oenb[94] = (~la_oe_storage[94]);
	la_oenb[95] = (~la_oe_storage[95]);
	la_oenb[96] = (~la_oe_storage[96]);
	la_oenb[97] = (~la_oe_storage[97]);
	la_oenb[98] = (~la_oe_storage[98]);
	la_oenb[99] = (~la_oe_storage[99]);
	la_oenb[100] = (~la_oe_storage[100]);
	la_oenb[101] = (~la_oe_storage[101]);
	la_oenb[102] = (~la_oe_storage[102]);
	la_oenb[103] = (~la_oe_storage[103]);
	la_oenb[104] = (~la_oe_storage[104]);
	la_oenb[105] = (~la_oe_storage[105]);
	la_oenb[106] = (~la_oe_storage[106]);
	la_oenb[107] = (~la_oe_storage[107]);
	la_oenb[108] = (~la_oe_storage[108]);
	la_oenb[109] = (~la_oe_storage[109]);
	la_oenb[110] = (~la_oe_storage[110]);
	la_oenb[111] = (~la_oe_storage[111]);
	la_oenb[112] = (~la_oe_storage[112]);
	la_oenb[113] = (~la_oe_storage[113]);
	la_oenb[114] = (~la_oe_storage[114]);
	la_oenb[115] = (~la_oe_storage[115]);
	la_oenb[116] = (~la_oe_storage[116]);
	la_oenb[117] = (~la_oe_storage[117]);
	la_oenb[118] = (~la_oe_storage[118]);
	la_oenb[119] = (~la_oe_storage[119]);
	la_oenb[120] = (~la_oe_storage[120]);
	la_oenb[121] = (~la_oe_storage[121]);
	la_oenb[122] = (~la_oe_storage[122]);
	la_oenb[123] = (~la_oe_storage[123]);
	la_oenb[124] = (~la_oe_storage[124]);
	la_oenb[125] = (~la_oe_storage[125]);
	la_oenb[126] = (~la_oe_storage[126]);
	la_oenb[127] = (~la_oe_storage[127]);
end
always @(*) begin
	la_output = 128'd0;
    // $display($time, "=> 1st la_output=%x", la_output); //tony_debug
	la_output[0] = la_out_storage[0];
	la_output[1] = la_out_storage[1];
	la_output[2] = la_out_storage[2];
	la_output[3] = la_out_storage[3];
	la_output[4] = la_out_storage[4];
	la_output[5] = la_out_storage[5];
	la_output[6] = la_out_storage[6];
	la_output[7] = la_out_storage[7];
	la_output[8] = la_out_storage[8];
	la_output[9] = la_out_storage[9];
	la_output[10] = la_out_storage[10];
	la_output[11] = la_out_storage[11];
	la_output[12] = la_out_storage[12];
	la_output[13] = la_out_storage[13];
	la_output[14] = la_out_storage[14];
	la_output[15] = la_out_storage[15];
	la_output[16] = la_out_storage[16];
	la_output[17] = la_out_storage[17];
	la_output[18] = la_out_storage[18];
	la_output[19] = la_out_storage[19];
	la_output[20] = la_out_storage[20];
	la_output[21] = la_out_storage[21];
	la_output[22] = la_out_storage[22];
	la_output[23] = la_out_storage[23];
	la_output[24] = la_out_storage[24];
	la_output[25] = la_out_storage[25];
	la_output[26] = la_out_storage[26];
	la_output[27] = la_out_storage[27];
	la_output[28] = la_out_storage[28];
	la_output[29] = la_out_storage[29];
	la_output[30] = la_out_storage[30];
	la_output[31] = la_out_storage[31];
	la_output[32] = la_out_storage[32];
	la_output[33] = la_out_storage[33];
	la_output[34] = la_out_storage[34];
	la_output[35] = la_out_storage[35];
	la_output[36] = la_out_storage[36];
	la_output[37] = la_out_storage[37];
	la_output[38] = la_out_storage[38];
	la_output[39] = la_out_storage[39];
	la_output[40] = la_out_storage[40];
	la_output[41] = la_out_storage[41];
	la_output[42] = la_out_storage[42];
	la_output[43] = la_out_storage[43];
	la_output[44] = la_out_storage[44];
	la_output[45] = la_out_storage[45];
	la_output[46] = la_out_storage[46];
	la_output[47] = la_out_storage[47];
	la_output[48] = la_out_storage[48];
	la_output[49] = la_out_storage[49];
	la_output[50] = la_out_storage[50];
	la_output[51] = la_out_storage[51];
	la_output[52] = la_out_storage[52];
	la_output[53] = la_out_storage[53];
	la_output[54] = la_out_storage[54];
	la_output[55] = la_out_storage[55];
	la_output[56] = la_out_storage[56];
	la_output[57] = la_out_storage[57];
	la_output[58] = la_out_storage[58];
	la_output[59] = la_out_storage[59];
	la_output[60] = la_out_storage[60];
	la_output[61] = la_out_storage[61];
	la_output[62] = la_out_storage[62];
	la_output[63] = la_out_storage[63];
	la_output[64] = la_out_storage[64];
	la_output[65] = la_out_storage[65];
	la_output[66] = la_out_storage[66];
	la_output[67] = la_out_storage[67];
	la_output[68] = la_out_storage[68];
	la_output[69] = la_out_storage[69];
	la_output[70] = la_out_storage[70];
	la_output[71] = la_out_storage[71];
	la_output[72] = la_out_storage[72];
	la_output[73] = la_out_storage[73];
	la_output[74] = la_out_storage[74];
	la_output[75] = la_out_storage[75];
	la_output[76] = la_out_storage[76];
	la_output[77] = la_out_storage[77];
	la_output[78] = la_out_storage[78];
	la_output[79] = la_out_storage[79];
	la_output[80] = la_out_storage[80];
	la_output[81] = la_out_storage[81];
	la_output[82] = la_out_storage[82];
	la_output[83] = la_out_storage[83];
	la_output[84] = la_out_storage[84];
	la_output[85] = la_out_storage[85];
	la_output[86] = la_out_storage[86];
	la_output[87] = la_out_storage[87];
	la_output[88] = la_out_storage[88];
	la_output[89] = la_out_storage[89];
	la_output[90] = la_out_storage[90];
	la_output[91] = la_out_storage[91];
	la_output[92] = la_out_storage[92];
	la_output[93] = la_out_storage[93];
	la_output[94] = la_out_storage[94];
	la_output[95] = la_out_storage[95];
	la_output[96] = la_out_storage[96];
	la_output[97] = la_out_storage[97];
	la_output[98] = la_out_storage[98];
	la_output[99] = la_out_storage[99];
	la_output[100] = la_out_storage[100];
	la_output[101] = la_out_storage[101];
	la_output[102] = la_out_storage[102];
	la_output[103] = la_out_storage[103];
	la_output[104] = la_out_storage[104];
	la_output[105] = la_out_storage[105];
	la_output[106] = la_out_storage[106];
	la_output[107] = la_out_storage[107];
	la_output[108] = la_out_storage[108];
	la_output[109] = la_out_storage[109];
	la_output[110] = la_out_storage[110];
	la_output[111] = la_out_storage[111];
	la_output[112] = la_out_storage[112];
	la_output[113] = la_out_storage[113];
	la_output[114] = la_out_storage[114];
	la_output[115] = la_out_storage[115];
	la_output[116] = la_out_storage[116];
	la_output[117] = la_out_storage[117];
	la_output[118] = la_out_storage[118];
	la_output[119] = la_out_storage[119];
	la_output[120] = la_out_storage[120];
	la_output[121] = la_out_storage[121];
	la_output[122] = la_out_storage[122];
	la_output[123] = la_out_storage[123];
	la_output[124] = la_out_storage[124];
	la_output[125] = la_out_storage[125];
	la_output[126] = la_out_storage[126];
	la_output[127] = la_out_storage[127];
    // $display($time, "=> 2nd la_output=%x", la_output); //tony_debug
end
assign spi_enabled = spi_enabled_storage;
assign user_irq_ena = user_irq_ena_storage;
always @(*) begin
	gpioin0_gpioin0_trigger = 1'd0;
	if (gpioin0_gpioin0_mode_storage) begin
		gpioin0_gpioin0_trigger = (gpioin0_in_status ^ gpioin0_gpioin0_in_pads_n_d);
	end else begin
		gpioin0_gpioin0_trigger = (gpioin0_in_status ^ gpioin0_gpioin0_edge_storage);
	end
end
assign gpioin0_i00 = gpioin0_gpioin0_status;
assign gpioin0_i01 = gpioin0_gpioin0_pending;
always @(*) begin
	gpioin0_gpioin0_clear = 1'd0;
	if ((gpioin0_pending_re & gpioin0_pending_r)) begin
		gpioin0_gpioin0_clear = 1'd1;
	end
end
assign gpioin0_gpioin0_irq = (gpioin0_pending_status & gpioin0_enable_storage);
assign gpioin0_gpioin0_status = gpioin0_gpioin0_trigger;
always @(*) begin
	gpioin1_gpioin1_trigger = 1'd0;
	if (gpioin1_gpioin1_mode_storage) begin
		gpioin1_gpioin1_trigger = (gpioin1_in_status ^ gpioin1_gpioin1_in_pads_n_d);
	end else begin
		gpioin1_gpioin1_trigger = (gpioin1_in_status ^ gpioin1_gpioin1_edge_storage);
	end
end
assign gpioin1_i00 = gpioin1_gpioin1_status;
assign gpioin1_i01 = gpioin1_gpioin1_pending;
always @(*) begin
	gpioin1_gpioin1_clear = 1'd0;
	if ((gpioin1_pending_re & gpioin1_pending_r)) begin
		gpioin1_gpioin1_clear = 1'd1;
	end
end
assign gpioin1_gpioin1_irq = (gpioin1_pending_status & gpioin1_enable_storage);
assign gpioin1_gpioin1_status = gpioin1_gpioin1_trigger;
always @(*) begin
	gpioin2_gpioin2_trigger = 1'd0;
	if (gpioin2_gpioin2_mode_storage) begin
		gpioin2_gpioin2_trigger = (gpioin2_in_status ^ gpioin2_gpioin2_in_pads_n_d);
	end else begin
		gpioin2_gpioin2_trigger = (gpioin2_in_status ^ gpioin2_gpioin2_edge_storage);
	end
end
assign gpioin2_i00 = gpioin2_gpioin2_status;
assign gpioin2_i01 = gpioin2_gpioin2_pending;
always @(*) begin
	gpioin2_gpioin2_clear = 1'd0;
	if ((gpioin2_pending_re & gpioin2_pending_r)) begin
		gpioin2_gpioin2_clear = 1'd1;
	end
end
assign gpioin2_gpioin2_irq = (gpioin2_pending_status & gpioin2_enable_storage);
assign gpioin2_gpioin2_status = gpioin2_gpioin2_trigger;
always @(*) begin
	gpioin3_gpioin3_trigger = 1'd0;
	if (gpioin3_gpioin3_mode_storage) begin
		gpioin3_gpioin3_trigger = (gpioin3_in_status ^ gpioin3_gpioin3_in_pads_n_d);
	end else begin
		gpioin3_gpioin3_trigger = (gpioin3_in_status ^ gpioin3_gpioin3_edge_storage);
	end
end
assign gpioin3_i00 = gpioin3_gpioin3_status;
assign gpioin3_i01 = gpioin3_gpioin3_pending;
always @(*) begin
	gpioin3_gpioin3_clear = 1'd0;
	if ((gpioin3_pending_re & gpioin3_pending_r)) begin
		gpioin3_gpioin3_clear = 1'd1;
	end
end
assign gpioin3_gpioin3_irq = (gpioin3_pending_status & gpioin3_enable_storage);
assign gpioin3_gpioin3_status = gpioin3_gpioin3_trigger;
always @(*) begin
	gpioin4_gpioin4_trigger = 1'd0;
	if (gpioin4_gpioin4_mode_storage) begin
		gpioin4_gpioin4_trigger = (gpioin4_in_status ^ gpioin4_gpioin4_in_pads_n_d);
	end else begin
		gpioin4_gpioin4_trigger = (gpioin4_in_status ^ gpioin4_gpioin4_edge_storage);
	end
end
assign gpioin4_i00 = gpioin4_gpioin4_status;
assign gpioin4_i01 = gpioin4_gpioin4_pending;
always @(*) begin
	gpioin4_gpioin4_clear = 1'd0;
	if ((gpioin4_pending_re & gpioin4_pending_r)) begin
		gpioin4_gpioin4_clear = 1'd1;
	end
end
assign gpioin4_gpioin4_irq = (gpioin4_pending_status & gpioin4_enable_storage);
assign gpioin4_gpioin4_status = gpioin4_gpioin4_trigger;
always @(*) begin
	gpioin5_gpioin5_trigger = 1'd0;
	if (gpioin5_gpioin5_mode_storage) begin
		gpioin5_gpioin5_trigger = (gpioin5_in_status ^ gpioin5_gpioin5_in_pads_n_d);
	end else begin
		gpioin5_gpioin5_trigger = (gpioin5_in_status ^ gpioin5_gpioin5_edge_storage);
	end
end
assign gpioin5_i00 = gpioin5_gpioin5_status;
assign gpioin5_i01 = gpioin5_gpioin5_pending;
always @(*) begin
	gpioin5_gpioin5_clear = 1'd0;
	if ((gpioin5_pending_re & gpioin5_pending_r)) begin
		gpioin5_gpioin5_clear = 1'd1;
	end
end
assign gpioin5_gpioin5_irq = (gpioin5_pending_status & gpioin5_enable_storage);
assign gpioin5_gpioin5_status = gpioin5_gpioin5_trigger;

// Patrick Hack
/*
always @(*) begin
	next_state = 1'd0;
	next_state = state;
	case (state)
		1'd1: begin
			next_state = 1'd0;
		end
		default: begin
			if ((mgmtsoc_wishbone_cyc & mgmtsoc_wishbone_stb)) begin
				next_state = 1'd1;
			end
		end
	endcase
end
*/
always @(*) begin
        if( state )
          next_state = 1'd0;
        else
          next_state = mgmtsoc_wishbone_cyc & mgmtsoc_wishbone_stb;
end

always @(*) begin
	mgmtsoc_dat_w = 32'd0;
	case (state)
		1'd1: begin
		end
		default: begin
			mgmtsoc_dat_w = mgmtsoc_wishbone_dat_w;
		end
	endcase
end
always @(*) begin
	mgmtsoc_wishbone_dat_r = 32'd0;
	case (state)
		1'd1: begin
			mgmtsoc_wishbone_dat_r = mgmtsoc_dat_r;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_wishbone_ack = 1'd0;
	case (state)
		1'd1: begin
			mgmtsoc_wishbone_ack = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_adr = 14'd0;
	case (state)
		1'd1: begin
		end
		default: begin
			if ((mgmtsoc_wishbone_cyc & mgmtsoc_wishbone_stb)) begin
				mgmtsoc_adr = mgmtsoc_wishbone_adr;
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_we = 1'd0;
	case (state)
		1'd1: begin
		end
		default: begin
			if ((mgmtsoc_wishbone_cyc & mgmtsoc_wishbone_stb)) begin
				mgmtsoc_we = (mgmtsoc_wishbone_we & (mgmtsoc_wishbone_sel != 1'd0));
			end
		end
	endcase
end
assign shared_adr = comb_array_muxed0;
assign shared_dat_w = comb_array_muxed1;
assign shared_sel = comb_array_muxed2;
assign shared_cyc = comb_array_muxed3;
assign shared_stb = comb_array_muxed4;
assign shared_we = comb_array_muxed5;
assign shared_cti = comb_array_muxed6;
assign shared_bte = comb_array_muxed7;
assign mgmtsoc_ibus_ibus_dat_r = shared_dat_r;
assign mgmtsoc_dbus_dbus_dat_r = shared_dat_r;
assign dbg_uart_wishbone_dat_r = shared_dat_r;
assign mgmtsoc_ibus_ibus_ack = (shared_ack & (grant == 1'd0));
assign mgmtsoc_dbus_dbus_ack = (shared_ack & (grant == 1'd1));
assign dbg_uart_wishbone_ack = (shared_ack & (grant == 2'd2));
assign mgmtsoc_ibus_ibus_err = (shared_err & (grant == 1'd0));
assign mgmtsoc_dbus_dbus_err = (shared_err & (grant == 1'd1));
assign dbg_uart_wishbone_err = (shared_err & (grant == 2'd2));
assign request = {dbg_uart_wishbone_cyc, mgmtsoc_dbus_dbus_cyc, mgmtsoc_ibus_ibus_cyc};
always @(*) begin
	slave_sel = 7'd0;
	slave_sel[0] = (shared_adr[29:6] == 24'd15732480);
	slave_sel[1] = (shared_adr[29:8] == 1'd0);
	slave_sel[2] = (shared_adr[29:7] == 2'd2);
	slave_sel[3] = (shared_adr[29:22] == 5'd16);
	slave_sel[4] = (shared_adr[29:26] == 2'd3);
	slave_sel[5] = (shared_adr[29:20] == 8'd152);
	slave_sel[6] = (shared_adr[29:14] == 16'd61440);
end
assign mgmtsoc_vexriscv_debug_bus_adr = shared_adr;
assign mgmtsoc_vexriscv_debug_bus_dat_w = shared_dat_w;
assign mgmtsoc_vexriscv_debug_bus_sel = shared_sel;
assign mgmtsoc_vexriscv_debug_bus_stb = shared_stb;
assign mgmtsoc_vexriscv_debug_bus_we = shared_we;
assign mgmtsoc_vexriscv_debug_bus_cti = shared_cti;
assign mgmtsoc_vexriscv_debug_bus_bte = shared_bte;
assign dff_bus_adr = shared_adr;
assign dff_bus_dat_w = shared_dat_w;
assign dff_bus_sel = shared_sel;
assign dff_bus_stb = shared_stb;
assign dff_bus_we = shared_we;
assign dff_bus_cti = shared_cti;
assign dff_bus_bte = shared_bte;
assign dff2_bus_adr = shared_adr;
assign dff2_bus_dat_w = shared_dat_w;
assign dff2_bus_sel = shared_sel;
assign dff2_bus_stb = shared_stb;
assign dff2_bus_we = shared_we;
assign dff2_bus_cti = shared_cti;
assign dff2_bus_bte = shared_bte;
assign mgmtsoc_litespimmap_bus_adr = shared_adr;
assign mgmtsoc_litespimmap_bus_dat_w = shared_dat_w;
assign mgmtsoc_litespimmap_bus_sel = shared_sel;
assign mgmtsoc_litespimmap_bus_stb = shared_stb;
assign mgmtsoc_litespimmap_bus_we = shared_we;
assign mgmtsoc_litespimmap_bus_cti = shared_cti;
assign mgmtsoc_litespimmap_bus_bte = shared_bte;
assign mprj_adr = shared_adr;
assign mprj_dat_w = shared_dat_w;
assign mprj_sel = shared_sel;
assign mprj_stb = shared_stb;
assign mprj_we = shared_we;
assign mprj_cti = shared_cti;
assign mprj_bte = shared_bte;
assign hk_adr = shared_adr;
assign hk_dat_w = shared_dat_w;
assign hk_sel = shared_sel;
assign hk_stb = shared_stb;
assign hk_we = shared_we;
assign hk_cti = shared_cti;
assign hk_bte = shared_bte;
assign mgmtsoc_wishbone_adr = shared_adr;
assign mgmtsoc_wishbone_dat_w = shared_dat_w;
assign mgmtsoc_wishbone_sel = shared_sel;
assign mgmtsoc_wishbone_stb = shared_stb;
assign mgmtsoc_wishbone_we = shared_we;
assign mgmtsoc_wishbone_cti = shared_cti;
assign mgmtsoc_wishbone_bte = shared_bte;
assign mgmtsoc_vexriscv_debug_bus_cyc = (shared_cyc & slave_sel[0]);
assign dff_bus_cyc = (shared_cyc & slave_sel[1]);
assign dff2_bus_cyc = (shared_cyc & slave_sel[2]);
assign mgmtsoc_litespimmap_bus_cyc = (shared_cyc & slave_sel[3]);
assign mprj_cyc = (shared_cyc & slave_sel[4]);
assign hk_cyc = (shared_cyc & slave_sel[5]);
assign mgmtsoc_wishbone_cyc = (shared_cyc & slave_sel[6]);
always @(*) begin
	shared_ack = 1'd0;
	shared_ack = ((((((mgmtsoc_vexriscv_debug_bus_ack | dff_bus_ack) | dff2_bus_ack) | mgmtsoc_litespimmap_bus_ack) | mprj_ack) | hk_ack) | mgmtsoc_wishbone_ack);
	if (done) begin
		shared_ack = 1'd1;
	end
end
assign shared_err = ((((((mgmtsoc_vexriscv_debug_bus_err | dff_bus_err) | dff2_bus_err) | mgmtsoc_litespimmap_bus_err) | mprj_err) | hk_err) | mgmtsoc_wishbone_err);
always @(*) begin
	shared_dat_r = 32'd0;
	shared_dat_r = ((((((({32{slave_sel_r[0]}} & mgmtsoc_vexriscv_debug_bus_dat_r) | ({32{slave_sel_r[1]}} & dff_bus_dat_r)) | ({32{slave_sel_r[2]}} & dff2_bus_dat_r)) | ({32{slave_sel_r[3]}} & mgmtsoc_litespimmap_bus_dat_r)) | ({32{slave_sel_r[4]}} & mprj_dat_r)) | ({32{slave_sel_r[5]}} & hk_dat_r)) | ({32{slave_sel_r[6]}} & mgmtsoc_wishbone_dat_r));
	if (done) begin
		shared_dat_r = 32'd4294967295;
	end
end
assign wait_1 = ((shared_stb & shared_cyc) & (~shared_ack));
always @(*) begin
	error = 1'd0;
	if (done) begin
		error = 1'd1;
	end
end
assign done = (count == 1'd0);
assign csrbank0_sel = (interface0_bank_bus_adr[13:9] == 1'd0);
assign csrbank0_reset0_r = interface0_bank_bus_dat_w[1:0];
always @(*) begin
	csrbank0_reset0_re = 1'd0;
	if ((csrbank0_sel & (interface0_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank0_reset0_re = interface0_bank_bus_we;
	end
end
always @(*) begin
	csrbank0_reset0_we = 1'd0;
	if ((csrbank0_sel & (interface0_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank0_reset0_we = (~interface0_bank_bus_we);
	end
end
assign csrbank0_scratch0_r = interface0_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank0_scratch0_we = 1'd0;
	if ((csrbank0_sel & (interface0_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank0_scratch0_we = (~interface0_bank_bus_we);
	end
end
always @(*) begin
	csrbank0_scratch0_re = 1'd0;
	if ((csrbank0_sel & (interface0_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank0_scratch0_re = interface0_bank_bus_we;
	end
end
assign csrbank0_bus_errors_r = interface0_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank0_bus_errors_re = 1'd0;
	if ((csrbank0_sel & (interface0_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank0_bus_errors_re = interface0_bank_bus_we;
	end
end
always @(*) begin
	csrbank0_bus_errors_we = 1'd0;
	if ((csrbank0_sel & (interface0_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank0_bus_errors_we = (~interface0_bank_bus_we);
	end
end
always @(*) begin
	mgmtsoc_soc_rst = 1'd0;
	if (mgmtsoc_reset_re) begin
		mgmtsoc_soc_rst = mgmtsoc_reset_storage[0];
	end
end
assign mgmtsoc_cpu_rst = mgmtsoc_reset_storage[1];
assign csrbank0_reset0_w = mgmtsoc_reset_storage[1:0];
assign csrbank0_scratch0_w = mgmtsoc_scratch_storage[31:0];
assign csrbank0_bus_errors_w = mgmtsoc_bus_errors_status[31:0];
assign mgmtsoc_bus_errors_we = csrbank0_bus_errors_we;
assign csrbank1_sel = (interface1_bank_bus_adr[13:9] == 1'd1);
assign csrbank1_out0_r = interface1_bank_bus_dat_w[0];
always @(*) begin
	csrbank1_out0_we = 1'd0;
	if ((csrbank1_sel & (interface1_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank1_out0_we = (~interface1_bank_bus_we);
	end
end
always @(*) begin
	csrbank1_out0_re = 1'd0;
	if ((csrbank1_sel & (interface1_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank1_out0_re = interface1_bank_bus_we;
	end
end
assign csrbank1_out0_w = debug_mode_storage;
assign csrbank2_sel = (interface2_bank_bus_adr[13:9] == 2'd2);
assign csrbank2_out0_r = interface2_bank_bus_dat_w[0];
always @(*) begin
	csrbank2_out0_we = 1'd0;
	if ((csrbank2_sel & (interface2_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank2_out0_we = (~interface2_bank_bus_we);
	end
end
always @(*) begin
	csrbank2_out0_re = 1'd0;
	if ((csrbank2_sel & (interface2_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank2_out0_re = interface2_bank_bus_we;
	end
end
assign csrbank2_out0_w = debug_oeb_storage;
assign csrbank3_sel = (interface3_bank_bus_adr[13:9] == 2'd3);
assign csrbank3_mmap_dummy_bits0_r = interface3_bank_bus_dat_w[7:0];
always @(*) begin
	csrbank3_mmap_dummy_bits0_re = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank3_mmap_dummy_bits0_re = interface3_bank_bus_we;
	end
end
always @(*) begin
	csrbank3_mmap_dummy_bits0_we = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank3_mmap_dummy_bits0_we = (~interface3_bank_bus_we);
	end
end
assign csrbank3_master_cs0_r = interface3_bank_bus_dat_w[0];
always @(*) begin
	csrbank3_master_cs0_re = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank3_master_cs0_re = interface3_bank_bus_we;
	end
end
always @(*) begin
	csrbank3_master_cs0_we = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank3_master_cs0_we = (~interface3_bank_bus_we);
	end
end
assign csrbank3_master_phyconfig0_r = interface3_bank_bus_dat_w[23:0];
always @(*) begin
	csrbank3_master_phyconfig0_we = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank3_master_phyconfig0_we = (~interface3_bank_bus_we);
	end
end
always @(*) begin
	csrbank3_master_phyconfig0_re = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank3_master_phyconfig0_re = interface3_bank_bus_we;
	end
end
assign mgmtsoc_master_rxtx_r = interface3_bank_bus_dat_w[31:0];
always @(*) begin
	mgmtsoc_master_rxtx_re = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 2'd3))) begin
		mgmtsoc_master_rxtx_re = interface3_bank_bus_we;
	end
end
always @(*) begin
	mgmtsoc_master_rxtx_we = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 2'd3))) begin
		mgmtsoc_master_rxtx_we = (~interface3_bank_bus_we);
	end
end
assign csrbank3_master_status_r = interface3_bank_bus_dat_w[1:0];
always @(*) begin
	csrbank3_master_status_re = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank3_master_status_re = interface3_bank_bus_we;
	end
end
always @(*) begin
	csrbank3_master_status_we = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank3_master_status_we = (~interface3_bank_bus_we);
	end
end
assign csrbank3_mmap_dummy_bits0_w = mgmtsoc_litespimmap_storage[7:0];
assign csrbank3_master_cs0_w = mgmtsoc_master_cs_storage;
assign mgmtsoc_master_len = mgmtsoc_master_phyconfig_storage[7:0];
assign mgmtsoc_master_width = mgmtsoc_master_phyconfig_storage[11:8];
assign mgmtsoc_master_mask = mgmtsoc_master_phyconfig_storage[23:16];
assign csrbank3_master_phyconfig0_w = mgmtsoc_master_phyconfig_storage[23:0];
always @(*) begin
	mgmtsoc_master_status_status = 2'd0;
	mgmtsoc_master_status_status[0] = mgmtsoc_master_tx_ready;
	mgmtsoc_master_status_status[1] = mgmtsoc_master_rx_ready;
end
assign csrbank3_master_status_w = mgmtsoc_master_status_status[1:0];
assign mgmtsoc_master_status_we = csrbank3_master_status_we;
assign csrbank4_sel = (interface4_bank_bus_adr[13:9] == 3'd4);
assign csrbank4_clk_divisor0_r = interface4_bank_bus_dat_w[7:0];
always @(*) begin
	csrbank4_clk_divisor0_we = 1'd0;
	if ((csrbank4_sel & (interface4_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank4_clk_divisor0_we = (~interface4_bank_bus_we);
	end
end
always @(*) begin
	csrbank4_clk_divisor0_re = 1'd0;
	if ((csrbank4_sel & (interface4_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank4_clk_divisor0_re = interface4_bank_bus_we;
	end
end
assign csrbank4_clk_divisor0_w = mgmtsoc_litespisdrphycore_storage[7:0];
assign csrbank5_sel = (interface5_bank_bus_adr[13:9] == 3'd5);
assign csrbank5_mode10_r = interface5_bank_bus_dat_w[0];
always @(*) begin
	csrbank5_mode10_we = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank5_mode10_we = (~interface5_bank_bus_we);
	end
end
always @(*) begin
	csrbank5_mode10_re = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank5_mode10_re = interface5_bank_bus_we;
	end
end
assign csrbank5_mode00_r = interface5_bank_bus_dat_w[0];
always @(*) begin
	csrbank5_mode00_re = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank5_mode00_re = interface5_bank_bus_we;
	end
end
always @(*) begin
	csrbank5_mode00_we = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank5_mode00_we = (~interface5_bank_bus_we);
	end
end
assign csrbank5_ien0_r = interface5_bank_bus_dat_w[0];
always @(*) begin
	csrbank5_ien0_we = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank5_ien0_we = (~interface5_bank_bus_we);
	end
end
always @(*) begin
	csrbank5_ien0_re = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank5_ien0_re = interface5_bank_bus_we;
	end
end
assign csrbank5_oe0_r = interface5_bank_bus_dat_w[0];
always @(*) begin
	csrbank5_oe0_we = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank5_oe0_we = (~interface5_bank_bus_we);
	end
end
always @(*) begin
	csrbank5_oe0_re = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank5_oe0_re = interface5_bank_bus_we;
	end
end
assign csrbank5_in_r = interface5_bank_bus_dat_w[0];
always @(*) begin
	csrbank5_in_re = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank5_in_re = interface5_bank_bus_we;
	end
end
always @(*) begin
	csrbank5_in_we = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank5_in_we = (~interface5_bank_bus_we);
	end
end
assign csrbank5_out0_r = interface5_bank_bus_dat_w[0];
always @(*) begin
	csrbank5_out0_we = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank5_out0_we = (~interface5_bank_bus_we);
	end
end
always @(*) begin
	csrbank5_out0_re = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank5_out0_re = interface5_bank_bus_we;
	end
end
assign csrbank5_mode10_w = gpio_mode1_storage;
assign csrbank5_mode00_w = gpio_mode0_storage;
assign csrbank5_ien0_w = gpio_ien_storage;
assign csrbank5_oe0_w = gpio_oe_storage;
assign csrbank5_in_w = gpio_in_status;
assign gpio_in_we = csrbank5_in_we;
assign csrbank5_out0_w = gpio_out_storage;
assign csrbank6_sel = (interface6_bank_bus_adr[13:9] == 3'd6);
assign csrbank6_ien3_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_ien3_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank6_ien3_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_ien3_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank6_ien3_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_ien2_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_ien2_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank6_ien2_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_ien2_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank6_ien2_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_ien1_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_ien1_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank6_ien1_we = (~interface6_bank_bus_we);
	end
end
always @(*) begin
	csrbank6_ien1_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank6_ien1_re = interface6_bank_bus_we;
	end
end
assign csrbank6_ien0_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_ien0_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank6_ien0_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_ien0_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank6_ien0_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_oe3_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_oe3_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank6_oe3_we = (~interface6_bank_bus_we);
	end
end
always @(*) begin
	csrbank6_oe3_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank6_oe3_re = interface6_bank_bus_we;
	end
end
assign csrbank6_oe2_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_oe2_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank6_oe2_we = (~interface6_bank_bus_we);
	end
end
always @(*) begin
	csrbank6_oe2_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank6_oe2_re = interface6_bank_bus_we;
	end
end
assign csrbank6_oe1_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_oe1_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank6_oe1_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_oe1_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank6_oe1_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_oe0_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_oe0_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd7))) begin
		csrbank6_oe0_we = (~interface6_bank_bus_we);
	end
end
always @(*) begin
	csrbank6_oe0_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd7))) begin
		csrbank6_oe0_re = interface6_bank_bus_we;
	end
end
assign csrbank6_in3_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_in3_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd8))) begin
		csrbank6_in3_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_in3_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd8))) begin
		csrbank6_in3_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_in2_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_in2_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd9))) begin
		csrbank6_in2_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_in2_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd9))) begin
		csrbank6_in2_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_in1_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_in1_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd10))) begin
		csrbank6_in1_we = (~interface6_bank_bus_we);
	end
end
always @(*) begin
	csrbank6_in1_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd10))) begin
		csrbank6_in1_re = interface6_bank_bus_we;
	end
end
assign csrbank6_in0_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_in0_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd11))) begin
		csrbank6_in0_we = (~interface6_bank_bus_we);
	end
end
always @(*) begin
	csrbank6_in0_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd11))) begin
		csrbank6_in0_re = interface6_bank_bus_we;
	end
end
assign csrbank6_out3_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_out3_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd12))) begin
		csrbank6_out3_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_out3_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd12))) begin
		csrbank6_out3_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_out2_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_out2_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd13))) begin
		csrbank6_out2_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_out2_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd13))) begin
		csrbank6_out2_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_out1_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_out1_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd14))) begin
		csrbank6_out1_we = (~interface6_bank_bus_we);
	end
end
always @(*) begin
	csrbank6_out1_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd14))) begin
		csrbank6_out1_re = interface6_bank_bus_we;
	end
end
assign csrbank6_out0_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_out0_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd15))) begin
		csrbank6_out0_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_out0_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd15))) begin
		csrbank6_out0_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_ien3_w = la_ien_storage[127:96];
assign csrbank6_ien2_w = la_ien_storage[95:64];
assign csrbank6_ien1_w = la_ien_storage[63:32];
assign csrbank6_ien0_w = la_ien_storage[31:0];
assign csrbank6_oe3_w = la_oe_storage[127:96];
assign csrbank6_oe2_w = la_oe_storage[95:64];
assign csrbank6_oe1_w = la_oe_storage[63:32];
assign csrbank6_oe0_w = la_oe_storage[31:0];
assign csrbank6_in3_w = la_in_status[127:96];
assign csrbank6_in2_w = la_in_status[95:64];
assign csrbank6_in1_w = la_in_status[63:32];
assign csrbank6_in0_w = la_in_status[31:0];
assign la_in_we = csrbank6_in0_we;
assign csrbank6_out3_w = la_out_storage[127:96];
assign csrbank6_out2_w = la_out_storage[95:64];
assign csrbank6_out1_w = la_out_storage[63:32];
assign csrbank6_out0_w = la_out_storage[31:0];
assign csrbank7_sel = (interface7_bank_bus_adr[13:9] == 3'd7);
assign csrbank7_out0_r = interface7_bank_bus_dat_w[0];
always @(*) begin
	csrbank7_out0_re = 1'd0;
	if ((csrbank7_sel & (interface7_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank7_out0_re = interface7_bank_bus_we;
	end
end
always @(*) begin
	csrbank7_out0_we = 1'd0;
	if ((csrbank7_sel & (interface7_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank7_out0_we = (~interface7_bank_bus_we);
	end
end
assign csrbank7_out0_w = mprj_wb_iena_storage;
assign csrbank8_sel = (interface8_bank_bus_adr[13:9] == 4'd8);
assign csrbank8_out0_r = interface8_bank_bus_dat_w[0];
always @(*) begin
	csrbank8_out0_we = 1'd0;
	if ((csrbank8_sel & (interface8_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank8_out0_we = (~interface8_bank_bus_we);
	end
end
always @(*) begin
	csrbank8_out0_re = 1'd0;
	if ((csrbank8_sel & (interface8_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank8_out0_re = interface8_bank_bus_we;
	end
end
assign csrbank8_out0_w = spi_enabled_storage;
assign csrbank9_sel = (interface9_bank_bus_adr[13:9] == 4'd9);
assign csrbank9_control0_r = interface9_bank_bus_dat_w[15:0];
always @(*) begin
	csrbank9_control0_we = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank9_control0_we = (~interface9_bank_bus_we);
	end
end
always @(*) begin
	csrbank9_control0_re = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank9_control0_re = interface9_bank_bus_we;
	end
end
assign csrbank9_status_r = interface9_bank_bus_dat_w[0];
always @(*) begin
	csrbank9_status_re = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank9_status_re = interface9_bank_bus_we;
	end
end
always @(*) begin
	csrbank9_status_we = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank9_status_we = (~interface9_bank_bus_we);
	end
end
assign csrbank9_mosi0_r = interface9_bank_bus_dat_w[7:0];
always @(*) begin
	csrbank9_mosi0_re = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank9_mosi0_re = interface9_bank_bus_we;
	end
end
always @(*) begin
	csrbank9_mosi0_we = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank9_mosi0_we = (~interface9_bank_bus_we);
	end
end
assign csrbank9_miso_r = interface9_bank_bus_dat_w[7:0];
always @(*) begin
	csrbank9_miso_we = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank9_miso_we = (~interface9_bank_bus_we);
	end
end
always @(*) begin
	csrbank9_miso_re = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank9_miso_re = interface9_bank_bus_we;
	end
end
assign csrbank9_cs0_r = interface9_bank_bus_dat_w[16:0];
always @(*) begin
	csrbank9_cs0_we = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank9_cs0_we = (~interface9_bank_bus_we);
	end
end
always @(*) begin
	csrbank9_cs0_re = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank9_cs0_re = interface9_bank_bus_we;
	end
end
assign csrbank9_loopback0_r = interface9_bank_bus_dat_w[0];
always @(*) begin
	csrbank9_loopback0_re = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank9_loopback0_re = interface9_bank_bus_we;
	end
end
always @(*) begin
	csrbank9_loopback0_we = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank9_loopback0_we = (~interface9_bank_bus_we);
	end
end
assign csrbank9_clk_divider0_r = interface9_bank_bus_dat_w[15:0];
always @(*) begin
	csrbank9_clk_divider0_we = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank9_clk_divider0_we = (~interface9_bank_bus_we);
	end
end
always @(*) begin
	csrbank9_clk_divider0_re = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank9_clk_divider0_re = interface9_bank_bus_we;
	end
end
always @(*) begin
	spi_master_start1 = 1'd0;
	if (spi_master_control_re) begin
		spi_master_start1 = spi_master_control_storage[0];
	end
end
assign spi_master_length1 = spi_master_control_storage[15:8];
assign csrbank9_control0_w = spi_master_control_storage[15:0];
assign spi_master_status_status = spi_master_done1;
assign csrbank9_status_w = spi_master_status_status;
assign spi_master_status_we = csrbank9_status_we;
assign csrbank9_mosi0_w = spi_master_mosi_storage[7:0];
assign csrbank9_miso_w = spi_master_miso_status[7:0];
assign spi_master_miso_we = csrbank9_miso_we;
assign spi_master_sel = spi_master_cs_storage[0];
assign spi_master_mode0 = spi_master_cs_storage[16];
assign csrbank9_cs0_w = spi_master_cs_storage[16:0];
assign spi_master_mode1 = spi_master_loopback_storage;
assign csrbank9_loopback0_w = spi_master_loopback_storage;
assign csrbank9_clk_divider0_w = spimaster_storage[15:0];
assign csrbank10_sel = (interface10_bank_bus_adr[13:9] == 4'd10);
assign csrbank10_load0_r = interface10_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank10_load0_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank10_load0_re = interface10_bank_bus_we;
	end
end
always @(*) begin
	csrbank10_load0_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank10_load0_we = (~interface10_bank_bus_we);
	end
end
assign csrbank10_reload0_r = interface10_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank10_reload0_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank10_reload0_re = interface10_bank_bus_we;
	end
end
always @(*) begin
	csrbank10_reload0_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank10_reload0_we = (~interface10_bank_bus_we);
	end
end
assign csrbank10_en0_r = interface10_bank_bus_dat_w[0];
always @(*) begin
	csrbank10_en0_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank10_en0_we = (~interface10_bank_bus_we);
	end
end
always @(*) begin
	csrbank10_en0_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank10_en0_re = interface10_bank_bus_we;
	end
end
assign csrbank10_update_value0_r = interface10_bank_bus_dat_w[0];
always @(*) begin
	csrbank10_update_value0_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank10_update_value0_re = interface10_bank_bus_we;
	end
end
always @(*) begin
	csrbank10_update_value0_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank10_update_value0_we = (~interface10_bank_bus_we);
	end
end
assign csrbank10_value_r = interface10_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank10_value_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank10_value_we = (~interface10_bank_bus_we);
	end
end
always @(*) begin
	csrbank10_value_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank10_value_re = interface10_bank_bus_we;
	end
end
assign csrbank10_ev_status_r = interface10_bank_bus_dat_w[0];
always @(*) begin
	csrbank10_ev_status_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank10_ev_status_we = (~interface10_bank_bus_we);
	end
end
always @(*) begin
	csrbank10_ev_status_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank10_ev_status_re = interface10_bank_bus_we;
	end
end
assign csrbank10_ev_pending_r = interface10_bank_bus_dat_w[0];
always @(*) begin
	csrbank10_ev_pending_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank10_ev_pending_re = interface10_bank_bus_we;
	end
end
always @(*) begin
	csrbank10_ev_pending_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank10_ev_pending_we = (~interface10_bank_bus_we);
	end
end
assign csrbank10_ev_enable0_r = interface10_bank_bus_dat_w[0];
always @(*) begin
	csrbank10_ev_enable0_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd7))) begin
		csrbank10_ev_enable0_re = interface10_bank_bus_we;
	end
end
always @(*) begin
	csrbank10_ev_enable0_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd7))) begin
		csrbank10_ev_enable0_we = (~interface10_bank_bus_we);
	end
end
assign csrbank10_load0_w = mgmtsoc_load_storage[31:0];
assign csrbank10_reload0_w = mgmtsoc_reload_storage[31:0];
assign csrbank10_en0_w = mgmtsoc_en_storage;
assign csrbank10_update_value0_w = mgmtsoc_update_value_storage;
assign csrbank10_value_w = mgmtsoc_value_status[31:0];
assign mgmtsoc_value_we = csrbank10_value_we;
assign mgmtsoc_status_status = mgmtsoc_zero0;
assign csrbank10_ev_status_w = mgmtsoc_status_status;
assign mgmtsoc_status_we = csrbank10_ev_status_we;
assign mgmtsoc_pending_status = mgmtsoc_zero1;
assign csrbank10_ev_pending_w = mgmtsoc_pending_status;
assign mgmtsoc_pending_we = csrbank10_ev_pending_we;
assign mgmtsoc_zero2 = mgmtsoc_enable_storage;
assign csrbank10_ev_enable0_w = mgmtsoc_enable_storage;
assign csrbank11_sel = (interface11_bank_bus_adr[13:9] == 4'd11);
assign uart_rxtx_r = interface11_bank_bus_dat_w[7:0];
always @(*) begin
	uart_rxtx_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 1'd0))) begin
		uart_rxtx_we = (~interface11_bank_bus_we);
	end
end
always @(*) begin
	uart_rxtx_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 1'd0))) begin
		uart_rxtx_re = interface11_bank_bus_we;
	end
end
assign csrbank11_txfull_r = interface11_bank_bus_dat_w[0];
always @(*) begin
	csrbank11_txfull_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank11_txfull_we = (~interface11_bank_bus_we);
	end
end
always @(*) begin
	csrbank11_txfull_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank11_txfull_re = interface11_bank_bus_we;
	end
end
assign csrbank11_rxempty_r = interface11_bank_bus_dat_w[0];
always @(*) begin
	csrbank11_rxempty_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank11_rxempty_we = (~interface11_bank_bus_we);
	end
end
always @(*) begin
	csrbank11_rxempty_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank11_rxempty_re = interface11_bank_bus_we;
	end
end
assign csrbank11_ev_status_r = interface11_bank_bus_dat_w[1:0];
always @(*) begin
	csrbank11_ev_status_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank11_ev_status_re = interface11_bank_bus_we;
	end
end
always @(*) begin
	csrbank11_ev_status_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank11_ev_status_we = (~interface11_bank_bus_we);
	end
end
assign csrbank11_ev_pending_r = interface11_bank_bus_dat_w[1:0];
always @(*) begin
	csrbank11_ev_pending_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank11_ev_pending_re = interface11_bank_bus_we;
	end
end
always @(*) begin
	csrbank11_ev_pending_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank11_ev_pending_we = (~interface11_bank_bus_we);
	end
end
assign csrbank11_ev_enable0_r = interface11_bank_bus_dat_w[1:0];
always @(*) begin
	csrbank11_ev_enable0_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank11_ev_enable0_we = (~interface11_bank_bus_we);
	end
end
always @(*) begin
	csrbank11_ev_enable0_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank11_ev_enable0_re = interface11_bank_bus_we;
	end
end
assign csrbank11_txempty_r = interface11_bank_bus_dat_w[0];
always @(*) begin
	csrbank11_txempty_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank11_txempty_re = interface11_bank_bus_we;
	end
end
always @(*) begin
	csrbank11_txempty_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank11_txempty_we = (~interface11_bank_bus_we);
	end
end
assign csrbank11_rxfull_r = interface11_bank_bus_dat_w[0];
always @(*) begin
	csrbank11_rxfull_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd7))) begin
		csrbank11_rxfull_re = interface11_bank_bus_we;
	end
end
always @(*) begin
	csrbank11_rxfull_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd7))) begin
		csrbank11_rxfull_we = (~interface11_bank_bus_we);
	end
end
assign csrbank11_txfull_w = uart_txfull_status;
assign uart_txfull_we = csrbank11_txfull_we;
assign csrbank11_rxempty_w = uart_rxempty_status;
assign uart_rxempty_we = csrbank11_rxempty_we;
always @(*) begin
	uart_status_status = 2'd0;
	uart_status_status[0] = uart_tx0;
	uart_status_status[1] = uart_rx0;
end
assign csrbank11_ev_status_w = uart_status_status[1:0];
assign uart_status_we = csrbank11_ev_status_we;
always @(*) begin
	uart_pending_status = 2'd0;
	uart_pending_status[0] = uart_tx1;
	uart_pending_status[1] = uart_rx1;
end
assign csrbank11_ev_pending_w = uart_pending_status[1:0];
assign uart_pending_we = csrbank11_ev_pending_we;
assign uart_tx2 = uart_enable_storage[0];
assign uart_rx2 = uart_enable_storage[1];
assign csrbank11_ev_enable0_w = uart_enable_storage[1:0];
assign csrbank11_txempty_w = uart_txempty_status;
assign uart_txempty_we = csrbank11_txempty_we;
assign csrbank11_rxfull_w = uart_rxfull_status;
assign uart_rxfull_we = csrbank11_rxfull_we;
assign csrbank12_sel = (interface12_bank_bus_adr[13:9] == 4'd12);
assign csrbank12_out0_r = interface12_bank_bus_dat_w[0];
always @(*) begin
	csrbank12_out0_we = 1'd0;
	if ((csrbank12_sel & (interface12_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank12_out0_we = (~interface12_bank_bus_we);
	end
end
always @(*) begin
	csrbank12_out0_re = 1'd0;
	if ((csrbank12_sel & (interface12_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank12_out0_re = interface12_bank_bus_we;
	end
end
assign csrbank12_out0_w = uart_enabled_storage;
assign csrbank13_sel = (interface13_bank_bus_adr[13:9] == 4'd13);
assign csrbank13_in_r = interface13_bank_bus_dat_w[0];
always @(*) begin
	csrbank13_in_we = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank13_in_we = (~interface13_bank_bus_we);
	end
end
always @(*) begin
	csrbank13_in_re = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank13_in_re = interface13_bank_bus_we;
	end
end
assign csrbank13_mode0_r = interface13_bank_bus_dat_w[0];
always @(*) begin
	csrbank13_mode0_we = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank13_mode0_we = (~interface13_bank_bus_we);
	end
end
always @(*) begin
	csrbank13_mode0_re = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank13_mode0_re = interface13_bank_bus_we;
	end
end
assign csrbank13_edge0_r = interface13_bank_bus_dat_w[0];
always @(*) begin
	csrbank13_edge0_re = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank13_edge0_re = interface13_bank_bus_we;
	end
end
always @(*) begin
	csrbank13_edge0_we = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank13_edge0_we = (~interface13_bank_bus_we);
	end
end
assign csrbank13_ev_status_r = interface13_bank_bus_dat_w[0];
always @(*) begin
	csrbank13_ev_status_we = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank13_ev_status_we = (~interface13_bank_bus_we);
	end
end
always @(*) begin
	csrbank13_ev_status_re = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank13_ev_status_re = interface13_bank_bus_we;
	end
end
assign csrbank13_ev_pending_r = interface13_bank_bus_dat_w[0];
always @(*) begin
	csrbank13_ev_pending_we = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank13_ev_pending_we = (~interface13_bank_bus_we);
	end
end
always @(*) begin
	csrbank13_ev_pending_re = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank13_ev_pending_re = interface13_bank_bus_we;
	end
end
assign csrbank13_ev_enable0_r = interface13_bank_bus_dat_w[0];
always @(*) begin
	csrbank13_ev_enable0_re = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank13_ev_enable0_re = interface13_bank_bus_we;
	end
end
always @(*) begin
	csrbank13_ev_enable0_we = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank13_ev_enable0_we = (~interface13_bank_bus_we);
	end
end
assign csrbank13_in_w = gpioin0_in_status;
assign gpioin0_in_we = csrbank13_in_we;
assign csrbank13_mode0_w = gpioin0_gpioin0_mode_storage;
assign csrbank13_edge0_w = gpioin0_gpioin0_edge_storage;
assign gpioin0_status_status = gpioin0_i00;
assign csrbank13_ev_status_w = gpioin0_status_status;
assign gpioin0_status_we = csrbank13_ev_status_we;
assign gpioin0_pending_status = gpioin0_i01;
assign csrbank13_ev_pending_w = gpioin0_pending_status;
assign gpioin0_pending_we = csrbank13_ev_pending_we;
assign gpioin0_i02 = gpioin0_enable_storage;
assign csrbank13_ev_enable0_w = gpioin0_enable_storage;
assign csrbank14_sel = (interface14_bank_bus_adr[13:9] == 4'd14);
assign csrbank14_in_r = interface14_bank_bus_dat_w[0];
always @(*) begin
	csrbank14_in_we = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank14_in_we = (~interface14_bank_bus_we);
	end
end
always @(*) begin
	csrbank14_in_re = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank14_in_re = interface14_bank_bus_we;
	end
end
assign csrbank14_mode0_r = interface14_bank_bus_dat_w[0];
always @(*) begin
	csrbank14_mode0_re = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank14_mode0_re = interface14_bank_bus_we;
	end
end
always @(*) begin
	csrbank14_mode0_we = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank14_mode0_we = (~interface14_bank_bus_we);
	end
end
assign csrbank14_edge0_r = interface14_bank_bus_dat_w[0];
always @(*) begin
	csrbank14_edge0_re = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank14_edge0_re = interface14_bank_bus_we;
	end
end
always @(*) begin
	csrbank14_edge0_we = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank14_edge0_we = (~interface14_bank_bus_we);
	end
end
assign csrbank14_ev_status_r = interface14_bank_bus_dat_w[0];
always @(*) begin
	csrbank14_ev_status_we = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank14_ev_status_we = (~interface14_bank_bus_we);
	end
end
always @(*) begin
	csrbank14_ev_status_re = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank14_ev_status_re = interface14_bank_bus_we;
	end
end
assign csrbank14_ev_pending_r = interface14_bank_bus_dat_w[0];
always @(*) begin
	csrbank14_ev_pending_re = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank14_ev_pending_re = interface14_bank_bus_we;
	end
end
always @(*) begin
	csrbank14_ev_pending_we = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank14_ev_pending_we = (~interface14_bank_bus_we);
	end
end
assign csrbank14_ev_enable0_r = interface14_bank_bus_dat_w[0];
always @(*) begin
	csrbank14_ev_enable0_re = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank14_ev_enable0_re = interface14_bank_bus_we;
	end
end
always @(*) begin
	csrbank14_ev_enable0_we = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank14_ev_enable0_we = (~interface14_bank_bus_we);
	end
end
assign csrbank14_in_w = gpioin1_in_status;
assign gpioin1_in_we = csrbank14_in_we;
assign csrbank14_mode0_w = gpioin1_gpioin1_mode_storage;
assign csrbank14_edge0_w = gpioin1_gpioin1_edge_storage;
assign gpioin1_status_status = gpioin1_i00;
assign csrbank14_ev_status_w = gpioin1_status_status;
assign gpioin1_status_we = csrbank14_ev_status_we;
assign gpioin1_pending_status = gpioin1_i01;
assign csrbank14_ev_pending_w = gpioin1_pending_status;
assign gpioin1_pending_we = csrbank14_ev_pending_we;
assign gpioin1_i02 = gpioin1_enable_storage;
assign csrbank14_ev_enable0_w = gpioin1_enable_storage;
assign csrbank15_sel = (interface15_bank_bus_adr[13:9] == 4'd15);
assign csrbank15_in_r = interface15_bank_bus_dat_w[0];
always @(*) begin
	csrbank15_in_we = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank15_in_we = (~interface15_bank_bus_we);
	end
end
always @(*) begin
	csrbank15_in_re = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank15_in_re = interface15_bank_bus_we;
	end
end
assign csrbank15_mode0_r = interface15_bank_bus_dat_w[0];
always @(*) begin
	csrbank15_mode0_re = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank15_mode0_re = interface15_bank_bus_we;
	end
end
always @(*) begin
	csrbank15_mode0_we = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank15_mode0_we = (~interface15_bank_bus_we);
	end
end
assign csrbank15_edge0_r = interface15_bank_bus_dat_w[0];
always @(*) begin
	csrbank15_edge0_we = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank15_edge0_we = (~interface15_bank_bus_we);
	end
end
always @(*) begin
	csrbank15_edge0_re = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank15_edge0_re = interface15_bank_bus_we;
	end
end
assign csrbank15_ev_status_r = interface15_bank_bus_dat_w[0];
always @(*) begin
	csrbank15_ev_status_we = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank15_ev_status_we = (~interface15_bank_bus_we);
	end
end
always @(*) begin
	csrbank15_ev_status_re = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank15_ev_status_re = interface15_bank_bus_we;
	end
end
assign csrbank15_ev_pending_r = interface15_bank_bus_dat_w[0];
always @(*) begin
	csrbank15_ev_pending_re = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank15_ev_pending_re = interface15_bank_bus_we;
	end
end
always @(*) begin
	csrbank15_ev_pending_we = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank15_ev_pending_we = (~interface15_bank_bus_we);
	end
end
assign csrbank15_ev_enable0_r = interface15_bank_bus_dat_w[0];
always @(*) begin
	csrbank15_ev_enable0_we = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank15_ev_enable0_we = (~interface15_bank_bus_we);
	end
end
always @(*) begin
	csrbank15_ev_enable0_re = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank15_ev_enable0_re = interface15_bank_bus_we;
	end
end
assign csrbank15_in_w = gpioin2_in_status;
assign gpioin2_in_we = csrbank15_in_we;
assign csrbank15_mode0_w = gpioin2_gpioin2_mode_storage;
assign csrbank15_edge0_w = gpioin2_gpioin2_edge_storage;
assign gpioin2_status_status = gpioin2_i00;
assign csrbank15_ev_status_w = gpioin2_status_status;
assign gpioin2_status_we = csrbank15_ev_status_we;
assign gpioin2_pending_status = gpioin2_i01;
assign csrbank15_ev_pending_w = gpioin2_pending_status;
assign gpioin2_pending_we = csrbank15_ev_pending_we;
assign gpioin2_i02 = gpioin2_enable_storage;
assign csrbank15_ev_enable0_w = gpioin2_enable_storage;
assign csrbank16_sel = (interface16_bank_bus_adr[13:9] == 5'd16);
assign csrbank16_in_r = interface16_bank_bus_dat_w[0];
always @(*) begin
	csrbank16_in_re = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank16_in_re = interface16_bank_bus_we;
	end
end
always @(*) begin
	csrbank16_in_we = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank16_in_we = (~interface16_bank_bus_we);
	end
end
assign csrbank16_mode0_r = interface16_bank_bus_dat_w[0];
always @(*) begin
	csrbank16_mode0_re = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank16_mode0_re = interface16_bank_bus_we;
	end
end
always @(*) begin
	csrbank16_mode0_we = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank16_mode0_we = (~interface16_bank_bus_we);
	end
end
assign csrbank16_edge0_r = interface16_bank_bus_dat_w[0];
always @(*) begin
	csrbank16_edge0_we = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank16_edge0_we = (~interface16_bank_bus_we);
	end
end
always @(*) begin
	csrbank16_edge0_re = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank16_edge0_re = interface16_bank_bus_we;
	end
end
assign csrbank16_ev_status_r = interface16_bank_bus_dat_w[0];
always @(*) begin
	csrbank16_ev_status_re = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank16_ev_status_re = interface16_bank_bus_we;
	end
end
always @(*) begin
	csrbank16_ev_status_we = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank16_ev_status_we = (~interface16_bank_bus_we);
	end
end
assign csrbank16_ev_pending_r = interface16_bank_bus_dat_w[0];
always @(*) begin
	csrbank16_ev_pending_re = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank16_ev_pending_re = interface16_bank_bus_we;
	end
end
always @(*) begin
	csrbank16_ev_pending_we = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank16_ev_pending_we = (~interface16_bank_bus_we);
	end
end
assign csrbank16_ev_enable0_r = interface16_bank_bus_dat_w[0];
always @(*) begin
	csrbank16_ev_enable0_we = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank16_ev_enable0_we = (~interface16_bank_bus_we);
	end
end
always @(*) begin
	csrbank16_ev_enable0_re = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank16_ev_enable0_re = interface16_bank_bus_we;
	end
end
assign csrbank16_in_w = gpioin3_in_status;
assign gpioin3_in_we = csrbank16_in_we;
assign csrbank16_mode0_w = gpioin3_gpioin3_mode_storage;
assign csrbank16_edge0_w = gpioin3_gpioin3_edge_storage;
assign gpioin3_status_status = gpioin3_i00;
assign csrbank16_ev_status_w = gpioin3_status_status;
assign gpioin3_status_we = csrbank16_ev_status_we;
assign gpioin3_pending_status = gpioin3_i01;
assign csrbank16_ev_pending_w = gpioin3_pending_status;
assign gpioin3_pending_we = csrbank16_ev_pending_we;
assign gpioin3_i02 = gpioin3_enable_storage;
assign csrbank16_ev_enable0_w = gpioin3_enable_storage;
assign csrbank17_sel = (interface17_bank_bus_adr[13:9] == 5'd17);
assign csrbank17_in_r = interface17_bank_bus_dat_w[0];
always @(*) begin
	csrbank17_in_re = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank17_in_re = interface17_bank_bus_we;
	end
end
always @(*) begin
	csrbank17_in_we = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank17_in_we = (~interface17_bank_bus_we);
	end
end
assign csrbank17_mode0_r = interface17_bank_bus_dat_w[0];
always @(*) begin
	csrbank17_mode0_re = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank17_mode0_re = interface17_bank_bus_we;
	end
end
always @(*) begin
	csrbank17_mode0_we = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank17_mode0_we = (~interface17_bank_bus_we);
	end
end
assign csrbank17_edge0_r = interface17_bank_bus_dat_w[0];
always @(*) begin
	csrbank17_edge0_we = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank17_edge0_we = (~interface17_bank_bus_we);
	end
end
always @(*) begin
	csrbank17_edge0_re = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank17_edge0_re = interface17_bank_bus_we;
	end
end
assign csrbank17_ev_status_r = interface17_bank_bus_dat_w[0];
always @(*) begin
	csrbank17_ev_status_re = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank17_ev_status_re = interface17_bank_bus_we;
	end
end
always @(*) begin
	csrbank17_ev_status_we = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank17_ev_status_we = (~interface17_bank_bus_we);
	end
end
assign csrbank17_ev_pending_r = interface17_bank_bus_dat_w[0];
always @(*) begin
	csrbank17_ev_pending_re = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank17_ev_pending_re = interface17_bank_bus_we;
	end
end
always @(*) begin
	csrbank17_ev_pending_we = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank17_ev_pending_we = (~interface17_bank_bus_we);
	end
end
assign csrbank17_ev_enable0_r = interface17_bank_bus_dat_w[0];
always @(*) begin
	csrbank17_ev_enable0_we = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank17_ev_enable0_we = (~interface17_bank_bus_we);
	end
end
always @(*) begin
	csrbank17_ev_enable0_re = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank17_ev_enable0_re = interface17_bank_bus_we;
	end
end
assign csrbank17_in_w = gpioin4_in_status;
assign gpioin4_in_we = csrbank17_in_we;
assign csrbank17_mode0_w = gpioin4_gpioin4_mode_storage;
assign csrbank17_edge0_w = gpioin4_gpioin4_edge_storage;
assign gpioin4_status_status = gpioin4_i00;
assign csrbank17_ev_status_w = gpioin4_status_status;
assign gpioin4_status_we = csrbank17_ev_status_we;
assign gpioin4_pending_status = gpioin4_i01;
assign csrbank17_ev_pending_w = gpioin4_pending_status;
assign gpioin4_pending_we = csrbank17_ev_pending_we;
assign gpioin4_i02 = gpioin4_enable_storage;
assign csrbank17_ev_enable0_w = gpioin4_enable_storage;
assign csrbank18_sel = (interface18_bank_bus_adr[13:9] == 5'd18);
assign csrbank18_in_r = interface18_bank_bus_dat_w[0];
always @(*) begin
	csrbank18_in_re = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank18_in_re = interface18_bank_bus_we;
	end
end
always @(*) begin
	csrbank18_in_we = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank18_in_we = (~interface18_bank_bus_we);
	end
end
assign csrbank18_mode0_r = interface18_bank_bus_dat_w[0];
always @(*) begin
	csrbank18_mode0_we = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank18_mode0_we = (~interface18_bank_bus_we);
	end
end
always @(*) begin
	csrbank18_mode0_re = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank18_mode0_re = interface18_bank_bus_we;
	end
end
assign csrbank18_edge0_r = interface18_bank_bus_dat_w[0];
always @(*) begin
	csrbank18_edge0_we = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank18_edge0_we = (~interface18_bank_bus_we);
	end
end
always @(*) begin
	csrbank18_edge0_re = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank18_edge0_re = interface18_bank_bus_we;
	end
end
assign csrbank18_ev_status_r = interface18_bank_bus_dat_w[0];
always @(*) begin
	csrbank18_ev_status_re = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank18_ev_status_re = interface18_bank_bus_we;
	end
end
always @(*) begin
	csrbank18_ev_status_we = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank18_ev_status_we = (~interface18_bank_bus_we);
	end
end
assign csrbank18_ev_pending_r = interface18_bank_bus_dat_w[0];
always @(*) begin
	csrbank18_ev_pending_we = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank18_ev_pending_we = (~interface18_bank_bus_we);
	end
end
always @(*) begin
	csrbank18_ev_pending_re = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank18_ev_pending_re = interface18_bank_bus_we;
	end
end
assign csrbank18_ev_enable0_r = interface18_bank_bus_dat_w[0];
always @(*) begin
	csrbank18_ev_enable0_we = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank18_ev_enable0_we = (~interface18_bank_bus_we);
	end
end
always @(*) begin
	csrbank18_ev_enable0_re = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank18_ev_enable0_re = interface18_bank_bus_we;
	end
end
assign csrbank18_in_w = gpioin5_in_status;
assign gpioin5_in_we = csrbank18_in_we;
assign csrbank18_mode0_w = gpioin5_gpioin5_mode_storage;
assign csrbank18_edge0_w = gpioin5_gpioin5_edge_storage;
assign gpioin5_status_status = gpioin5_i00;
assign csrbank18_ev_status_w = gpioin5_status_status;
assign gpioin5_status_we = csrbank18_ev_status_we;
assign gpioin5_pending_status = gpioin5_i01;
assign csrbank18_ev_pending_w = gpioin5_pending_status;
assign gpioin5_pending_we = csrbank18_ev_pending_we;
assign gpioin5_i02 = gpioin5_enable_storage;
assign csrbank18_ev_enable0_w = gpioin5_enable_storage;
assign csrbank19_sel = (interface19_bank_bus_adr[13:9] == 5'd19);
assign csrbank19_out0_r = interface19_bank_bus_dat_w[2:0];
always @(*) begin
	csrbank19_out0_re = 1'd0;
	if ((csrbank19_sel & (interface19_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank19_out0_re = interface19_bank_bus_we;
	end
end
always @(*) begin
	csrbank19_out0_we = 1'd0;
	if ((csrbank19_sel & (interface19_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank19_out0_we = (~interface19_bank_bus_we);
	end
end
assign csrbank19_out0_w = user_irq_ena_storage[2:0];
assign csr_interconnect_adr = mgmtsoc_adr;
assign csr_interconnect_we = mgmtsoc_we;
assign csr_interconnect_dat_w = mgmtsoc_dat_w;
assign mgmtsoc_dat_r = csr_interconnect_dat_r;
assign interface0_bank_bus_adr = csr_interconnect_adr;
assign interface1_bank_bus_adr = csr_interconnect_adr;
assign interface2_bank_bus_adr = csr_interconnect_adr;
assign interface3_bank_bus_adr = csr_interconnect_adr;
assign interface4_bank_bus_adr = csr_interconnect_adr;
assign interface5_bank_bus_adr = csr_interconnect_adr;
assign interface6_bank_bus_adr = csr_interconnect_adr;
assign interface7_bank_bus_adr = csr_interconnect_adr;
assign interface8_bank_bus_adr = csr_interconnect_adr;
assign interface9_bank_bus_adr = csr_interconnect_adr;
assign interface10_bank_bus_adr = csr_interconnect_adr;
assign interface11_bank_bus_adr = csr_interconnect_adr;
assign interface12_bank_bus_adr = csr_interconnect_adr;
assign interface13_bank_bus_adr = csr_interconnect_adr;
assign interface14_bank_bus_adr = csr_interconnect_adr;
assign interface15_bank_bus_adr = csr_interconnect_adr;
assign interface16_bank_bus_adr = csr_interconnect_adr;
assign interface17_bank_bus_adr = csr_interconnect_adr;
assign interface18_bank_bus_adr = csr_interconnect_adr;
assign interface19_bank_bus_adr = csr_interconnect_adr;
assign interface0_bank_bus_we = csr_interconnect_we;
assign interface1_bank_bus_we = csr_interconnect_we;
assign interface2_bank_bus_we = csr_interconnect_we;
assign interface3_bank_bus_we = csr_interconnect_we;
assign interface4_bank_bus_we = csr_interconnect_we;
assign interface5_bank_bus_we = csr_interconnect_we;
assign interface6_bank_bus_we = csr_interconnect_we;
assign interface7_bank_bus_we = csr_interconnect_we;
assign interface8_bank_bus_we = csr_interconnect_we;
assign interface9_bank_bus_we = csr_interconnect_we;
assign interface10_bank_bus_we = csr_interconnect_we;
assign interface11_bank_bus_we = csr_interconnect_we;
assign interface12_bank_bus_we = csr_interconnect_we;
assign interface13_bank_bus_we = csr_interconnect_we;
assign interface14_bank_bus_we = csr_interconnect_we;
assign interface15_bank_bus_we = csr_interconnect_we;
assign interface16_bank_bus_we = csr_interconnect_we;
assign interface17_bank_bus_we = csr_interconnect_we;
assign interface18_bank_bus_we = csr_interconnect_we;
assign interface19_bank_bus_we = csr_interconnect_we;
assign interface0_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface1_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface2_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface3_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface4_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface5_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface6_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface7_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface8_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface9_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface10_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface11_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface12_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface13_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface14_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface15_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface16_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface17_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface18_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface19_bank_bus_dat_w = csr_interconnect_dat_w;
assign csr_interconnect_dat_r = (((((((((((((((((((interface0_bank_bus_dat_r | interface1_bank_bus_dat_r) | interface2_bank_bus_dat_r) | interface3_bank_bus_dat_r) | interface4_bank_bus_dat_r) | interface5_bank_bus_dat_r) | interface6_bank_bus_dat_r) | interface7_bank_bus_dat_r) | interface8_bank_bus_dat_r) | interface9_bank_bus_dat_r) | interface10_bank_bus_dat_r) | interface11_bank_bus_dat_r) | interface12_bank_bus_dat_r) | interface13_bank_bus_dat_r) | interface14_bank_bus_dat_r) | interface15_bank_bus_dat_r) | interface16_bank_bus_dat_r) | interface17_bank_bus_dat_r) | interface18_bank_bus_dat_r) | interface19_bank_bus_dat_r);
always @(*) begin
	comb_array_muxed0 = 30'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed0 = mgmtsoc_ibus_ibus_adr;
		end
		1'd1: begin
			comb_array_muxed0 = mgmtsoc_dbus_dbus_adr;
		end
		default: begin
			comb_array_muxed0 = dbg_uart_wishbone_adr;
		end
	endcase
end
always @(*) begin
	comb_array_muxed1 = 32'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed1 = mgmtsoc_ibus_ibus_dat_w;
		end
		1'd1: begin
			comb_array_muxed1 = mgmtsoc_dbus_dbus_dat_w;
		end
		default: begin
			comb_array_muxed1 = dbg_uart_wishbone_dat_w;
		end
	endcase
end
always @(*) begin
	comb_array_muxed2 = 4'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed2 = mgmtsoc_ibus_ibus_sel;
		end
		1'd1: begin
			comb_array_muxed2 = mgmtsoc_dbus_dbus_sel;
		end
		default: begin
			comb_array_muxed2 = dbg_uart_wishbone_sel;
		end
	endcase
end
always @(*) begin
	comb_array_muxed3 = 1'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed3 = mgmtsoc_ibus_ibus_cyc;
		end
		1'd1: begin
			comb_array_muxed3 = mgmtsoc_dbus_dbus_cyc;
		end
		default: begin
			comb_array_muxed3 = dbg_uart_wishbone_cyc;
		end
	endcase
end
always @(*) begin
	comb_array_muxed4 = 1'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed4 = mgmtsoc_ibus_ibus_stb;
		end
		1'd1: begin
			comb_array_muxed4 = mgmtsoc_dbus_dbus_stb;
		end
		default: begin
			comb_array_muxed4 = dbg_uart_wishbone_stb;
		end
	endcase
end
always @(*) begin
	comb_array_muxed5 = 1'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed5 = mgmtsoc_ibus_ibus_we;
		end
		1'd1: begin
			comb_array_muxed5 = mgmtsoc_dbus_dbus_we;
		end
		default: begin
			comb_array_muxed5 = dbg_uart_wishbone_we;
		end
	endcase
end
always @(*) begin
	comb_array_muxed6 = 3'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed6 = mgmtsoc_ibus_ibus_cti;
		end
		1'd1: begin
			comb_array_muxed6 = mgmtsoc_dbus_dbus_cti;
		end
		default: begin
			comb_array_muxed6 = dbg_uart_wishbone_cti;
		end
	endcase
end
always @(*) begin
	comb_array_muxed7 = 2'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed7 = mgmtsoc_ibus_ibus_bte;
		end
		1'd1: begin
			comb_array_muxed7 = mgmtsoc_dbus_dbus_bte;
		end
		default: begin
			comb_array_muxed7 = dbg_uart_wishbone_bte;
		end
	endcase
end
always @(*) begin
	sync_array_muxed = 1'd0;
	case (spi_master_mosi_sel)
		1'd0: begin
			sync_array_muxed = spi_master_mosi_data[0];
		end
		1'd1: begin
			sync_array_muxed = spi_master_mosi_data[1];
		end
		2'd2: begin
			sync_array_muxed = spi_master_mosi_data[2];
		end
		2'd3: begin
			sync_array_muxed = spi_master_mosi_data[3];
		end
		3'd4: begin
			sync_array_muxed = spi_master_mosi_data[4];
		end
		3'd5: begin
			sync_array_muxed = spi_master_mosi_data[5];
		end
		3'd6: begin
			sync_array_muxed = spi_master_mosi_data[6];
		end
		default: begin
			sync_array_muxed = spi_master_mosi_data[7];
		end
	endcase
end
assign sdrio_clk = sys_clk;
assign sdrio_clk_1 = sys_clk;
assign sdrio_clk_2 = sys_clk;
assign sdrio_clk_3 = sys_clk;
assign uart_phy_rx_rx = multiregimpl0_regs1;
assign dbg_uart_rx_rx = multiregimpl1_regs1;
assign gpio_in_status = multiregimpl2_regs1;
always @(*) begin
	la_in_status = 128'd0;
	la_in_status[0] = multiregimpl3_regs1;
	la_in_status[1] = multiregimpl4_regs1;
	la_in_status[2] = multiregimpl5_regs1;
	la_in_status[3] = multiregimpl6_regs1;
	la_in_status[4] = multiregimpl7_regs1;
	la_in_status[5] = multiregimpl8_regs1;
	la_in_status[6] = multiregimpl9_regs1;
	la_in_status[7] = multiregimpl10_regs1;
	la_in_status[8] = multiregimpl11_regs1;
	la_in_status[9] = multiregimpl12_regs1;
	la_in_status[10] = multiregimpl13_regs1;
	la_in_status[11] = multiregimpl14_regs1;
	la_in_status[12] = multiregimpl15_regs1;
	la_in_status[13] = multiregimpl16_regs1;
	la_in_status[14] = multiregimpl17_regs1;
	la_in_status[15] = multiregimpl18_regs1;
	la_in_status[16] = multiregimpl19_regs1;
	la_in_status[17] = multiregimpl20_regs1;
	la_in_status[18] = multiregimpl21_regs1;
	la_in_status[19] = multiregimpl22_regs1;
	la_in_status[20] = multiregimpl23_regs1;
	la_in_status[21] = multiregimpl24_regs1;
	la_in_status[22] = multiregimpl25_regs1;
	la_in_status[23] = multiregimpl26_regs1;
	la_in_status[24] = multiregimpl27_regs1;
	la_in_status[25] = multiregimpl28_regs1;
	la_in_status[26] = multiregimpl29_regs1;
	la_in_status[27] = multiregimpl30_regs1;
	la_in_status[28] = multiregimpl31_regs1;
	la_in_status[29] = multiregimpl32_regs1;
	la_in_status[30] = multiregimpl33_regs1;
	la_in_status[31] = multiregimpl34_regs1;
	la_in_status[32] = multiregimpl35_regs1;
	la_in_status[33] = multiregimpl36_regs1;
	la_in_status[34] = multiregimpl37_regs1;
	la_in_status[35] = multiregimpl38_regs1;
	la_in_status[36] = multiregimpl39_regs1;
	la_in_status[37] = multiregimpl40_regs1;
	la_in_status[38] = multiregimpl41_regs1;
	la_in_status[39] = multiregimpl42_regs1;
	la_in_status[40] = multiregimpl43_regs1;
	la_in_status[41] = multiregimpl44_regs1;
	la_in_status[42] = multiregimpl45_regs1;
	la_in_status[43] = multiregimpl46_regs1;
	la_in_status[44] = multiregimpl47_regs1;
	la_in_status[45] = multiregimpl48_regs1;
	la_in_status[46] = multiregimpl49_regs1;
	la_in_status[47] = multiregimpl50_regs1;
	la_in_status[48] = multiregimpl51_regs1;
	la_in_status[49] = multiregimpl52_regs1;
	la_in_status[50] = multiregimpl53_regs1;
	la_in_status[51] = multiregimpl54_regs1;
	la_in_status[52] = multiregimpl55_regs1;
	la_in_status[53] = multiregimpl56_regs1;
	la_in_status[54] = multiregimpl57_regs1;
	la_in_status[55] = multiregimpl58_regs1;
	la_in_status[56] = multiregimpl59_regs1;
	la_in_status[57] = multiregimpl60_regs1;
	la_in_status[58] = multiregimpl61_regs1;
	la_in_status[59] = multiregimpl62_regs1;
	la_in_status[60] = multiregimpl63_regs1;
	la_in_status[61] = multiregimpl64_regs1;
	la_in_status[62] = multiregimpl65_regs1;
	la_in_status[63] = multiregimpl66_regs1;
	la_in_status[64] = multiregimpl67_regs1;
	la_in_status[65] = multiregimpl68_regs1;
	la_in_status[66] = multiregimpl69_regs1;
	la_in_status[67] = multiregimpl70_regs1;
	la_in_status[68] = multiregimpl71_regs1;
	la_in_status[69] = multiregimpl72_regs1;
	la_in_status[70] = multiregimpl73_regs1;
	la_in_status[71] = multiregimpl74_regs1;
	la_in_status[72] = multiregimpl75_regs1;
	la_in_status[73] = multiregimpl76_regs1;
	la_in_status[74] = multiregimpl77_regs1;
	la_in_status[75] = multiregimpl78_regs1;
	la_in_status[76] = multiregimpl79_regs1;
	la_in_status[77] = multiregimpl80_regs1;
	la_in_status[78] = multiregimpl81_regs1;
	la_in_status[79] = multiregimpl82_regs1;
	la_in_status[80] = multiregimpl83_regs1;
	la_in_status[81] = multiregimpl84_regs1;
	la_in_status[82] = multiregimpl85_regs1;
	la_in_status[83] = multiregimpl86_regs1;
	la_in_status[84] = multiregimpl87_regs1;
	la_in_status[85] = multiregimpl88_regs1;
	la_in_status[86] = multiregimpl89_regs1;
	la_in_status[87] = multiregimpl90_regs1;
	la_in_status[88] = multiregimpl91_regs1;
	la_in_status[89] = multiregimpl92_regs1;
	la_in_status[90] = multiregimpl93_regs1;
	la_in_status[91] = multiregimpl94_regs1;
	la_in_status[92] = multiregimpl95_regs1;
	la_in_status[93] = multiregimpl96_regs1;
	la_in_status[94] = multiregimpl97_regs1;
	la_in_status[95] = multiregimpl98_regs1;
	la_in_status[96] = multiregimpl99_regs1;
	la_in_status[97] = multiregimpl100_regs1;
	la_in_status[98] = multiregimpl101_regs1;
	la_in_status[99] = multiregimpl102_regs1;
	la_in_status[100] = multiregimpl103_regs1;
	la_in_status[101] = multiregimpl104_regs1;
	la_in_status[102] = multiregimpl105_regs1;
	la_in_status[103] = multiregimpl106_regs1;
	la_in_status[104] = multiregimpl107_regs1;
	la_in_status[105] = multiregimpl108_regs1;
	la_in_status[106] = multiregimpl109_regs1;
	la_in_status[107] = multiregimpl110_regs1;
	la_in_status[108] = multiregimpl111_regs1;
	la_in_status[109] = multiregimpl112_regs1;
	la_in_status[110] = multiregimpl113_regs1;
	la_in_status[111] = multiregimpl114_regs1;
	la_in_status[112] = multiregimpl115_regs1;
	la_in_status[113] = multiregimpl116_regs1;
	la_in_status[114] = multiregimpl117_regs1;
	la_in_status[115] = multiregimpl118_regs1;
	la_in_status[116] = multiregimpl119_regs1;
	la_in_status[117] = multiregimpl120_regs1;
	la_in_status[118] = multiregimpl121_regs1;
	la_in_status[119] = multiregimpl122_regs1;
	la_in_status[120] = multiregimpl123_regs1;
	la_in_status[121] = multiregimpl124_regs1;
	la_in_status[122] = multiregimpl125_regs1;
	la_in_status[123] = multiregimpl126_regs1;
	la_in_status[124] = multiregimpl127_regs1;
	la_in_status[125] = multiregimpl128_regs1;
	la_in_status[126] = multiregimpl129_regs1;
	la_in_status[127] = multiregimpl130_regs1;
end
assign gpioin0_in_status = multiregimpl131_regs1;
assign gpioin1_in_status = multiregimpl132_regs1;
assign gpioin2_in_status = multiregimpl133_regs1;
assign gpioin3_in_status = multiregimpl134_regs1;
assign gpioin4_in_status = multiregimpl135_regs1;
assign gpioin5_in_status = multiregimpl136_regs1;

always @(posedge por_clk) begin
	int_rst <= core_rst;
end

always @(posedge sdrio_clk) begin
	flash_clk <= mgmtsoc_litespisdrphycore_clk;
	flash_io0_oeb <= (~mgmtsoc_litespisdrphycore_dq_oe);
	flash_io0_do <= mgmtsoc_litespisdrphycore_dq_o;
	mgmtsoc_litespisdrphycore_dq_i[1] <= flash_io1_di;
end

always @(posedge sys_clk) begin
	if ((mgmtsoc_bus_errors != 32'd4294967295)) begin
		if (mgmtsoc_bus_error) begin
			mgmtsoc_bus_errors <= (mgmtsoc_bus_errors + 1'd1);
		end
	end
	mgmtsoc_vexriscv_debug_bus_dat_r <= mgmtsoc_vexriscv_o_rsp_data;
	mgmtsoc_vexriscv_debug_reset <= (mgmtsoc_vexriscv_reset_debug_logic | sys_rst);
	if (((((mgmtsoc_vexriscv_debug_bus_stb & mgmtsoc_vexriscv_debug_bus_cyc) & (~mgmtsoc_vexriscv_transfer_in_progress)) & (~mgmtsoc_vexriscv_transfer_complete)) & (~mgmtsoc_vexriscv_transfer_wait_for_ack))) begin
		mgmtsoc_vexriscv_i_cmd_payload_data <= mgmtsoc_vexriscv_debug_bus_dat_w;
		mgmtsoc_vexriscv_i_cmd_payload_address <= ((mgmtsoc_vexriscv_debug_bus_adr[5:0] <<< 2'd2) | 1'd0);
		mgmtsoc_vexriscv_i_cmd_payload_wr <= mgmtsoc_vexriscv_debug_bus_we;
		mgmtsoc_vexriscv_i_cmd_valid <= 1'd1;
		mgmtsoc_vexriscv_transfer_in_progress <= 1'd1;
		mgmtsoc_vexriscv_transfer_complete <= 1'd0;
		mgmtsoc_vexriscv_debug_bus_ack <= 1'd0;
	end else begin
		if (mgmtsoc_vexriscv_transfer_in_progress) begin
			if (mgmtsoc_vexriscv_o_cmd_ready) begin
				mgmtsoc_vexriscv_i_cmd_valid <= 1'd0;
				mgmtsoc_vexriscv_i_cmd_payload_wr <= 1'd0;
				mgmtsoc_vexriscv_transfer_complete <= 1'd1;
				mgmtsoc_vexriscv_transfer_in_progress <= 1'd0;
			end
		end else begin
			if (mgmtsoc_vexriscv_transfer_complete) begin
				mgmtsoc_vexriscv_transfer_complete <= 1'd0;
				mgmtsoc_vexriscv_debug_bus_ack <= 1'd1;
				mgmtsoc_vexriscv_transfer_wait_for_ack <= 1'd1;
			end else begin
				if ((mgmtsoc_vexriscv_transfer_wait_for_ack & (~(mgmtsoc_vexriscv_debug_bus_stb & mgmtsoc_vexriscv_debug_bus_cyc)))) begin
					mgmtsoc_vexriscv_transfer_wait_for_ack <= 1'd0;
					mgmtsoc_vexriscv_debug_bus_ack <= 1'd0;
				end
			end
		end
	end
	if (mgmtsoc_vexriscv_o_resetOut) begin
		if ((mgmtsoc_ibus_ibus_cyc & mgmtsoc_ibus_ibus_stb)) begin
			mgmtsoc_vexriscv_ibus_err <= 1'd1;
		end else begin
			mgmtsoc_vexriscv_ibus_err <= 1'd0;
		end
		if ((mgmtsoc_dbus_dbus_cyc & mgmtsoc_dbus_dbus_stb)) begin
			mgmtsoc_vexriscv_dbus_err <= 1'd1;
		end else begin
			mgmtsoc_vexriscv_dbus_err <= 1'd0;
		end
		mgmtsoc_vexriscv_reset_debug_logic <= 1'd1;
	end else begin
		mgmtsoc_vexriscv_reset_debug_logic <= 1'd0;
	end
	if (mgmtsoc_en_storage) begin
		if ((mgmtsoc_value == 1'd0)) begin
			mgmtsoc_value <= mgmtsoc_reload_storage;
		end else begin
			mgmtsoc_value <= (mgmtsoc_value - 1'd1);
		end
	end else begin
		mgmtsoc_value <= mgmtsoc_load_storage;
	end
	if (mgmtsoc_update_value_re) begin
		mgmtsoc_value_status <= mgmtsoc_value;
	end
	if (mgmtsoc_zero_clear) begin
		mgmtsoc_zero_pending <= 1'd0;
	end
	mgmtsoc_zero_trigger_d <= mgmtsoc_zero_trigger;
	if ((mgmtsoc_zero_trigger & (~mgmtsoc_zero_trigger_d))) begin
		mgmtsoc_zero_pending <= 1'd1;
	end
	dff_bus_ack <= ((dff_bus_stb & dff_bus_cyc) & (~dff_bus_ack));
	dff2_bus_ack <= ((dff2_bus_stb & dff2_bus_cyc) & (~dff2_bus_ack));
	if (mgmtsoc_litespisdrphycore_sr_out_load) begin
		mgmtsoc_litespisdrphycore_sr_out <= (mgmtsoc_litespisdrphycore_sink_payload_data <<< (6'd32 - mgmtsoc_litespisdrphycore_sink_payload_len));
	end
	if (mgmtsoc_litespisdrphycore_sr_out_shift) begin
		case (mgmtsoc_litespisdrphycore_sink_payload_width)
			1'd1: begin
				mgmtsoc_litespisdrphycore_sr_out <= {mgmtsoc_litespisdrphycore_sr_out, mgmtsoc_litespisdrphycore0};
			end
			2'd2: begin
				mgmtsoc_litespisdrphycore_sr_out <= {mgmtsoc_litespisdrphycore_sr_out, mgmtsoc_litespisdrphycore1};
			end
			3'd4: begin
				mgmtsoc_litespisdrphycore_sr_out <= {mgmtsoc_litespisdrphycore_sr_out, mgmtsoc_litespisdrphycore2};
			end
			4'd8: begin
				mgmtsoc_litespisdrphycore_sr_out <= {mgmtsoc_litespisdrphycore_sr_out, mgmtsoc_litespisdrphycore3};
			end
		endcase
	end
	if (mgmtsoc_litespisdrphycore_sr_in_shift) begin
		case (mgmtsoc_litespisdrphycore_sink_payload_width)
			1'd1: begin
				mgmtsoc_litespisdrphycore_sr_in <= {mgmtsoc_litespisdrphycore_sr_in, mgmtsoc_litespisdrphycore_dq_i[1]};
			end
			2'd2: begin
				mgmtsoc_litespisdrphycore_sr_in <= {mgmtsoc_litespisdrphycore_sr_in, mgmtsoc_litespisdrphycore_dq_i[1:0]};
			end
			3'd4: begin
				mgmtsoc_litespisdrphycore_sr_in <= {mgmtsoc_litespisdrphycore_sr_in, mgmtsoc_litespisdrphycore_dq_i[1:0]};
			end
			4'd8: begin
				mgmtsoc_litespisdrphycore_sr_in <= {mgmtsoc_litespisdrphycore_sr_in, mgmtsoc_litespisdrphycore_dq_i[1:0]};
			end
		endcase
	end
	mgmtsoc_litespisdrphycore_posedge_reg <= mgmtsoc_litespisdrphycore_posedge;
	mgmtsoc_litespisdrphycore_posedge_reg2 <= mgmtsoc_litespisdrphycore_posedge_reg;
	if ((mgmtsoc_litespisdrphycore_en | mgmtsoc_litespisdrphycore_en_int)) begin
		if ((mgmtsoc_litespisdrphycore_cnt < mgmtsoc_litespisdrphycore_div)) begin
			mgmtsoc_litespisdrphycore_cnt <= (mgmtsoc_litespisdrphycore_cnt + 1'd1);
		end else begin
			mgmtsoc_litespisdrphycore_cnt <= 1'd0;
			mgmtsoc_litespisdrphycore_clk <= (~mgmtsoc_litespisdrphycore_clk);
		end
	end else begin
		mgmtsoc_litespisdrphycore_clk <= 1'd0;
		mgmtsoc_litespisdrphycore_cnt <= 1'd0;
	end
	if (mgmtsoc_litespisdrphycore_wait) begin
		if ((~mgmtsoc_litespisdrphycore_done)) begin
			mgmtsoc_litespisdrphycore_count <= (mgmtsoc_litespisdrphycore_count - 1'd1);
		end
	end else begin
		mgmtsoc_litespisdrphycore_count <= 4'd11;
	end
	litespiphy_state <= litespiphy_next_state;
	if (mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value_ce) begin
		mgmtsoc_litespisdrphycore_sr_cnt <= mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value;
	end
	case (litespi_grant)
		1'd0: begin
			if ((~litespi_request[0])) begin
				if (litespi_request[1]) begin
					litespi_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~litespi_request[1])) begin
				if (litespi_request[0]) begin
					litespi_grant <= 1'd0;
				end
			end
		end
	endcase
	if (mgmtsoc_litespimmap_wait) begin
		if ((~mgmtsoc_litespimmap_done)) begin
			mgmtsoc_litespimmap_count <= (mgmtsoc_litespimmap_count - 1'd1);
		end
	end else begin
		mgmtsoc_litespimmap_count <= 9'd256;
	end
	litespi_state <= litespi_next_state;
	if (mgmtsoc_litespimmap_burst_cs_litespi_next_value_ce0) begin
		mgmtsoc_litespimmap_burst_cs <= mgmtsoc_litespimmap_burst_cs_litespi_next_value0;
	end
	if (mgmtsoc_litespimmap_burst_adr_litespi_next_value_ce1) begin
		mgmtsoc_litespimmap_burst_adr <= mgmtsoc_litespimmap_burst_adr_litespi_next_value1;
	end
	if (((~mgmtsoc_master_tx_fifo_source_valid) | mgmtsoc_master_tx_fifo_source_ready)) begin
		mgmtsoc_master_tx_fifo_source_valid <= mgmtsoc_master_tx_fifo_sink_valid;
		mgmtsoc_master_tx_fifo_source_first <= mgmtsoc_master_tx_fifo_sink_first;
		mgmtsoc_master_tx_fifo_source_last <= mgmtsoc_master_tx_fifo_sink_last;
		mgmtsoc_master_tx_fifo_source_payload_data <= mgmtsoc_master_tx_fifo_sink_payload_data;
		mgmtsoc_master_tx_fifo_source_payload_len <= mgmtsoc_master_tx_fifo_sink_payload_len;
		mgmtsoc_master_tx_fifo_source_payload_width <= mgmtsoc_master_tx_fifo_sink_payload_width;
		mgmtsoc_master_tx_fifo_source_payload_mask <= mgmtsoc_master_tx_fifo_sink_payload_mask;
	end
	if (((~mgmtsoc_master_rx_fifo_source_valid) | mgmtsoc_master_rx_fifo_source_ready)) begin
		mgmtsoc_master_rx_fifo_source_valid <= mgmtsoc_master_rx_fifo_sink_valid;
		mgmtsoc_master_rx_fifo_source_first <= mgmtsoc_master_rx_fifo_sink_first;
		mgmtsoc_master_rx_fifo_source_last <= mgmtsoc_master_rx_fifo_sink_last;
		mgmtsoc_master_rx_fifo_source_payload_data <= mgmtsoc_master_rx_fifo_sink_payload_data;
	end
	spi_master_clk_divider1 <= (spi_master_clk_divider1 + 1'd1);
	if (spi_master_clk_rise) begin
		spi_clk <= spi_master_clk_enable;
	end else begin
		if (spi_master_clk_fall) begin
			spi_master_clk_divider1 <= 1'd0;
			spi_clk <= 1'd0;
		end
	end
	spi_cs_n <= (~(spi_master_cs & (spi_master_xfer_enable | (spi_master_cs_mode == 1'd1))));
	if (spi_master_mosi_latch) begin
		spi_master_mosi_data <= spi_master_mosi;
		spi_master_mosi_sel <= 3'd7;
	end else begin
		if (spi_master_clk_fall) begin
			if (spi_master_xfer_enable) begin
				spi_mosi <= sync_array_muxed;
			end
			spi_master_mosi_sel <= (spi_master_mosi_sel - 1'd1);
		end
	end
	if (spi_master_clk_rise) begin
		if (spi_master_loopback) begin
			spi_master_miso_data <= {spi_master_miso_data, spi_mosi};
		end else begin
			spi_master_miso_data <= {spi_master_miso_data, spi_miso};
		end
	end
	if (spi_master_miso_latch) begin
		spi_master_miso <= spi_master_miso_data;
	end
	spimaster_state <= spimaster_next_state;
	if (spi_master_count_spimaster_next_value_ce) begin
		spi_master_count <= spi_master_count_spimaster_next_value;
	end
	{uart_phy_tx_tick, uart_phy_tx_phase} <= 22'd4123168;
	if (uart_phy_tx_enable) begin
		{uart_phy_tx_tick, uart_phy_tx_phase} <= (uart_phy_tx_phase + 22'd4123168);
	end
	rs232phy_rs232phytx_state <= rs232phy_rs232phytx_next_state;
	if (uart_phy_tx_count_rs232phy_rs232phytx_next_value_ce0) begin
		uart_phy_tx_count <= uart_phy_tx_count_rs232phy_rs232phytx_next_value0;
	end
	if (sys_uart_tx_rs232phy_rs232phytx_next_value_ce1) begin
		sys_uart_tx <= sys_uart_tx_rs232phy_rs232phytx_next_value1;
	end
	if (uart_phy_tx_data_rs232phy_rs232phytx_next_value_ce2) begin
		uart_phy_tx_data <= uart_phy_tx_data_rs232phy_rs232phytx_next_value2;
	end
	uart_phy_rx_rx_d <= uart_phy_rx_rx;
	{uart_phy_rx_tick, uart_phy_rx_phase} <= 32'd2147483648;
	if (uart_phy_rx_enable) begin
		{uart_phy_rx_tick, uart_phy_rx_phase} <= (uart_phy_rx_phase + 22'd4123168);
	end
	rs232phy_rs232phyrx_state <= rs232phy_rs232phyrx_next_state;
	if (uart_phy_rx_count_rs232phy_rs232phyrx_next_value_ce0) begin
		uart_phy_rx_count <= uart_phy_rx_count_rs232phy_rs232phyrx_next_value0;
	end
	if (uart_phy_rx_data_rs232phy_rs232phyrx_next_value_ce1) begin
		uart_phy_rx_data <= uart_phy_rx_data_rs232phy_rs232phyrx_next_value1;
	end
	if (uart_tx_clear) begin
		uart_tx_pending <= 1'd0;
	end
	uart_tx_trigger_d <= uart_tx_trigger;
	if ((uart_tx_trigger & (~uart_tx_trigger_d))) begin
		uart_tx_pending <= 1'd1;
	end
	if (uart_rx_clear) begin
		uart_rx_pending <= 1'd0;
	end
	uart_rx_trigger_d <= uart_rx_trigger;
	if ((uart_rx_trigger & (~uart_rx_trigger_d))) begin
		uart_rx_pending <= 1'd1;
	end
	if (uart_tx_fifo_syncfifo_re) begin
		uart_tx_fifo_readable <= 1'd1;
	end else begin
		if (uart_tx_fifo_re) begin
			uart_tx_fifo_readable <= 1'd0;
		end
	end
	if (((uart_tx_fifo_syncfifo_we & uart_tx_fifo_syncfifo_writable) & (~uart_tx_fifo_replace))) begin
		uart_tx_fifo_produce <= (uart_tx_fifo_produce + 1'd1);
	end
	if (uart_tx_fifo_do_read) begin
		uart_tx_fifo_consume <= (uart_tx_fifo_consume + 1'd1);
	end
	if (((uart_tx_fifo_syncfifo_we & uart_tx_fifo_syncfifo_writable) & (~uart_tx_fifo_replace))) begin
		if ((~uart_tx_fifo_do_read)) begin
			uart_tx_fifo_level0 <= (uart_tx_fifo_level0 + 1'd1);
		end
	end else begin
		if (uart_tx_fifo_do_read) begin
			uart_tx_fifo_level0 <= (uart_tx_fifo_level0 - 1'd1);
		end
	end
	if (uart_rx_fifo_syncfifo_re) begin
		uart_rx_fifo_readable <= 1'd1;
	end else begin
		if (uart_rx_fifo_re) begin
			uart_rx_fifo_readable <= 1'd0;
		end
	end
	if (((uart_rx_fifo_syncfifo_we & uart_rx_fifo_syncfifo_writable) & (~uart_rx_fifo_replace))) begin
		uart_rx_fifo_produce <= (uart_rx_fifo_produce + 1'd1);
	end
	if (uart_rx_fifo_do_read) begin
		uart_rx_fifo_consume <= (uart_rx_fifo_consume + 1'd1);
	end
	if (((uart_rx_fifo_syncfifo_we & uart_rx_fifo_syncfifo_writable) & (~uart_rx_fifo_replace))) begin
		if ((~uart_rx_fifo_do_read)) begin
			uart_rx_fifo_level0 <= (uart_rx_fifo_level0 + 1'd1);
		end
	end else begin
		if (uart_rx_fifo_do_read) begin
			uart_rx_fifo_level0 <= (uart_rx_fifo_level0 - 1'd1);
		end
	end
	{dbg_uart_tx_tick, dbg_uart_tx_phase} <= 26'd49478023;
	if (dbg_uart_tx_enable) begin
		{dbg_uart_tx_tick, dbg_uart_tx_phase} <= (dbg_uart_tx_phase + 26'd49478023);
	end
	uartwishbonebridge_rs232phytx_state <= uartwishbonebridge_rs232phytx_next_state;
	if (dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value_ce0) begin
		dbg_uart_tx_count <= dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value0;
	end
	if (dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value_ce1) begin
		dbg_uart_dbg_uart_tx <= dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value1;
	end
	if (dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value_ce2) begin
		dbg_uart_tx_data <= dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value2;
	end
	dbg_uart_rx_rx_d <= dbg_uart_rx_rx;
	{dbg_uart_rx_tick, dbg_uart_rx_phase} <= 32'd2147483648;
	if (dbg_uart_rx_enable) begin
		{dbg_uart_rx_tick, dbg_uart_rx_phase} <= (dbg_uart_rx_phase + 26'd49478023);
	end
	uartwishbonebridge_rs232phyrx_state <= uartwishbonebridge_rs232phyrx_next_state;
	if (dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value_ce0) begin
		dbg_uart_rx_count <= dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value0;
	end
	if (dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value_ce1) begin
		dbg_uart_rx_data <= dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value1;
	end
	uartwishbonebridge_state <= uartwishbonebridge_next_state;
	if (dbg_uart_bytes_count_uartwishbonebridge_next_value_ce0) begin
		dbg_uart_bytes_count <= dbg_uart_bytes_count_uartwishbonebridge_next_value0;
	end
	if (dbg_uart_words_count_uartwishbonebridge_next_value_ce1) begin
		dbg_uart_words_count <= dbg_uart_words_count_uartwishbonebridge_next_value1;
	end
	if (dbg_uart_cmd_uartwishbonebridge_next_value_ce2) begin
		dbg_uart_cmd <= dbg_uart_cmd_uartwishbonebridge_next_value2;
	end
	if (dbg_uart_length_uartwishbonebridge_next_value_ce3) begin
		dbg_uart_length <= dbg_uart_length_uartwishbonebridge_next_value3;
	end
	if (dbg_uart_address_uartwishbonebridge_next_value_ce4) begin
		dbg_uart_address <= dbg_uart_address_uartwishbonebridge_next_value4;
	end
	if (dbg_uart_incr_uartwishbonebridge_next_value_ce5) begin
		dbg_uart_incr <= dbg_uart_incr_uartwishbonebridge_next_value5;
	end
	if (dbg_uart_data_uartwishbonebridge_next_value_ce6) begin
		dbg_uart_data <= dbg_uart_data_uartwishbonebridge_next_value6;
	end
	if (dbg_uart_reset) begin
		dbg_uart_incr <= 1'd0;
		uartwishbonebridge_state <= 3'd0;
	end
	if (dbg_uart_wait) begin
		if ((~dbg_uart_done)) begin
			dbg_uart_count <= (dbg_uart_count - 1'd1);
		end
	end else begin
		dbg_uart_count <= 20'd1000000;
	end
	gpioin0_gpioin0_in_pads_n_d <= gpioin0_in_status;
	if (gpioin0_gpioin0_clear) begin
		gpioin0_gpioin0_pending <= 1'd0;
	end
	gpioin0_gpioin0_trigger_d <= gpioin0_gpioin0_trigger;
	if ((gpioin0_gpioin0_trigger & (~gpioin0_gpioin0_trigger_d))) begin
		gpioin0_gpioin0_pending <= 1'd1;
	end
	gpioin1_gpioin1_in_pads_n_d <= gpioin1_in_status;
	if (gpioin1_gpioin1_clear) begin
		gpioin1_gpioin1_pending <= 1'd0;
	end
	gpioin1_gpioin1_trigger_d <= gpioin1_gpioin1_trigger;
	if ((gpioin1_gpioin1_trigger & (~gpioin1_gpioin1_trigger_d))) begin
		gpioin1_gpioin1_pending <= 1'd1;
	end
	gpioin2_gpioin2_in_pads_n_d <= gpioin2_in_status;
	if (gpioin2_gpioin2_clear) begin
		gpioin2_gpioin2_pending <= 1'd0;
	end
	gpioin2_gpioin2_trigger_d <= gpioin2_gpioin2_trigger;
	if ((gpioin2_gpioin2_trigger & (~gpioin2_gpioin2_trigger_d))) begin
		gpioin2_gpioin2_pending <= 1'd1;
	end
	gpioin3_gpioin3_in_pads_n_d <= gpioin3_in_status;
	if (gpioin3_gpioin3_clear) begin
		gpioin3_gpioin3_pending <= 1'd0;
	end
	gpioin3_gpioin3_trigger_d <= gpioin3_gpioin3_trigger;
	if ((gpioin3_gpioin3_trigger & (~gpioin3_gpioin3_trigger_d))) begin
		gpioin3_gpioin3_pending <= 1'd1;
	end
	gpioin4_gpioin4_in_pads_n_d <= gpioin4_in_status;
	if (gpioin4_gpioin4_clear) begin
		gpioin4_gpioin4_pending <= 1'd0;
	end
	gpioin4_gpioin4_trigger_d <= gpioin4_gpioin4_trigger;
	if ((gpioin4_gpioin4_trigger & (~gpioin4_gpioin4_trigger_d))) begin
		gpioin4_gpioin4_pending <= 1'd1;
	end
	gpioin5_gpioin5_in_pads_n_d <= gpioin5_in_status;
	if (gpioin5_gpioin5_clear) begin
		gpioin5_gpioin5_pending <= 1'd0;
	end
	gpioin5_gpioin5_trigger_d <= gpioin5_gpioin5_trigger;
	if ((gpioin5_gpioin5_trigger & (~gpioin5_gpioin5_trigger_d))) begin
		gpioin5_gpioin5_pending <= 1'd1;
	end
	state <= next_state;
	case (grant)
		1'd0: begin
			if ((~request[0])) begin
				if (request[1]) begin
					grant <= 1'd1;
				end else begin
					if (request[2]) begin
						grant <= 2'd2;
					end
				end
			end
		end
		1'd1: begin
			if ((~request[1])) begin
				if (request[2]) begin
					grant <= 2'd2;
				end else begin
					if (request[0]) begin
						grant <= 1'd0;
					end
				end
			end
		end
		2'd2: begin
			if ((~request[2])) begin
				if (request[0]) begin
					grant <= 1'd0;
				end else begin
					if (request[1]) begin
						grant <= 1'd1;
					end
				end
			end
		end
	endcase
	slave_sel_r <= slave_sel;
	if (wait_1) begin
		if ((~done)) begin
			count <= (count - 1'd1);
		end
	end else begin
		count <= 20'd1000000;
	end
	interface0_bank_bus_dat_r <= 1'd0;
	if (csrbank0_sel) begin
		case (interface0_bank_bus_adr[8:0])
			1'd0: begin
				interface0_bank_bus_dat_r <= csrbank0_reset0_w;
			end
			1'd1: begin
				interface0_bank_bus_dat_r <= csrbank0_scratch0_w;
			end
			2'd2: begin
				interface0_bank_bus_dat_r <= csrbank0_bus_errors_w;
			end
		endcase
	end
	if (csrbank0_reset0_re) begin
		mgmtsoc_reset_storage[1:0] <= csrbank0_reset0_r;
	end
	mgmtsoc_reset_re <= csrbank0_reset0_re;
	if (csrbank0_scratch0_re) begin
		mgmtsoc_scratch_storage[31:0] <= csrbank0_scratch0_r;
	end
	mgmtsoc_scratch_re <= csrbank0_scratch0_re;
	mgmtsoc_bus_errors_re <= csrbank0_bus_errors_re;
	interface1_bank_bus_dat_r <= 1'd0;
	if (csrbank1_sel) begin
		case (interface1_bank_bus_adr[8:0])
			1'd0: begin
				interface1_bank_bus_dat_r <= csrbank1_out0_w;
			end
		endcase
	end
	if (csrbank1_out0_re) begin
		debug_mode_storage <= csrbank1_out0_r;
	end
	debug_mode_re <= csrbank1_out0_re;
	interface2_bank_bus_dat_r <= 1'd0;
	if (csrbank2_sel) begin
		case (interface2_bank_bus_adr[8:0])
			1'd0: begin
				interface2_bank_bus_dat_r <= csrbank2_out0_w;
			end
		endcase
	end
	if (csrbank2_out0_re) begin
		debug_oeb_storage <= csrbank2_out0_r;
	end
	debug_oeb_re <= csrbank2_out0_re;
	interface3_bank_bus_dat_r <= 1'd0;
	if (csrbank3_sel) begin
		case (interface3_bank_bus_adr[8:0])
			1'd0: begin
				interface3_bank_bus_dat_r <= csrbank3_mmap_dummy_bits0_w;
			end
			1'd1: begin
				interface3_bank_bus_dat_r <= csrbank3_master_cs0_w;
			end
			2'd2: begin
				interface3_bank_bus_dat_r <= csrbank3_master_phyconfig0_w;
			end
			2'd3: begin
				interface3_bank_bus_dat_r <= mgmtsoc_master_rxtx_w;
			end
			3'd4: begin
				interface3_bank_bus_dat_r <= csrbank3_master_status_w;
			end
		endcase
	end
	if (csrbank3_mmap_dummy_bits0_re) begin
		mgmtsoc_litespimmap_storage[7:0] <= csrbank3_mmap_dummy_bits0_r;
	end
	mgmtsoc_litespimmap_re <= csrbank3_mmap_dummy_bits0_re;
	if (csrbank3_master_cs0_re) begin
		mgmtsoc_master_cs_storage <= csrbank3_master_cs0_r;
	end
	mgmtsoc_master_cs_re <= csrbank3_master_cs0_re;
	if (csrbank3_master_phyconfig0_re) begin
		mgmtsoc_master_phyconfig_storage[23:0] <= csrbank3_master_phyconfig0_r;
	end
	mgmtsoc_master_phyconfig_re <= csrbank3_master_phyconfig0_re;
	mgmtsoc_master_status_re <= csrbank3_master_status_re;
	interface4_bank_bus_dat_r <= 1'd0;
	if (csrbank4_sel) begin
		case (interface4_bank_bus_adr[8:0])
			1'd0: begin
				interface4_bank_bus_dat_r <= csrbank4_clk_divisor0_w;
			end
		endcase
	end
	if (csrbank4_clk_divisor0_re) begin
		mgmtsoc_litespisdrphycore_storage[7:0] <= csrbank4_clk_divisor0_r;
	end
	mgmtsoc_litespisdrphycore_re <= csrbank4_clk_divisor0_re;
	interface5_bank_bus_dat_r <= 1'd0;
	if (csrbank5_sel) begin
		case (interface5_bank_bus_adr[8:0])
			1'd0: begin
				interface5_bank_bus_dat_r <= csrbank5_mode10_w;
			end
			1'd1: begin
				interface5_bank_bus_dat_r <= csrbank5_mode00_w;
			end
			2'd2: begin
				interface5_bank_bus_dat_r <= csrbank5_ien0_w;
			end
			2'd3: begin
				interface5_bank_bus_dat_r <= csrbank5_oe0_w;
			end
			3'd4: begin
				interface5_bank_bus_dat_r <= csrbank5_in_w;
			end
			3'd5: begin
				interface5_bank_bus_dat_r <= csrbank5_out0_w;
			end
		endcase
	end
	if (csrbank5_mode10_re) begin
		gpio_mode1_storage <= csrbank5_mode10_r;
	end
	gpio_mode1_re <= csrbank5_mode10_re;
	if (csrbank5_mode00_re) begin
		gpio_mode0_storage <= csrbank5_mode00_r;
	end
	gpio_mode0_re <= csrbank5_mode00_re;
	if (csrbank5_ien0_re) begin
		gpio_ien_storage <= csrbank5_ien0_r;
	end
	gpio_ien_re <= csrbank5_ien0_re;
	if (csrbank5_oe0_re) begin
		gpio_oe_storage <= csrbank5_oe0_r;
	end
	gpio_oe_re <= csrbank5_oe0_re;
	gpio_in_re <= csrbank5_in_re;
	if (csrbank5_out0_re) begin
		gpio_out_storage <= csrbank5_out0_r;
	end
	gpio_out_re <= csrbank5_out0_re;
	interface6_bank_bus_dat_r <= 1'd0;
	if (csrbank6_sel) begin
		case (interface6_bank_bus_adr[8:0])
			1'd0: begin
				interface6_bank_bus_dat_r <= csrbank6_ien3_w;
			end
			1'd1: begin
				interface6_bank_bus_dat_r <= csrbank6_ien2_w;
			end
			2'd2: begin
				interface6_bank_bus_dat_r <= csrbank6_ien1_w;
			end
			2'd3: begin
				interface6_bank_bus_dat_r <= csrbank6_ien0_w;
			end
			3'd4: begin
				interface6_bank_bus_dat_r <= csrbank6_oe3_w;
			end
			3'd5: begin
				interface6_bank_bus_dat_r <= csrbank6_oe2_w;
			end
			3'd6: begin
				interface6_bank_bus_dat_r <= csrbank6_oe1_w;
			end
			3'd7: begin
				interface6_bank_bus_dat_r <= csrbank6_oe0_w;
			end
			4'd8: begin
				interface6_bank_bus_dat_r <= csrbank6_in3_w;
			end
			4'd9: begin
				interface6_bank_bus_dat_r <= csrbank6_in2_w;
			end
			4'd10: begin
				interface6_bank_bus_dat_r <= csrbank6_in1_w;
			end
			4'd11: begin
				interface6_bank_bus_dat_r <= csrbank6_in0_w;
			end
			4'd12: begin
				interface6_bank_bus_dat_r <= csrbank6_out3_w;
			end
			4'd13: begin
				interface6_bank_bus_dat_r <= csrbank6_out2_w;
			end
			4'd14: begin
				interface6_bank_bus_dat_r <= csrbank6_out1_w;
			end
			4'd15: begin
				interface6_bank_bus_dat_r <= csrbank6_out0_w;
			end
		endcase
	end
	if (csrbank6_ien3_re) begin
		la_ien_storage[127:96] <= csrbank6_ien3_r;
	end
	if (csrbank6_ien2_re) begin
		la_ien_storage[95:64] <= csrbank6_ien2_r;
	end
	if (csrbank6_ien1_re) begin
		la_ien_storage[63:32] <= csrbank6_ien1_r;
	end
	if (csrbank6_ien0_re) begin
		la_ien_storage[31:0] <= csrbank6_ien0_r;
	end
	la_ien_re <= csrbank6_ien0_re;
	if (csrbank6_oe3_re) begin
		la_oe_storage[127:96] <= csrbank6_oe3_r;
	end
	if (csrbank6_oe2_re) begin
		la_oe_storage[95:64] <= csrbank6_oe2_r;
	end
	if (csrbank6_oe1_re) begin
		la_oe_storage[63:32] <= csrbank6_oe1_r;
	end
	if (csrbank6_oe0_re) begin
		la_oe_storage[31:0] <= csrbank6_oe0_r;
	end
	la_oe_re <= csrbank6_oe0_re;
	la_in_re <= csrbank6_in0_re;
	if (csrbank6_out3_re) begin
		la_out_storage[127:96] <= csrbank6_out3_r;
	end
	if (csrbank6_out2_re) begin
		la_out_storage[95:64] <= csrbank6_out2_r;
	end
	if (csrbank6_out1_re) begin
		la_out_storage[63:32] <= csrbank6_out1_r;
	end
	if (csrbank6_out0_re) begin
		la_out_storage[31:0] <= csrbank6_out0_r;
	end
	la_out_re <= csrbank6_out0_re;
	interface7_bank_bus_dat_r <= 1'd0;
	if (csrbank7_sel) begin
		case (interface7_bank_bus_adr[8:0])
			1'd0: begin
				interface7_bank_bus_dat_r <= csrbank7_out0_w;
			end
		endcase
	end
	if (csrbank7_out0_re) begin
		mprj_wb_iena_storage <= csrbank7_out0_r;
	end
	mprj_wb_iena_re <= csrbank7_out0_re;
	interface8_bank_bus_dat_r <= 1'd0;
	if (csrbank8_sel) begin
		case (interface8_bank_bus_adr[8:0])
			1'd0: begin
				interface8_bank_bus_dat_r <= csrbank8_out0_w;
			end
		endcase
	end
	if (csrbank8_out0_re) begin
		spi_enabled_storage <= csrbank8_out0_r;
	end
	spi_enabled_re <= csrbank8_out0_re;
	interface9_bank_bus_dat_r <= 1'd0;
	if (csrbank9_sel) begin
		case (interface9_bank_bus_adr[8:0])
			1'd0: begin
				interface9_bank_bus_dat_r <= csrbank9_control0_w;
			end
			1'd1: begin
				interface9_bank_bus_dat_r <= csrbank9_status_w;
			end
			2'd2: begin
				interface9_bank_bus_dat_r <= csrbank9_mosi0_w;
			end
			2'd3: begin
				interface9_bank_bus_dat_r <= csrbank9_miso_w;
			end
			3'd4: begin
				interface9_bank_bus_dat_r <= csrbank9_cs0_w;
			end
			3'd5: begin
				interface9_bank_bus_dat_r <= csrbank9_loopback0_w;
			end
			3'd6: begin
				interface9_bank_bus_dat_r <= csrbank9_clk_divider0_w;
			end
		endcase
	end
	if (csrbank9_control0_re) begin
		spi_master_control_storage[15:0] <= csrbank9_control0_r;
	end
	spi_master_control_re <= csrbank9_control0_re;
	spi_master_status_re <= csrbank9_status_re;
	if (csrbank9_mosi0_re) begin
		spi_master_mosi_storage[7:0] <= csrbank9_mosi0_r;
	end
	spi_master_mosi_re <= csrbank9_mosi0_re;
	spi_master_miso_re <= csrbank9_miso_re;
	if (csrbank9_cs0_re) begin
		spi_master_cs_storage[16:0] <= csrbank9_cs0_r;
	end
	spi_master_cs_re <= csrbank9_cs0_re;
	if (csrbank9_loopback0_re) begin
		spi_master_loopback_storage <= csrbank9_loopback0_r;
	end
	spi_master_loopback_re <= csrbank9_loopback0_re;
	if (csrbank9_clk_divider0_re) begin
		spimaster_storage[15:0] <= csrbank9_clk_divider0_r;
	end
	spimaster_re <= csrbank9_clk_divider0_re;
	interface10_bank_bus_dat_r <= 1'd0;
	if (csrbank10_sel) begin
		case (interface10_bank_bus_adr[8:0])
			1'd0: begin
				interface10_bank_bus_dat_r <= csrbank10_load0_w;
			end
			1'd1: begin
				interface10_bank_bus_dat_r <= csrbank10_reload0_w;
			end
			2'd2: begin
				interface10_bank_bus_dat_r <= csrbank10_en0_w;
			end
			2'd3: begin
				interface10_bank_bus_dat_r <= csrbank10_update_value0_w;
			end
			3'd4: begin
				interface10_bank_bus_dat_r <= csrbank10_value_w;
			end
			3'd5: begin
				interface10_bank_bus_dat_r <= csrbank10_ev_status_w;
			end
			3'd6: begin
				interface10_bank_bus_dat_r <= csrbank10_ev_pending_w;
			end
			3'd7: begin
				interface10_bank_bus_dat_r <= csrbank10_ev_enable0_w;
			end
		endcase
	end
	if (csrbank10_load0_re) begin
		mgmtsoc_load_storage[31:0] <= csrbank10_load0_r;
	end
	mgmtsoc_load_re <= csrbank10_load0_re;
	if (csrbank10_reload0_re) begin
		mgmtsoc_reload_storage[31:0] <= csrbank10_reload0_r;
	end
	mgmtsoc_reload_re <= csrbank10_reload0_re;
	if (csrbank10_en0_re) begin
		mgmtsoc_en_storage <= csrbank10_en0_r;
	end
	mgmtsoc_en_re <= csrbank10_en0_re;
	if (csrbank10_update_value0_re) begin
		mgmtsoc_update_value_storage <= csrbank10_update_value0_r;
	end
	mgmtsoc_update_value_re <= csrbank10_update_value0_re;
	mgmtsoc_value_re <= csrbank10_value_re;
	mgmtsoc_status_re <= csrbank10_ev_status_re;
	if (csrbank10_ev_pending_re) begin
		mgmtsoc_pending_r <= csrbank10_ev_pending_r;
	end
	mgmtsoc_pending_re <= csrbank10_ev_pending_re;
	if (csrbank10_ev_enable0_re) begin
		mgmtsoc_enable_storage <= csrbank10_ev_enable0_r;
	end
	mgmtsoc_enable_re <= csrbank10_ev_enable0_re;
	interface11_bank_bus_dat_r <= 1'd0;
	if (csrbank11_sel) begin
		case (interface11_bank_bus_adr[8:0])
			1'd0: begin
				interface11_bank_bus_dat_r <= uart_rxtx_w;
			end
			1'd1: begin
				interface11_bank_bus_dat_r <= csrbank11_txfull_w;
			end
			2'd2: begin
				interface11_bank_bus_dat_r <= csrbank11_rxempty_w;
			end
			2'd3: begin
				interface11_bank_bus_dat_r <= csrbank11_ev_status_w;
			end
			3'd4: begin
				interface11_bank_bus_dat_r <= csrbank11_ev_pending_w;
			end
			3'd5: begin
				interface11_bank_bus_dat_r <= csrbank11_ev_enable0_w;
			end
			3'd6: begin
				interface11_bank_bus_dat_r <= csrbank11_txempty_w;
			end
			3'd7: begin
				interface11_bank_bus_dat_r <= csrbank11_rxfull_w;
			end
		endcase
	end
	uart_txfull_re <= csrbank11_txfull_re;
	uart_rxempty_re <= csrbank11_rxempty_re;
	uart_status_re <= csrbank11_ev_status_re;
	if (csrbank11_ev_pending_re) begin
		uart_pending_r[1:0] <= csrbank11_ev_pending_r;
	end
	uart_pending_re <= csrbank11_ev_pending_re;
	if (csrbank11_ev_enable0_re) begin
		uart_enable_storage[1:0] <= csrbank11_ev_enable0_r;
	end
	uart_enable_re <= csrbank11_ev_enable0_re;
	uart_txempty_re <= csrbank11_txempty_re;
	uart_rxfull_re <= csrbank11_rxfull_re;
	interface12_bank_bus_dat_r <= 1'd0;
	if (csrbank12_sel) begin
		case (interface12_bank_bus_adr[8:0])
			1'd0: begin
				interface12_bank_bus_dat_r <= csrbank12_out0_w;
			end
		endcase
	end
	if (csrbank12_out0_re) begin
		uart_enabled_storage <= csrbank12_out0_r;
	end
	uart_enabled_re <= csrbank12_out0_re;
	interface13_bank_bus_dat_r <= 1'd0;
	if (csrbank13_sel) begin
		case (interface13_bank_bus_adr[8:0])
			1'd0: begin
				interface13_bank_bus_dat_r <= csrbank13_in_w;
			end
			1'd1: begin
				interface13_bank_bus_dat_r <= csrbank13_mode0_w;
			end
			2'd2: begin
				interface13_bank_bus_dat_r <= csrbank13_edge0_w;
			end
			2'd3: begin
				interface13_bank_bus_dat_r <= csrbank13_ev_status_w;
			end
			3'd4: begin
				interface13_bank_bus_dat_r <= csrbank13_ev_pending_w;
			end
			3'd5: begin
				interface13_bank_bus_dat_r <= csrbank13_ev_enable0_w;
			end
		endcase
	end
	gpioin0_in_re <= csrbank13_in_re;
	if (csrbank13_mode0_re) begin
		gpioin0_gpioin0_mode_storage <= csrbank13_mode0_r;
	end
	gpioin0_gpioin0_mode_re <= csrbank13_mode0_re;
	if (csrbank13_edge0_re) begin
		gpioin0_gpioin0_edge_storage <= csrbank13_edge0_r;
	end
	gpioin0_gpioin0_edge_re <= csrbank13_edge0_re;
	gpioin0_status_re <= csrbank13_ev_status_re;
	if (csrbank13_ev_pending_re) begin
		gpioin0_pending_r <= csrbank13_ev_pending_r;
	end
	gpioin0_pending_re <= csrbank13_ev_pending_re;
	if (csrbank13_ev_enable0_re) begin
		gpioin0_enable_storage <= csrbank13_ev_enable0_r;
	end
	gpioin0_enable_re <= csrbank13_ev_enable0_re;
	interface14_bank_bus_dat_r <= 1'd0;
	if (csrbank14_sel) begin
		case (interface14_bank_bus_adr[8:0])
			1'd0: begin
				interface14_bank_bus_dat_r <= csrbank14_in_w;
			end
			1'd1: begin
				interface14_bank_bus_dat_r <= csrbank14_mode0_w;
			end
			2'd2: begin
				interface14_bank_bus_dat_r <= csrbank14_edge0_w;
			end
			2'd3: begin
				interface14_bank_bus_dat_r <= csrbank14_ev_status_w;
			end
			3'd4: begin
				interface14_bank_bus_dat_r <= csrbank14_ev_pending_w;
			end
			3'd5: begin
				interface14_bank_bus_dat_r <= csrbank14_ev_enable0_w;
			end
		endcase
	end
	gpioin1_in_re <= csrbank14_in_re;
	if (csrbank14_mode0_re) begin
		gpioin1_gpioin1_mode_storage <= csrbank14_mode0_r;
	end
	gpioin1_gpioin1_mode_re <= csrbank14_mode0_re;
	if (csrbank14_edge0_re) begin
		gpioin1_gpioin1_edge_storage <= csrbank14_edge0_r;
	end
	gpioin1_gpioin1_edge_re <= csrbank14_edge0_re;
	gpioin1_status_re <= csrbank14_ev_status_re;
	if (csrbank14_ev_pending_re) begin
		gpioin1_pending_r <= csrbank14_ev_pending_r;
	end
	gpioin1_pending_re <= csrbank14_ev_pending_re;
	if (csrbank14_ev_enable0_re) begin
		gpioin1_enable_storage <= csrbank14_ev_enable0_r;
	end
	gpioin1_enable_re <= csrbank14_ev_enable0_re;
	interface15_bank_bus_dat_r <= 1'd0;
	if (csrbank15_sel) begin
		case (interface15_bank_bus_adr[8:0])
			1'd0: begin
				interface15_bank_bus_dat_r <= csrbank15_in_w;
			end
			1'd1: begin
				interface15_bank_bus_dat_r <= csrbank15_mode0_w;
			end
			2'd2: begin
				interface15_bank_bus_dat_r <= csrbank15_edge0_w;
			end
			2'd3: begin
				interface15_bank_bus_dat_r <= csrbank15_ev_status_w;
			end
			3'd4: begin
				interface15_bank_bus_dat_r <= csrbank15_ev_pending_w;
			end
			3'd5: begin
				interface15_bank_bus_dat_r <= csrbank15_ev_enable0_w;
			end
		endcase
	end
	gpioin2_in_re <= csrbank15_in_re;
	if (csrbank15_mode0_re) begin
		gpioin2_gpioin2_mode_storage <= csrbank15_mode0_r;
	end
	gpioin2_gpioin2_mode_re <= csrbank15_mode0_re;
	if (csrbank15_edge0_re) begin
		gpioin2_gpioin2_edge_storage <= csrbank15_edge0_r;
	end
	gpioin2_gpioin2_edge_re <= csrbank15_edge0_re;
	gpioin2_status_re <= csrbank15_ev_status_re;
	if (csrbank15_ev_pending_re) begin
		gpioin2_pending_r <= csrbank15_ev_pending_r;
	end
	gpioin2_pending_re <= csrbank15_ev_pending_re;
	if (csrbank15_ev_enable0_re) begin
		gpioin2_enable_storage <= csrbank15_ev_enable0_r;
	end
	gpioin2_enable_re <= csrbank15_ev_enable0_re;
	interface16_bank_bus_dat_r <= 1'd0;
	if (csrbank16_sel) begin
		case (interface16_bank_bus_adr[8:0])
			1'd0: begin
				interface16_bank_bus_dat_r <= csrbank16_in_w;
			end
			1'd1: begin
				interface16_bank_bus_dat_r <= csrbank16_mode0_w;
			end
			2'd2: begin
				interface16_bank_bus_dat_r <= csrbank16_edge0_w;
			end
			2'd3: begin
				interface16_bank_bus_dat_r <= csrbank16_ev_status_w;
			end
			3'd4: begin
				interface16_bank_bus_dat_r <= csrbank16_ev_pending_w;
			end
			3'd5: begin
				interface16_bank_bus_dat_r <= csrbank16_ev_enable0_w;
			end
		endcase
	end
	gpioin3_in_re <= csrbank16_in_re;
	if (csrbank16_mode0_re) begin
		gpioin3_gpioin3_mode_storage <= csrbank16_mode0_r;
	end
	gpioin3_gpioin3_mode_re <= csrbank16_mode0_re;
	if (csrbank16_edge0_re) begin
		gpioin3_gpioin3_edge_storage <= csrbank16_edge0_r;
	end
	gpioin3_gpioin3_edge_re <= csrbank16_edge0_re;
	gpioin3_status_re <= csrbank16_ev_status_re;
	if (csrbank16_ev_pending_re) begin
		gpioin3_pending_r <= csrbank16_ev_pending_r;
	end
	gpioin3_pending_re <= csrbank16_ev_pending_re;
	if (csrbank16_ev_enable0_re) begin
		gpioin3_enable_storage <= csrbank16_ev_enable0_r;
	end
	gpioin3_enable_re <= csrbank16_ev_enable0_re;
	interface17_bank_bus_dat_r <= 1'd0;
	if (csrbank17_sel) begin
		case (interface17_bank_bus_adr[8:0])
			1'd0: begin
				interface17_bank_bus_dat_r <= csrbank17_in_w;
			end
			1'd1: begin
				interface17_bank_bus_dat_r <= csrbank17_mode0_w;
			end
			2'd2: begin
				interface17_bank_bus_dat_r <= csrbank17_edge0_w;
			end
			2'd3: begin
				interface17_bank_bus_dat_r <= csrbank17_ev_status_w;
			end
			3'd4: begin
				interface17_bank_bus_dat_r <= csrbank17_ev_pending_w;
			end
			3'd5: begin
				interface17_bank_bus_dat_r <= csrbank17_ev_enable0_w;
			end
		endcase
	end
	gpioin4_in_re <= csrbank17_in_re;
	if (csrbank17_mode0_re) begin
		gpioin4_gpioin4_mode_storage <= csrbank17_mode0_r;
	end
	gpioin4_gpioin4_mode_re <= csrbank17_mode0_re;
	if (csrbank17_edge0_re) begin
		gpioin4_gpioin4_edge_storage <= csrbank17_edge0_r;
	end
	gpioin4_gpioin4_edge_re <= csrbank17_edge0_re;
	gpioin4_status_re <= csrbank17_ev_status_re;
	if (csrbank17_ev_pending_re) begin
		gpioin4_pending_r <= csrbank17_ev_pending_r;
	end
	gpioin4_pending_re <= csrbank17_ev_pending_re;
	if (csrbank17_ev_enable0_re) begin
		gpioin4_enable_storage <= csrbank17_ev_enable0_r;
	end
	gpioin4_enable_re <= csrbank17_ev_enable0_re;
	interface18_bank_bus_dat_r <= 1'd0;
	if (csrbank18_sel) begin
		case (interface18_bank_bus_adr[8:0])
			1'd0: begin
				interface18_bank_bus_dat_r <= csrbank18_in_w;
			end
			1'd1: begin
				interface18_bank_bus_dat_r <= csrbank18_mode0_w;
			end
			2'd2: begin
				interface18_bank_bus_dat_r <= csrbank18_edge0_w;
			end
			2'd3: begin
				interface18_bank_bus_dat_r <= csrbank18_ev_status_w;
			end
			3'd4: begin
				interface18_bank_bus_dat_r <= csrbank18_ev_pending_w;
			end
			3'd5: begin
				interface18_bank_bus_dat_r <= csrbank18_ev_enable0_w;
			end
		endcase
	end
	gpioin5_in_re <= csrbank18_in_re;
	if (csrbank18_mode0_re) begin
		gpioin5_gpioin5_mode_storage <= csrbank18_mode0_r;
	end
	gpioin5_gpioin5_mode_re <= csrbank18_mode0_re;
	if (csrbank18_edge0_re) begin
		gpioin5_gpioin5_edge_storage <= csrbank18_edge0_r;
	end
	gpioin5_gpioin5_edge_re <= csrbank18_edge0_re;
	gpioin5_status_re <= csrbank18_ev_status_re;
	if (csrbank18_ev_pending_re) begin
		gpioin5_pending_r <= csrbank18_ev_pending_r;
	end
	gpioin5_pending_re <= csrbank18_ev_pending_re;
	if (csrbank18_ev_enable0_re) begin
		gpioin5_enable_storage <= csrbank18_ev_enable0_r;
	end
	gpioin5_enable_re <= csrbank18_ev_enable0_re;
	interface19_bank_bus_dat_r <= 1'd0;
	if (csrbank19_sel) begin
		case (interface19_bank_bus_adr[8:0])
			1'd0: begin
				interface19_bank_bus_dat_r <= csrbank19_out0_w;
			end
		endcase
	end
	if (csrbank19_out0_re) begin
		user_irq_ena_storage[2:0] <= csrbank19_out0_r;
	end
	user_irq_ena_re <= csrbank19_out0_re;
	if (sys_rst) begin
	    // ****** added to correct GL testbench failure
        dbg_uart_tx_data <= 8'd0;
        dbg_uart_tx_count <= 4'd0;
        dbg_uart_tx_tick <= 1'd0;
        dbg_uart_tx_phase <= 32'd0;
        dbg_uart_rx_tick <= 1'd0;
        dbg_uart_rx_phase <= 32'd0;
        dbg_uart_rx_rx_d <= 1'd0;
        dbg_uart_cmd <= 8'd0;
        dbg_uart_incr <= 1'd0;
        dbg_uart_address <= 32'd0;
        dbg_uart_data <= 32'd0;
        dbg_uart_bytes_count <= 2'd0;
        dbg_uart_words_count <= 8'd0;
        dbg_uart_count <= 20'd1000000;
	    // ******
		mgmtsoc_reset_storage <= 2'd0;
		mgmtsoc_reset_re <= 1'd0;
		mgmtsoc_scratch_storage <= 32'd305419896;
		mgmtsoc_scratch_re <= 1'd0;
		mgmtsoc_bus_errors_re <= 1'd0;
		mgmtsoc_bus_errors <= 32'd0;
		mgmtsoc_vexriscv_debug_reset <= 1'd0;
		mgmtsoc_vexriscv_ibus_err <= 1'd0;
		mgmtsoc_vexriscv_dbus_err <= 1'd0;
		mgmtsoc_vexriscv_i_cmd_valid <= 1'd0;
		mgmtsoc_vexriscv_i_cmd_payload_wr <= 1'd0;
		mgmtsoc_vexriscv_i_cmd_payload_address <= 8'd0;
		mgmtsoc_vexriscv_i_cmd_payload_data <= 32'd0;
		mgmtsoc_vexriscv_reset_debug_logic <= 1'd0;
		mgmtsoc_vexriscv_transfer_complete <= 1'd0;
		mgmtsoc_vexriscv_transfer_in_progress <= 1'd0;
		mgmtsoc_vexriscv_transfer_wait_for_ack <= 1'd0;
		mgmtsoc_vexriscv_debug_bus_ack <= 1'd0;
		mgmtsoc_load_storage <= 32'd0;
		mgmtsoc_load_re <= 1'd0;
		mgmtsoc_reload_storage <= 32'd0;
		mgmtsoc_reload_re <= 1'd0;
		mgmtsoc_en_storage <= 1'd0;
		mgmtsoc_en_re <= 1'd0;
		mgmtsoc_update_value_storage <= 1'd0;
		mgmtsoc_update_value_re <= 1'd0;
		mgmtsoc_value_status <= 32'd0;
		mgmtsoc_value_re <= 1'd0;
		mgmtsoc_zero_pending <= 1'd0;
		mgmtsoc_zero_trigger_d <= 1'd0;
		mgmtsoc_status_re <= 1'd0;
		mgmtsoc_pending_re <= 1'd0;
		mgmtsoc_pending_r <= 1'd0;
		mgmtsoc_enable_storage <= 1'd0;
		mgmtsoc_enable_re <= 1'd0;
		mgmtsoc_value <= 32'd0;
		dff_bus_ack <= 1'd0;
		dff2_bus_ack <= 1'd0;
		mgmtsoc_litespisdrphycore_storage <= 8'd1;
		mgmtsoc_litespisdrphycore_re <= 1'd0;
		mgmtsoc_litespisdrphycore_cnt <= 8'd0;
		mgmtsoc_litespisdrphycore_clk <= 1'd0;
		mgmtsoc_litespisdrphycore_posedge_reg <= 1'd0;
		mgmtsoc_litespisdrphycore_posedge_reg2 <= 1'd0;
		mgmtsoc_litespisdrphycore_count <= 4'd11;
		mgmtsoc_litespimmap_burst_cs <= 1'd0;
		mgmtsoc_litespimmap_count <= 9'd256;
		mgmtsoc_litespimmap_storage <= 8'd0;
		mgmtsoc_litespimmap_re <= 1'd0;
		mgmtsoc_master_cs_storage <= 1'd0;
		mgmtsoc_master_cs_re <= 1'd0;
		mgmtsoc_master_phyconfig_storage <= 24'd0;
		mgmtsoc_master_phyconfig_re <= 1'd0;
		mgmtsoc_master_status_re <= 1'd0;
		mgmtsoc_master_tx_fifo_source_valid <= 1'd0;
		mgmtsoc_master_tx_fifo_source_payload_data <= 32'd0;
		mgmtsoc_master_tx_fifo_source_payload_len <= 6'd0;
		mgmtsoc_master_tx_fifo_source_payload_width <= 4'd0;
		mgmtsoc_master_tx_fifo_source_payload_mask <= 8'd0;
		mgmtsoc_master_rx_fifo_source_valid <= 1'd0;
		mgmtsoc_master_rx_fifo_source_payload_data <= 32'd0;
		spi_clk <= 1'd0;
		spi_cs_n <= 1'd0;
		spi_mosi <= 1'd0;
		spi_master_miso <= 8'd0;
		spi_master_control_storage <= 16'd0;
		spi_master_control_re <= 1'd0;
		spi_master_status_re <= 1'd0;
		spi_master_mosi_re <= 1'd0;
		spi_master_miso_re <= 1'd0;
		spi_master_cs_storage <= 17'd1;
		spi_master_cs_re <= 1'd0;
		spi_master_loopback_storage <= 1'd0;
		spi_master_loopback_re <= 1'd0;
		spi_master_count <= 3'd0;
		spi_master_clk_divider1 <= 16'd0;
		spi_master_mosi_data <= 8'd0;
		spi_master_mosi_sel <= 3'd0;
		spi_master_miso_data <= 8'd0;
		spimaster_storage <= 16'd100;
		spimaster_re <= 1'd0;
		mprj_wb_iena_storage <= 1'd0;
		mprj_wb_iena_re <= 1'd0;
		sys_uart_tx <= 1'd1;
		uart_phy_tx_tick <= 1'd0;
		uart_phy_rx_tick <= 1'd0;
		uart_phy_rx_rx_d <= 1'd0;
		uart_txfull_re <= 1'd0;
		uart_rxempty_re <= 1'd0;
		uart_tx_pending <= 1'd0;
		uart_tx_trigger_d <= 1'd0;
		uart_rx_pending <= 1'd0;
		uart_rx_trigger_d <= 1'd0;
		uart_status_re <= 1'd0;
		uart_pending_re <= 1'd0;
		uart_pending_r <= 2'd0;
		uart_enable_storage <= 2'd0;
		uart_enable_re <= 1'd0;
		uart_txempty_re <= 1'd0;
		uart_rxfull_re <= 1'd0;
		uart_tx_fifo_readable <= 1'd0;
		uart_tx_fifo_level0 <= 5'd0;
		uart_tx_fifo_produce <= 4'd0;
		uart_tx_fifo_consume <= 4'd0;
		uart_rx_fifo_readable <= 1'd0;
		uart_rx_fifo_level0 <= 5'd0;
		uart_rx_fifo_produce <= 4'd0;
		uart_rx_fifo_consume <= 4'd0;
		dbg_uart_dbg_uart_tx <= 1'd1;
		dbg_uart_tx_tick <= 1'd0;
		dbg_uart_rx_tick <= 1'd0;
		dbg_uart_rx_rx_d <= 1'd0;
		dbg_uart_incr <= 1'd0;
		dbg_uart_count <= 20'd1000000;
		debug_oeb_storage <= 1'd0;
		debug_oeb_re <= 1'd0;
		debug_mode_storage <= 1'd0;
		debug_mode_re <= 1'd0;
		uart_enabled_storage <= 1'd0;
		uart_enabled_re <= 1'd0;
		gpio_mode1_storage <= 1'd0;
		gpio_mode1_re <= 1'd0;
		gpio_mode0_storage <= 1'd0;
		gpio_mode0_re <= 1'd0;
		gpio_ien_storage <= 1'd0;
		gpio_ien_re <= 1'd0;
		gpio_oe_storage <= 1'd0;
		gpio_oe_re <= 1'd0;
		gpio_in_re <= 1'd0;
		gpio_out_storage <= 1'd0;
		gpio_out_re <= 1'd0;
		la_ien_storage <= 128'd0;
		la_ien_re <= 1'd0;
		la_oe_storage <= 128'd0;
		la_oe_re <= 1'd0;
		la_in_re <= 1'd0;
		la_out_storage <= 128'd0;
		la_out_re <= 1'd0;
		spi_enabled_storage <= 1'd0;
		spi_enabled_re <= 1'd0;
		user_irq_ena_storage <= 3'd0;
		user_irq_ena_re <= 1'd0;
		gpioin0_in_re <= 1'd0;
		gpioin0_gpioin0_mode_storage <= 1'd0;
		gpioin0_gpioin0_mode_re <= 1'd0;
		gpioin0_gpioin0_edge_storage <= 1'd0;
		gpioin0_gpioin0_edge_re <= 1'd0;
		gpioin0_gpioin0_in_pads_n_d <= 1'd0;
		gpioin0_gpioin0_pending <= 1'd0;
		gpioin0_gpioin0_trigger_d <= 1'd0;
		gpioin1_in_re <= 1'd0;
		gpioin1_gpioin1_mode_storage <= 1'd0;
		gpioin1_gpioin1_mode_re <= 1'd0;
		gpioin1_gpioin1_edge_storage <= 1'd0;
		gpioin1_gpioin1_edge_re <= 1'd0;
		gpioin1_gpioin1_in_pads_n_d <= 1'd0;
		gpioin1_gpioin1_pending <= 1'd0;
		gpioin1_gpioin1_trigger_d <= 1'd0;
		gpioin2_in_re <= 1'd0;
		gpioin2_gpioin2_mode_storage <= 1'd0;
		gpioin2_gpioin2_mode_re <= 1'd0;
		gpioin2_gpioin2_edge_storage <= 1'd0;
		gpioin2_gpioin2_edge_re <= 1'd0;
		gpioin2_gpioin2_in_pads_n_d <= 1'd0;
		gpioin2_gpioin2_pending <= 1'd0;
		gpioin2_gpioin2_trigger_d <= 1'd0;
		gpioin3_in_re <= 1'd0;
		gpioin3_gpioin3_mode_storage <= 1'd0;
		gpioin3_gpioin3_mode_re <= 1'd0;
		gpioin3_gpioin3_edge_storage <= 1'd0;
		gpioin3_gpioin3_edge_re <= 1'd0;
		gpioin3_gpioin3_in_pads_n_d <= 1'd0;
		gpioin3_gpioin3_pending <= 1'd0;
		gpioin3_gpioin3_trigger_d <= 1'd0;
		gpioin4_in_re <= 1'd0;
		gpioin4_gpioin4_mode_storage <= 1'd0;
		gpioin4_gpioin4_mode_re <= 1'd0;
		gpioin4_gpioin4_edge_storage <= 1'd0;
		gpioin4_gpioin4_edge_re <= 1'd0;
		gpioin4_gpioin4_in_pads_n_d <= 1'd0;
		gpioin4_gpioin4_pending <= 1'd0;
		gpioin4_gpioin4_trigger_d <= 1'd0;
		gpioin5_in_re <= 1'd0;
		gpioin5_gpioin5_mode_storage <= 1'd0;
		gpioin5_gpioin5_mode_re <= 1'd0;
		gpioin5_gpioin5_edge_storage <= 1'd0;
		gpioin5_gpioin5_edge_re <= 1'd0;
		gpioin5_gpioin5_in_pads_n_d <= 1'd0;
		gpioin5_gpioin5_pending <= 1'd0;
		gpioin5_gpioin5_trigger_d <= 1'd0;
		litespiphy_state <= 2'd0;
		litespi_grant <= 1'd0;
		litespi_state <= 4'd0;
		spimaster_state <= 2'd0;
		rs232phy_rs232phytx_state <= 1'd0;
		rs232phy_rs232phyrx_state <= 1'd0;
		uartwishbonebridge_rs232phytx_state <= 1'd0;
		uartwishbonebridge_rs232phyrx_state <= 1'd0;
		uartwishbonebridge_state <= 3'd0;
		gpioin0_status_re <= 1'd0;
		gpioin0_pending_re <= 1'd0;
		gpioin0_pending_r <= 1'd0;
		gpioin0_enable_storage <= 1'd0;
		gpioin0_enable_re <= 1'd0;
		gpioin1_status_re <= 1'd0;
		gpioin1_pending_re <= 1'd0;
		gpioin1_pending_r <= 1'd0;
		gpioin1_enable_storage <= 1'd0;
		gpioin1_enable_re <= 1'd0;
		gpioin2_status_re <= 1'd0;
		gpioin2_pending_re <= 1'd0;
		gpioin2_pending_r <= 1'd0;
		gpioin2_enable_storage <= 1'd0;
		gpioin2_enable_re <= 1'd0;
		gpioin3_status_re <= 1'd0;
		gpioin3_pending_re <= 1'd0;
		gpioin3_pending_r <= 1'd0;
		gpioin3_enable_storage <= 1'd0;
		gpioin3_enable_re <= 1'd0;
		gpioin4_status_re <= 1'd0;
		gpioin4_pending_re <= 1'd0;
		gpioin4_pending_r <= 1'd0;
		gpioin4_enable_storage <= 1'd0;
		gpioin4_enable_re <= 1'd0;
		gpioin5_status_re <= 1'd0;
		gpioin5_pending_re <= 1'd0;
		gpioin5_pending_r <= 1'd0;
		gpioin5_enable_storage <= 1'd0;
		gpioin5_enable_re <= 1'd0;
		grant <= 2'd0;
		slave_sel_r <= 7'd0;
		count <= 20'd1000000;
		state <= 1'd0;
	end
	multiregimpl0_regs0 <= sys_uart_rx;
	multiregimpl0_regs1 <= multiregimpl0_regs0;
	multiregimpl1_regs0 <= dbg_uart_dbg_uart_rx;
	multiregimpl1_regs1 <= multiregimpl1_regs0;
	multiregimpl2_regs0 <= gpio_in_pad;
	multiregimpl2_regs1 <= multiregimpl2_regs0;
	multiregimpl3_regs0 <= la_input[0];
	multiregimpl3_regs1 <= multiregimpl3_regs0;
	multiregimpl4_regs0 <= la_input[1];
	multiregimpl4_regs1 <= multiregimpl4_regs0;
	multiregimpl5_regs0 <= la_input[2];
	multiregimpl5_regs1 <= multiregimpl5_regs0;
	multiregimpl6_regs0 <= la_input[3];
	multiregimpl6_regs1 <= multiregimpl6_regs0;
	multiregimpl7_regs0 <= la_input[4];
	multiregimpl7_regs1 <= multiregimpl7_regs0;
	multiregimpl8_regs0 <= la_input[5];
	multiregimpl8_regs1 <= multiregimpl8_regs0;
	multiregimpl9_regs0 <= la_input[6];
	multiregimpl9_regs1 <= multiregimpl9_regs0;
	multiregimpl10_regs0 <= la_input[7];
	multiregimpl10_regs1 <= multiregimpl10_regs0;
	multiregimpl11_regs0 <= la_input[8];
	multiregimpl11_regs1 <= multiregimpl11_regs0;
	multiregimpl12_regs0 <= la_input[9];
	multiregimpl12_regs1 <= multiregimpl12_regs0;
	multiregimpl13_regs0 <= la_input[10];
	multiregimpl13_regs1 <= multiregimpl13_regs0;
	multiregimpl14_regs0 <= la_input[11];
	multiregimpl14_regs1 <= multiregimpl14_regs0;
	multiregimpl15_regs0 <= la_input[12];
	multiregimpl15_regs1 <= multiregimpl15_regs0;
	multiregimpl16_regs0 <= la_input[13];
	multiregimpl16_regs1 <= multiregimpl16_regs0;
	multiregimpl17_regs0 <= la_input[14];
	multiregimpl17_regs1 <= multiregimpl17_regs0;
	multiregimpl18_regs0 <= la_input[15];
	multiregimpl18_regs1 <= multiregimpl18_regs0;
	multiregimpl19_regs0 <= la_input[16];
	multiregimpl19_regs1 <= multiregimpl19_regs0;
	multiregimpl20_regs0 <= la_input[17];
	multiregimpl20_regs1 <= multiregimpl20_regs0;
	multiregimpl21_regs0 <= la_input[18];
	multiregimpl21_regs1 <= multiregimpl21_regs0;
	multiregimpl22_regs0 <= la_input[19];
	multiregimpl22_regs1 <= multiregimpl22_regs0;
	multiregimpl23_regs0 <= la_input[20];
	multiregimpl23_regs1 <= multiregimpl23_regs0;
	multiregimpl24_regs0 <= la_input[21];
	multiregimpl24_regs1 <= multiregimpl24_regs0;
	multiregimpl25_regs0 <= la_input[22];
	multiregimpl25_regs1 <= multiregimpl25_regs0;
	multiregimpl26_regs0 <= la_input[23];
	multiregimpl26_regs1 <= multiregimpl26_regs0;
	multiregimpl27_regs0 <= la_input[24];
	multiregimpl27_regs1 <= multiregimpl27_regs0;
	multiregimpl28_regs0 <= la_input[25];
	multiregimpl28_regs1 <= multiregimpl28_regs0;
	multiregimpl29_regs0 <= la_input[26];
	multiregimpl29_regs1 <= multiregimpl29_regs0;
	multiregimpl30_regs0 <= la_input[27];
	multiregimpl30_regs1 <= multiregimpl30_regs0;
	multiregimpl31_regs0 <= la_input[28];
	multiregimpl31_regs1 <= multiregimpl31_regs0;
	multiregimpl32_regs0 <= la_input[29];
	multiregimpl32_regs1 <= multiregimpl32_regs0;
	multiregimpl33_regs0 <= la_input[30];
	multiregimpl33_regs1 <= multiregimpl33_regs0;
	multiregimpl34_regs0 <= la_input[31];
	multiregimpl34_regs1 <= multiregimpl34_regs0;
	multiregimpl35_regs0 <= la_input[32];
	multiregimpl35_regs1 <= multiregimpl35_regs0;
	multiregimpl36_regs0 <= la_input[33];
	multiregimpl36_regs1 <= multiregimpl36_regs0;
	multiregimpl37_regs0 <= la_input[34];
	multiregimpl37_regs1 <= multiregimpl37_regs0;
	multiregimpl38_regs0 <= la_input[35];
	multiregimpl38_regs1 <= multiregimpl38_regs0;
	multiregimpl39_regs0 <= la_input[36];
	multiregimpl39_regs1 <= multiregimpl39_regs0;
	multiregimpl40_regs0 <= la_input[37];
	multiregimpl40_regs1 <= multiregimpl40_regs0;
	multiregimpl41_regs0 <= la_input[38];
	multiregimpl41_regs1 <= multiregimpl41_regs0;
	multiregimpl42_regs0 <= la_input[39];
	multiregimpl42_regs1 <= multiregimpl42_regs0;
	multiregimpl43_regs0 <= la_input[40];
	multiregimpl43_regs1 <= multiregimpl43_regs0;
	multiregimpl44_regs0 <= la_input[41];
	multiregimpl44_regs1 <= multiregimpl44_regs0;
	multiregimpl45_regs0 <= la_input[42];
	multiregimpl45_regs1 <= multiregimpl45_regs0;
	multiregimpl46_regs0 <= la_input[43];
	multiregimpl46_regs1 <= multiregimpl46_regs0;
	multiregimpl47_regs0 <= la_input[44];
	multiregimpl47_regs1 <= multiregimpl47_regs0;
	multiregimpl48_regs0 <= la_input[45];
	multiregimpl48_regs1 <= multiregimpl48_regs0;
	multiregimpl49_regs0 <= la_input[46];
	multiregimpl49_regs1 <= multiregimpl49_regs0;
	multiregimpl50_regs0 <= la_input[47];
	multiregimpl50_regs1 <= multiregimpl50_regs0;
	multiregimpl51_regs0 <= la_input[48];
	multiregimpl51_regs1 <= multiregimpl51_regs0;
	multiregimpl52_regs0 <= la_input[49];
	multiregimpl52_regs1 <= multiregimpl52_regs0;
	multiregimpl53_regs0 <= la_input[50];
	multiregimpl53_regs1 <= multiregimpl53_regs0;
	multiregimpl54_regs0 <= la_input[51];
	multiregimpl54_regs1 <= multiregimpl54_regs0;
	multiregimpl55_regs0 <= la_input[52];
	multiregimpl55_regs1 <= multiregimpl55_regs0;
	multiregimpl56_regs0 <= la_input[53];
	multiregimpl56_regs1 <= multiregimpl56_regs0;
	multiregimpl57_regs0 <= la_input[54];
	multiregimpl57_regs1 <= multiregimpl57_regs0;
	multiregimpl58_regs0 <= la_input[55];
	multiregimpl58_regs1 <= multiregimpl58_regs0;
	multiregimpl59_regs0 <= la_input[56];
	multiregimpl59_regs1 <= multiregimpl59_regs0;
	multiregimpl60_regs0 <= la_input[57];
	multiregimpl60_regs1 <= multiregimpl60_regs0;
	multiregimpl61_regs0 <= la_input[58];
	multiregimpl61_regs1 <= multiregimpl61_regs0;
	multiregimpl62_regs0 <= la_input[59];
	multiregimpl62_regs1 <= multiregimpl62_regs0;
	multiregimpl63_regs0 <= la_input[60];
	multiregimpl63_regs1 <= multiregimpl63_regs0;
	multiregimpl64_regs0 <= la_input[61];
	multiregimpl64_regs1 <= multiregimpl64_regs0;
	multiregimpl65_regs0 <= la_input[62];
	multiregimpl65_regs1 <= multiregimpl65_regs0;
	multiregimpl66_regs0 <= la_input[63];
	multiregimpl66_regs1 <= multiregimpl66_regs0;
	multiregimpl67_regs0 <= la_input[64];
	multiregimpl67_regs1 <= multiregimpl67_regs0;
	multiregimpl68_regs0 <= la_input[65];
	multiregimpl68_regs1 <= multiregimpl68_regs0;
	multiregimpl69_regs0 <= la_input[66];
	multiregimpl69_regs1 <= multiregimpl69_regs0;
	multiregimpl70_regs0 <= la_input[67];
	multiregimpl70_regs1 <= multiregimpl70_regs0;
	multiregimpl71_regs0 <= la_input[68];
	multiregimpl71_regs1 <= multiregimpl71_regs0;
	multiregimpl72_regs0 <= la_input[69];
	multiregimpl72_regs1 <= multiregimpl72_regs0;
	multiregimpl73_regs0 <= la_input[70];
	multiregimpl73_regs1 <= multiregimpl73_regs0;
	multiregimpl74_regs0 <= la_input[71];
	multiregimpl74_regs1 <= multiregimpl74_regs0;
	multiregimpl75_regs0 <= la_input[72];
	multiregimpl75_regs1 <= multiregimpl75_regs0;
	multiregimpl76_regs0 <= la_input[73];
	multiregimpl76_regs1 <= multiregimpl76_regs0;
	multiregimpl77_regs0 <= la_input[74];
	multiregimpl77_regs1 <= multiregimpl77_regs0;
	multiregimpl78_regs0 <= la_input[75];
	multiregimpl78_regs1 <= multiregimpl78_regs0;
	multiregimpl79_regs0 <= la_input[76];
	multiregimpl79_regs1 <= multiregimpl79_regs0;
	multiregimpl80_regs0 <= la_input[77];
	multiregimpl80_regs1 <= multiregimpl80_regs0;
	multiregimpl81_regs0 <= la_input[78];
	multiregimpl81_regs1 <= multiregimpl81_regs0;
	multiregimpl82_regs0 <= la_input[79];
	multiregimpl82_regs1 <= multiregimpl82_regs0;
	multiregimpl83_regs0 <= la_input[80];
	multiregimpl83_regs1 <= multiregimpl83_regs0;
	multiregimpl84_regs0 <= la_input[81];
	multiregimpl84_regs1 <= multiregimpl84_regs0;
	multiregimpl85_regs0 <= la_input[82];
	multiregimpl85_regs1 <= multiregimpl85_regs0;
	multiregimpl86_regs0 <= la_input[83];
	multiregimpl86_regs1 <= multiregimpl86_regs0;
	multiregimpl87_regs0 <= la_input[84];
	multiregimpl87_regs1 <= multiregimpl87_regs0;
	multiregimpl88_regs0 <= la_input[85];
	multiregimpl88_regs1 <= multiregimpl88_regs0;
	multiregimpl89_regs0 <= la_input[86];
	multiregimpl89_regs1 <= multiregimpl89_regs0;
	multiregimpl90_regs0 <= la_input[87];
	multiregimpl90_regs1 <= multiregimpl90_regs0;
	multiregimpl91_regs0 <= la_input[88];
	multiregimpl91_regs1 <= multiregimpl91_regs0;
	multiregimpl92_regs0 <= la_input[89];
	multiregimpl92_regs1 <= multiregimpl92_regs0;
	multiregimpl93_regs0 <= la_input[90];
	multiregimpl93_regs1 <= multiregimpl93_regs0;
	multiregimpl94_regs0 <= la_input[91];
	multiregimpl94_regs1 <= multiregimpl94_regs0;
	multiregimpl95_regs0 <= la_input[92];
	multiregimpl95_regs1 <= multiregimpl95_regs0;
	multiregimpl96_regs0 <= la_input[93];
	multiregimpl96_regs1 <= multiregimpl96_regs0;
	multiregimpl97_regs0 <= la_input[94];
	multiregimpl97_regs1 <= multiregimpl97_regs0;
	multiregimpl98_regs0 <= la_input[95];
	multiregimpl98_regs1 <= multiregimpl98_regs0;
	multiregimpl99_regs0 <= la_input[96];
	multiregimpl99_regs1 <= multiregimpl99_regs0;
	multiregimpl100_regs0 <= la_input[97];
	multiregimpl100_regs1 <= multiregimpl100_regs0;
	multiregimpl101_regs0 <= la_input[98];
	multiregimpl101_regs1 <= multiregimpl101_regs0;
	multiregimpl102_regs0 <= la_input[99];
	multiregimpl102_regs1 <= multiregimpl102_regs0;
	multiregimpl103_regs0 <= la_input[100];
	multiregimpl103_regs1 <= multiregimpl103_regs0;
	multiregimpl104_regs0 <= la_input[101];
	multiregimpl104_regs1 <= multiregimpl104_regs0;
	multiregimpl105_regs0 <= la_input[102];
	multiregimpl105_regs1 <= multiregimpl105_regs0;
	multiregimpl106_regs0 <= la_input[103];
	multiregimpl106_regs1 <= multiregimpl106_regs0;
	multiregimpl107_regs0 <= la_input[104];
	multiregimpl107_regs1 <= multiregimpl107_regs0;
	multiregimpl108_regs0 <= la_input[105];
	multiregimpl108_regs1 <= multiregimpl108_regs0;
	multiregimpl109_regs0 <= la_input[106];
	multiregimpl109_regs1 <= multiregimpl109_regs0;
	multiregimpl110_regs0 <= la_input[107];
	multiregimpl110_regs1 <= multiregimpl110_regs0;
	multiregimpl111_regs0 <= la_input[108];
	multiregimpl111_regs1 <= multiregimpl111_regs0;
	multiregimpl112_regs0 <= la_input[109];
	multiregimpl112_regs1 <= multiregimpl112_regs0;
	multiregimpl113_regs0 <= la_input[110];
	multiregimpl113_regs1 <= multiregimpl113_regs0;
	multiregimpl114_regs0 <= la_input[111];
	multiregimpl114_regs1 <= multiregimpl114_regs0;
	multiregimpl115_regs0 <= la_input[112];
	multiregimpl115_regs1 <= multiregimpl115_regs0;
	multiregimpl116_regs0 <= la_input[113];
	multiregimpl116_regs1 <= multiregimpl116_regs0;
	multiregimpl117_regs0 <= la_input[114];
	multiregimpl117_regs1 <= multiregimpl117_regs0;
	multiregimpl118_regs0 <= la_input[115];
	multiregimpl118_regs1 <= multiregimpl118_regs0;
	multiregimpl119_regs0 <= la_input[116];
	multiregimpl119_regs1 <= multiregimpl119_regs0;
	multiregimpl120_regs0 <= la_input[117];
	multiregimpl120_regs1 <= multiregimpl120_regs0;
	multiregimpl121_regs0 <= la_input[118];
	multiregimpl121_regs1 <= multiregimpl121_regs0;
	multiregimpl122_regs0 <= la_input[119];
	multiregimpl122_regs1 <= multiregimpl122_regs0;
	multiregimpl123_regs0 <= la_input[120];
	multiregimpl123_regs1 <= multiregimpl123_regs0;
	multiregimpl124_regs0 <= la_input[121];
	multiregimpl124_regs1 <= multiregimpl124_regs0;
	multiregimpl125_regs0 <= la_input[122];
	multiregimpl125_regs1 <= multiregimpl125_regs0;
	multiregimpl126_regs0 <= la_input[123];
	multiregimpl126_regs1 <= multiregimpl126_regs0;
	multiregimpl127_regs0 <= la_input[124];
	multiregimpl127_regs1 <= multiregimpl127_regs0;
	multiregimpl128_regs0 <= la_input[125];
	multiregimpl128_regs1 <= multiregimpl128_regs0;
	multiregimpl129_regs0 <= la_input[126];
	multiregimpl129_regs1 <= multiregimpl129_regs0;
	multiregimpl130_regs0 <= la_input[127];
	multiregimpl130_regs1 <= multiregimpl130_regs0;
	multiregimpl131_regs0 <= user_irq[0];
	multiregimpl131_regs1 <= multiregimpl131_regs0;
	multiregimpl132_regs0 <= user_irq[1];
	multiregimpl132_regs1 <= multiregimpl132_regs0;
	multiregimpl133_regs0 <= user_irq[2];
	multiregimpl133_regs1 <= multiregimpl133_regs0;
	multiregimpl134_regs0 <= user_irq[3];
	multiregimpl134_regs1 <= multiregimpl134_regs0;
	multiregimpl135_regs0 <= user_irq[4];
	multiregimpl135_regs1 <= multiregimpl135_regs0;
	multiregimpl136_regs0 <= user_irq[5];
	multiregimpl136_regs1 <= multiregimpl136_regs0;
end

RAM256 RAM256(
	.A0(dff_bus_adr[7:0]),
	.CLK(sys_clk),
	.Di0(dff_di),
	.EN0(dff_en),
	.WE0(dff_we),
	.Do0(dff_do)
);

RAM128 RAM128(
	.A0(dff2_bus_adr[6:0]),
	.CLK(sys_clk),
	.Di0(dff2_di),
	.EN0(dff2_en),
	.WE0(dff2_we),
	.Do0(dff2_do)
);

reg [9:0] storage[0:15];
reg [9:0] memdat;
reg [9:0] memdat_1;
always @(posedge sys_clk) begin
	if (uart_tx_fifo_wrport_we)
		storage[uart_tx_fifo_wrport_adr] <= uart_tx_fifo_wrport_dat_w;
	memdat <= storage[uart_tx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
	if (uart_tx_fifo_rdport_re)
		memdat_1 <= storage[uart_tx_fifo_rdport_adr];
end

assign uart_tx_fifo_wrport_dat_r = memdat;
assign uart_tx_fifo_rdport_dat_r = memdat_1;

reg [9:0] storage_1[0:15];
reg [9:0] memdat_2;
reg [9:0] memdat_3;
always @(posedge sys_clk) begin
	if (uart_rx_fifo_wrport_we)
		storage_1[uart_rx_fifo_wrport_adr] <= uart_rx_fifo_wrport_dat_w;
	memdat_2 <= storage_1[uart_rx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
	if (uart_rx_fifo_rdport_re)
		memdat_3 <= storage_1[uart_rx_fifo_rdport_adr];
end

assign uart_rx_fifo_wrport_dat_r = memdat_2;
assign uart_rx_fifo_rdport_dat_r = memdat_3;

VexRiscv VexRiscv(
	.clk(sys_clk),
	.dBusWishbone_ACK(mgmtsoc_dbus_dbus_ack),
	.dBusWishbone_DAT_MISO(mgmtsoc_dbus_dbus_dat_r),
	.dBusWishbone_ERR((mgmtsoc_dbus_dbus_err | mgmtsoc_vexriscv_dbus_err)),
	.debugReset(sys_rst),
	.debug_bus_cmd_payload_address(mgmtsoc_vexriscv_i_cmd_payload_address),
	.debug_bus_cmd_payload_data(mgmtsoc_vexriscv_i_cmd_payload_data),
	.debug_bus_cmd_payload_wr(mgmtsoc_vexriscv_i_cmd_payload_wr),
	.debug_bus_cmd_valid(mgmtsoc_vexriscv_i_cmd_valid),
	.externalInterruptArray(mgmtsoc_interrupt),
	.externalResetVector(mgmtsoc_vexriscv),
	.iBusWishbone_ACK(mgmtsoc_ibus_ibus_ack),
	.iBusWishbone_DAT_MISO(mgmtsoc_ibus_ibus_dat_r),
	.iBusWishbone_ERR((mgmtsoc_ibus_ibus_err | mgmtsoc_vexriscv_ibus_err)),
	.reset(((sys_rst | mgmtsoc_reset) | mgmtsoc_vexriscv_debug_reset)),
	.softwareInterrupt(1'd0),
	.timerInterrupt(1'd0),
	.dBusWishbone_ADR(mgmtsoc_dbus_dbus_adr),
	.dBusWishbone_BTE(mgmtsoc_dbus_dbus_bte),
	.dBusWishbone_CTI(mgmtsoc_dbus_dbus_cti),
	.dBusWishbone_CYC(mgmtsoc_dbus_dbus_cyc),
	.dBusWishbone_DAT_MOSI(mgmtsoc_dbus_dbus_dat_w),
	.dBusWishbone_SEL(mgmtsoc_dbus_dbus_sel),
	.dBusWishbone_STB(mgmtsoc_dbus_dbus_stb),
	.dBusWishbone_WE(mgmtsoc_dbus_dbus_we),
	.debug_bus_cmd_ready(mgmtsoc_vexriscv_o_cmd_ready),
	.debug_bus_rsp_data(mgmtsoc_vexriscv_o_rsp_data),
	.debug_resetOut(mgmtsoc_vexriscv_o_resetOut),
	.iBusWishbone_ADR(mgmtsoc_ibus_ibus_adr),
	.iBusWishbone_BTE(mgmtsoc_ibus_ibus_bte),
	.iBusWishbone_CTI(mgmtsoc_ibus_ibus_cti),
	.iBusWishbone_CYC(mgmtsoc_ibus_ibus_cyc),
	.iBusWishbone_DAT_MOSI(mgmtsoc_ibus_ibus_dat_w),
	.iBusWishbone_SEL(mgmtsoc_ibus_ibus_sel),
	.iBusWishbone_STB(mgmtsoc_ibus_ibus_stb),
	.iBusWishbone_WE(mgmtsoc_ibus_ibus_we)
);

endmodule
/*
 *  SPDX-FileCopyrightText: 2015 Clifford Wolf
 *  PicoSoC - A simple example SoC using PicoRV32
 *
 *  Copyright (C) 2017  Clifford Wolf <clifford@clifford.at>
 *
 *  Permission to use, copy, modify, and/or distribute this software for any
 *  purpose with or without fee is hereby granted, provided that the above
 *  copyright notice and this permission notice appear in all copies.
 *
 *  THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
 *  WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
 *  MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
 *  ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
 *  WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
 *  ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
 *  OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 *
 *  Revision 1,  July 2019:  Added signals to drive flash_clk and flash_csb
 *  output enable (inverted), tied to reset so that the flash is completely
 *  isolated from the processor when the processor is in reset.
 *
 *  Also: Made ram_wenb a 4-bit bus so that the memory access can be made
 *  byte-wide for byte-wide instructions.
 *
 *  SPDX-License-Identifier: ISC
 */


//`default_nettype none



/* Wrapper module around management SoC core for pin compatibility  */
/* with the Caravel harness chip. */    

module mgmt_core_wrapper (
    // Clock and reset
    input core_clk,
    input core_rstn,

    // Pass-thru signals
    input clk_in,
    input resetn_in,
    output clk_out,
    output resetn_out,

    input serial_load_in,
    input serial_data_2_in,
    input serial_resetn_in,
    input serial_clock_in,
    input rstb_l_in,
    //input por_l_in,
    //input porb_h_in,

    output serial_load_out,
    output serial_data_2_out,
    output serial_resetn_out,
    output serial_clock_out,
    output rstb_l_out,
    //output por_l_out,
    //output porb_h_out,

    // GPIO (one pin)
    output gpio_out_pad,    // Connect to out on gpio pad
    input  gpio_in_pad,     // Connect to in on gpio pad
    output gpio_mode0_pad,  // Connect to dm[0] on gpio pad
    output gpio_mode1_pad,  // Connect to dm[2] on gpio pad
    output gpio_outenb_pad, // Connect to oe_n on gpio pad
    output gpio_inenb_pad,  // Connect to inp_dis on gpio pad

    // Logic analyzer signals
    input  [127:0] la_input,            // From user project to CPU
    output [127:0] la_output,           // From CPU to user project
    output [127:0] la_oenb,             // Logic analyzer output enable
    output [127:0] la_iena,             // Logic analyzer input enable

    // Flash memory control (SPI master)
    output flash_csb,
    output flash_clk,

    output flash_io0_oeb,
    output flash_io1_oeb,
    output flash_io2_oeb,
    output flash_io3_oeb,

    output flash_io0_do,
    output flash_io1_do,
    output flash_io2_do,
    output flash_io3_do,

    input  flash_io0_di,
    input  flash_io1_di,
    input  flash_io2_di,
    input  flash_io3_di,

    // Exported Wishboned bus
    output    mprj_wb_iena, // Enable for the user wishbone return signals
    output    mprj_cyc_o,
    output    mprj_stb_o,
    output    mprj_we_o,
    output [3:0]  mprj_sel_o,
    output [31:0] mprj_adr_o,
    output [31:0] mprj_dat_o,
    input     mprj_ack_i,
    input  [31:0] mprj_dat_i,

    output    hk_cyc_o,
    output    hk_stb_o,
    input  [31:0] hk_dat_i,
    input     hk_ack_i,

    // IRQ
    input  [5:0] irq,       // IRQ from SPI and user project
    output [2:0] user_irq_ena,  // Enables for user project IRQ

    // Module status
    output qspi_enabled,
    output uart_enabled,
    output spi_enabled,
    output debug_mode,

    // Module I/O
    output ser_tx,
    input  ser_rx,
    output spi_csb,
    output spi_sck,
    output spi_sdo,
    output spi_sdoenb,
    input  spi_sdi,
    input  debug_in,
    output debug_out,
    output debug_oeb,

    // Trap state from CPU
    output trap
);


// Signals below are sram_ro ports that left no_connect
// as they are tied down inside mgmt_core

    /* Implement the PicoSoC core */

    mgmt_core core (
        .core_clk(core_clk),
        .core_rstn(core_rstn),

        // Pass-thru signals
        .clk_in(clk_in),
        .clk_out(clk_out),
        .resetn_in(resetn_in),
        .resetn_out(resetn_out),

        .serial_load_in(serial_load_in),
        .serial_load_out(serial_load_out),
        .serial_data_2_in(serial_data_2_in),
        .serial_data_2_out(serial_data_2_out),
        .serial_resetn_in(serial_resetn_in),
        .serial_resetn_out(serial_resetn_out),
        .serial_clock_in(serial_clock_in),
        .serial_clock_out(serial_clock_out),

        .rstb_l_in(rstb_l_in),
        .rstb_l_out(rstb_l_out),
        // [Vic]: POR is useless here
        //.por_l_in(por_l_in),
        //.por_l_out(por_l_out),
        //.porb_h_in(porb_h_in),
        //.porb_h_out(porb_h_out),

        // Trap state from CPU
        .trap(trap),

        // GPIO (one pin)
        .gpio_out_pad(gpio_out_pad),        // Connect to out on gpio pad
        .gpio_in_pad(gpio_in_pad),      // Connect to in on gpio pad
        .gpio_mode0_pad(gpio_mode0_pad),    // Connect to dm[0] on gpio pad
        .gpio_mode1_pad(gpio_mode1_pad),    // Connect to dm[2] on gpio pad
        .gpio_outenb_pad(gpio_outenb_pad),  // Connect to oe_n on gpio pad
        .gpio_inenb_pad(gpio_inenb_pad),    // Connect to inp_dis on gpio pad

        .la_input(la_input),            // From user project to CPU
        .la_output(la_output),          // From CPU to user project
        .la_oenb(la_oenb),          // Logic analyzer output enable
        .la_iena(la_iena),          // Logic analyzer input enable

        // IRQ
        .user_irq(irq),     // IRQ from SPI and user project
        .user_irq_ena(user_irq_ena),

        // Flash memory control (SPI master)
        .flash_cs_n(flash_csb),
        .flash_clk(flash_clk),

        .flash_io0_oeb(flash_io0_oeb),
        .flash_io1_oeb(flash_io1_oeb),
        .flash_io2_oeb(flash_io2_oeb),
        .flash_io3_oeb(flash_io3_oeb),

        .flash_io0_do(flash_io0_do),
        .flash_io1_do(flash_io1_do),
        .flash_io2_do(flash_io2_do),
        .flash_io3_do(flash_io3_do),

        .flash_io0_di(flash_io0_di),
        .flash_io1_di(flash_io1_di),
        .flash_io2_di(flash_io2_di),
        .flash_io3_di(flash_io3_di),

        // Exported wishbone bus (User project)
        .mprj_wb_iena(mprj_wb_iena),
        .mprj_ack_i(mprj_ack_i),
        .mprj_dat_i(mprj_dat_i),
        .mprj_cyc_o(mprj_cyc_o),
        .mprj_stb_o(mprj_stb_o),
        .mprj_we_o(mprj_we_o),
        .mprj_sel_o(mprj_sel_o),
        .mprj_adr_o(mprj_adr_o),
        .mprj_dat_o(mprj_dat_o),

        .hk_cyc_o(hk_cyc_o),
        .hk_stb_o(hk_stb_o),
        .hk_dat_i(hk_dat_i),
        .hk_ack_i(hk_ack_i),

        // Module status
        .qspi_enabled(qspi_enabled),
        .uart_enabled(uart_enabled),
        .spi_enabled(spi_enabled),
        .debug_mode(debug_mode),

        // Module I/O
//      .ser_tx(ser_tx),
//      .ser_rx(ser_rx),
        .serial_tx(ser_tx),
        .serial_rx(ser_rx),
        .spi_cs_n(spi_csb),
        .spi_clk(spi_sck),
        .spi_miso(spi_sdi),
        .spi_sdoenb(spi_sdoenb),
        .spi_mosi(spi_sdo),
        .debug_in(debug_in),
        .debug_out(debug_out),
        .debug_oeb(debug_oeb)

    );


endmodule
//`default_nettype wire



/* Copyright (C) 1991-2020 Free Software Foundation, Inc.
   This file is part of the GNU C Library.

   The GNU C Library is free software; you can redistribute it and/or
   modify it under the terms of the GNU Lesser General Public
   License as published by the Free Software Foundation; either
   version 2.1 of the License, or (at your option) any later version.

   The GNU C Library is distributed in the hope that it will be useful,
   but WITHOUT ANY WARRANTY; without even the implied warranty of
   MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
   Lesser General Public License for more details.

   You should have received a copy of the GNU Lesser General Public
   License along with the GNU C Library; if not, see
   <https://www.gnu.org/licenses/>.  */




/* This header is separate from features.h so that the compiler can
   include it implicitly at the start of every compilation.  It must
   not itself include <features.h> or any other header that includes
   <features.h> because the implicit include comes before any feature
   test macros that may be defined in a source file before it first
   explicitly includes a system header.  GCC knows the name of this
   header in order to preinclude it.  */

/* glibc's intent is to support the IEC 559 math functionality, real
   and complex.  If the GCC (4.9 and later) predefined macros
   specifying compiler intent are available, use them to determine
   whether the overall intent is to support these features; otherwise,
   presume an older compiler has intent to support these features and
   define these macros by default.  */
/* wchar_t uses Unicode 10.0.0.  Version 10.0 of the Unicode Standard is
   synchronized with ISO/IEC 10646:2017, fifth edition, plus
   the following additions from Amendment 1 to the fifth edition:
   - 56 emoji characters
   - 285 hentaigana
   - 3 additional Zanabazar Square characters */

// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

// `default_nettype none

/* Define the array of GPIO pads.  Note that the analog project support
 * version of caravel (caravan) defines fewer GPIO and replaces them
 * with analog in the chip_io_alt module.  Because the pad signalling
 * remains the same, `MPRJ_IO_PADS does not change, so a local parameter
 * is made that can be made smaller than `MPRJ_IO_PADS to accommodate
 * the analog pads.
 */

module mprj_io #(
    parameter AREA1PADS = `MPRJ_IO_PADS_1,
    parameter TOTAL_PADS = `MPRJ_IO_PADS
) (
    inout vddio,
    inout vssio,
    inout vdda,
    inout vssa,
    inout vccd,
    inout vssd,

    inout vdda1,
    inout vdda2,
    inout vssa1,
    inout vssa2,

    input vddio_q,
    input vssio_q,
    input analog_a,
    input analog_b,
    input porb_h,
    input [TOTAL_PADS-1:0] vccd_conb,
    inout [TOTAL_PADS-1:0] io,
    input [TOTAL_PADS-1:0] io_out,
    input [TOTAL_PADS-1:0] oeb,
    input [TOTAL_PADS-1:0] enh,
    input [TOTAL_PADS-1:0] inp_dis,
    input [TOTAL_PADS-1:0] ib_mode_sel,
    input [TOTAL_PADS-1:0] vtrip_sel,
    input [TOTAL_PADS-1:0] slow_sel,
    input [TOTAL_PADS-1:0] holdover,
    input [TOTAL_PADS-1:0] analog_en,
    input [TOTAL_PADS-1:0] analog_sel,
    input [TOTAL_PADS-1:0] analog_pol,
    input [TOTAL_PADS*3-1:0] dm,
    output [TOTAL_PADS-1:0] io_in,
    output [TOTAL_PADS-1:0] io_in_3v3,
    inout [TOTAL_PADS-10:0] analog_io,
    inout [TOTAL_PADS-10:0] analog_noesd_io
);

    wire [TOTAL_PADS-1:0] loop0_io; // Internal loopback to 3.3V domain ground
    wire [TOTAL_PADS-1:0] loop1_io; // Internal loopback to 3.3V domain power
    wire [6:0] no_connect_1a, no_connect_1b;
    wire [1:0] no_connect_2a, no_connect_2b;
boledu_io io_pad[TOTAL_PADS -1: 0] (
 .io(io[TOTAL_PADS-1:0]),
 .io_out (io_out[TOTAL_PADS - 1:0]),
 .oeb( oeb[TOTAL_PADS-1:0]),
 .io_in ( io_in[TOTAL_PADS-1:0])
);


endmodule


module boledu_io( inout io,
       input io_out,
       input oeb,
   output io_in);
 // bufif0(io_in, io, oeb);
 assign io_in = io;
 bufif0(io, io_out, oeb);
 //pullup (io);

endmodule


// `default_nettype wire
// Generator : SpinalHDL v1.6.0    git head : 73c8d8e2b86b45646e9d0b2e729291f2b65e6be3
// Component : VexRiscv
// Git hash  : c4eca1837ebca20b637a0a61e3a93d9446488459


`define EnvCtrlEnum_binary_sequential_type [1:0]
`define EnvCtrlEnum_binary_sequential_NONE 2'b00
`define EnvCtrlEnum_binary_sequential_XRET 2'b01
`define EnvCtrlEnum_binary_sequential_ECALL 2'b10

`define BranchCtrlEnum_binary_sequential_type [1:0]
`define BranchCtrlEnum_binary_sequential_INC 2'b00
`define BranchCtrlEnum_binary_sequential_B 2'b01
`define BranchCtrlEnum_binary_sequential_JAL 2'b10
`define BranchCtrlEnum_binary_sequential_JALR 2'b11

`define ShiftCtrlEnum_binary_sequential_type [1:0]
`define ShiftCtrlEnum_binary_sequential_DISABLE_1 2'b00
`define ShiftCtrlEnum_binary_sequential_SLL_1 2'b01
`define ShiftCtrlEnum_binary_sequential_SRL_1 2'b10
`define ShiftCtrlEnum_binary_sequential_SRA_1 2'b11

`define AluBitwiseCtrlEnum_binary_sequential_type [1:0]
`define AluBitwiseCtrlEnum_binary_sequential_XOR_1 2'b00
`define AluBitwiseCtrlEnum_binary_sequential_OR_1 2'b01
`define AluBitwiseCtrlEnum_binary_sequential_AND_1 2'b10

`define Src2CtrlEnum_binary_sequential_type [1:0]
`define Src2CtrlEnum_binary_sequential_RS 2'b00
`define Src2CtrlEnum_binary_sequential_IMI 2'b01
`define Src2CtrlEnum_binary_sequential_IMS 2'b10
`define Src2CtrlEnum_binary_sequential_PC 2'b11

`define AluCtrlEnum_binary_sequential_type [1:0]
`define AluCtrlEnum_binary_sequential_ADD_SUB 2'b00
`define AluCtrlEnum_binary_sequential_SLT_SLTU 2'b01
`define AluCtrlEnum_binary_sequential_BITWISE 2'b10

`define Src1CtrlEnum_binary_sequential_type [1:0]
`define Src1CtrlEnum_binary_sequential_RS 2'b00
`define Src1CtrlEnum_binary_sequential_IMU 2'b01
`define Src1CtrlEnum_binary_sequential_PC_INCREMENT 2'b10
`define Src1CtrlEnum_binary_sequential_URS1 2'b11


module VexRiscv (

  input      [31:0]   externalResetVector,
  input               timerInterrupt,
  input               softwareInterrupt,
  input      [31:0]   externalInterruptArray,
  input               debug_bus_cmd_valid,
  output reg          debug_bus_cmd_ready,
  input               debug_bus_cmd_payload_wr,
  input      [7:0]    debug_bus_cmd_payload_address,
  input      [31:0]   debug_bus_cmd_payload_data,
  output reg [31:0]   debug_bus_rsp_data,
  output              debug_resetOut,
  output reg          iBusWishbone_CYC,
  output reg          iBusWishbone_STB,
  input               iBusWishbone_ACK,
  output              iBusWishbone_WE,
  output     [29:0]   iBusWishbone_ADR,
  input      [31:0]   iBusWishbone_DAT_MISO,
  output     [31:0]   iBusWishbone_DAT_MOSI,
  output     [3:0]    iBusWishbone_SEL,
  input               iBusWishbone_ERR,
  output     [2:0]    iBusWishbone_CTI,
  output     [1:0]    iBusWishbone_BTE,
  output              dBusWishbone_CYC,
  output              dBusWishbone_STB,
  input               dBusWishbone_ACK,
  output              dBusWishbone_WE,
  output     [29:0]   dBusWishbone_ADR,
  input      [31:0]   dBusWishbone_DAT_MISO,
  output     [31:0]   dBusWishbone_DAT_MOSI,
  output reg [3:0]    dBusWishbone_SEL,
  input               dBusWishbone_ERR,
  output     [2:0]    dBusWishbone_CTI,
  output     [1:0]    dBusWishbone_BTE,
  input               clk,
  input               reset,
  input               debugReset
);
  wire                IBusCachedPlugin_cache_io_flush;
  wire                IBusCachedPlugin_cache_io_cpu_prefetch_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isStuck;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isRemoved;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isStuck;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isUser;
  reg                 IBusCachedPlugin_cache_io_cpu_fill_valid;
  reg        [31:0]   _zz_RegFilePlugin_regFile_port0;
  reg        [31:0]   _zz_RegFilePlugin_regFile_port1;
  wire                IBusCachedPlugin_cache_io_cpu_prefetch_haltIt;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_fetch_data;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_fetch_physicalAddress;
  wire                IBusCachedPlugin_cache_io_cpu_decode_error;
  wire                IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling;
  wire                IBusCachedPlugin_cache_io_cpu_decode_mmuException;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_decode_data;
  wire                IBusCachedPlugin_cache_io_cpu_decode_cacheMiss;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_decode_physicalAddress;
  wire                IBusCachedPlugin_cache_io_mem_cmd_valid;
  wire       [31:0]   IBusCachedPlugin_cache_io_mem_cmd_payload_address;
  wire       [2:0]    IBusCachedPlugin_cache_io_mem_cmd_payload_size;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_1;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_2;
  wire                _zz_decode_LEGAL_INSTRUCTION_3;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_4;
  wire       [12:0]   _zz_decode_LEGAL_INSTRUCTION_5;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_6;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_7;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_8;
  wire                _zz_decode_LEGAL_INSTRUCTION_9;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_10;
  wire       [6:0]    _zz_decode_LEGAL_INSTRUCTION_11;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_12;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_13;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_14;
  wire                _zz_decode_LEGAL_INSTRUCTION_15;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_16;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_17;
  wire       [1:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload_1;
  wire       [1:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload_2;
  wire       [31:0]   _zz_IBusCachedPlugin_fetchPc_pc;
  wire       [2:0]    _zz_IBusCachedPlugin_fetchPc_pc_1;
  wire       [2:0]    _zz_DBusSimplePlugin_memoryExceptionPort_payload_code;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_1;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_2;
  wire                _zz__zz_decode_ENV_CTRL_2_3;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_4;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_5;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_6;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_7;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_8;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_9;
  wire                _zz__zz_decode_ENV_CTRL_2_10;
  wire                _zz__zz_decode_ENV_CTRL_2_11;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_12;
  wire                _zz__zz_decode_ENV_CTRL_2_13;
  wire       [21:0]   _zz__zz_decode_ENV_CTRL_2_14;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_15;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_16;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_17;
  wire                _zz__zz_decode_ENV_CTRL_2_18;
  wire                _zz__zz_decode_ENV_CTRL_2_19;
  wire                _zz__zz_decode_ENV_CTRL_2_20;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_21;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_22;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_23;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_24;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_25;
  wire       [18:0]   _zz__zz_decode_ENV_CTRL_2_26;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_27;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_28;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_29;
  wire                _zz__zz_decode_ENV_CTRL_2_30;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_31;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_32;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_33;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_34;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_35;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_36;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_37;
  wire       [15:0]   _zz__zz_decode_ENV_CTRL_2_38;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_39;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_40;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_41;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_42;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_43;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_44;
  wire                _zz__zz_decode_ENV_CTRL_2_45;
  wire                _zz__zz_decode_ENV_CTRL_2_46;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_47;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_48;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_49;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_50;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_51;
  wire                _zz__zz_decode_ENV_CTRL_2_52;
  wire       [12:0]   _zz__zz_decode_ENV_CTRL_2_53;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_54;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_55;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_56;
  wire                _zz__zz_decode_ENV_CTRL_2_57;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_58;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_59;
  wire       [4:0]    _zz__zz_decode_ENV_CTRL_2_60;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_61;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_62;
  wire                _zz__zz_decode_ENV_CTRL_2_63;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_64;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_65;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_66;
  wire                _zz__zz_decode_ENV_CTRL_2_67;
  wire                _zz__zz_decode_ENV_CTRL_2_68;
  wire       [9:0]    _zz__zz_decode_ENV_CTRL_2_69;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_70;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_71;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_72;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_73;
  wire                _zz__zz_decode_ENV_CTRL_2_74;
  wire                _zz__zz_decode_ENV_CTRL_2_75;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_76;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_77;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_78;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_79;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_80;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_81;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_82;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_83;
  wire       [6:0]    _zz__zz_decode_ENV_CTRL_2_84;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_85;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_86;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_87;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_88;
  wire                _zz__zz_decode_ENV_CTRL_2_89;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_90;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_91;
  wire       [2:0]    _zz__zz_decode_ENV_CTRL_2_92;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_93;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_94;
  wire                _zz__zz_decode_ENV_CTRL_2_95;
  wire                _zz__zz_decode_ENV_CTRL_2_96;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_97;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_98;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_99;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_100;
  wire       [3:0]    _zz__zz_decode_ENV_CTRL_2_101;
  wire                _zz__zz_decode_ENV_CTRL_2_102;
  wire                _zz__zz_decode_ENV_CTRL_2_103;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_104;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_105;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_106;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_107;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_108;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_109;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_110;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_111;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_112;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_113;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_114;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_115;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_116;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_117;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_118;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_119;
  wire                _zz_RegFilePlugin_regFile_port;
  wire                _zz_decode_RegFilePlugin_rs1Data;
  wire                _zz_RegFilePlugin_regFile_port_1;
  wire                _zz_decode_RegFilePlugin_rs2Data;
  wire       [0:0]    _zz__zz_execute_REGFILE_WRITE_DATA;
  wire       [2:0]    _zz__zz_execute_SRC1;
  wire       [4:0]    _zz__zz_execute_SRC1_1;
  wire       [11:0]   _zz__zz_execute_SRC2_3;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_1;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_2;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_3;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_4;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_5;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_6;
  wire       [31:0]   _zz__zz_execute_to_memory_REGFILE_WRITE_DATA_1;
  wire       [32:0]   _zz__zz_execute_to_memory_REGFILE_WRITE_DATA_1_1;
  wire       [19:0]   _zz__zz_execute_BranchPlugin_branch_src2;
  wire       [11:0]   _zz__zz_execute_BranchPlugin_branch_src2_4;
  wire       [1:0]    _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1;
  wire       [1:0]    _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1;
  wire       [1:0]    _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3;
  wire       [1:0]    _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3_1;
  wire                _zz_when;
  wire                _zz_when_1;
  wire       [26:0]   _zz_iBusWishbone_ADR_1;
  wire       [31:0]   memory_MEMORY_READ_DATA;
  wire       [31:0]   execute_BRANCH_CALC;
  wire                execute_BRANCH_DO;
  wire       [31:0]   writeBack_REGFILE_WRITE_DATA;
  wire       [31:0]   execute_REGFILE_WRITE_DATA;
  wire       [1:0]    memory_MEMORY_ADDRESS_LOW;
  wire       [1:0]    execute_MEMORY_ADDRESS_LOW;
  wire                decode_DO_EBREAK;
  wire                decode_CSR_READ_OPCODE;
  wire                decode_CSR_WRITE_OPCODE;
  wire                decode_SRC2_FORCE_ZERO;
  wire       [31:0]   decode_RS2;
  wire       [31:0]   decode_RS1;
  wire       `EnvCtrlEnum_binary_sequential_type _zz_memory_to_writeBack_ENV_CTRL;
  wire       `EnvCtrlEnum_binary_sequential_type _zz_memory_to_writeBack_ENV_CTRL_1;
  wire       `EnvCtrlEnum_binary_sequential_type _zz_execute_to_memory_ENV_CTRL;
  wire       `EnvCtrlEnum_binary_sequential_type _zz_execute_to_memory_ENV_CTRL_1;
  wire       `EnvCtrlEnum_binary_sequential_type decode_ENV_CTRL;
  wire       `EnvCtrlEnum_binary_sequential_type _zz_decode_ENV_CTRL;
  wire       `EnvCtrlEnum_binary_sequential_type _zz_decode_to_execute_ENV_CTRL;
  wire       `EnvCtrlEnum_binary_sequential_type _zz_decode_to_execute_ENV_CTRL_1;
  wire                decode_IS_CSR;
  wire       `BranchCtrlEnum_binary_sequential_type decode_BRANCH_CTRL;
  wire       `BranchCtrlEnum_binary_sequential_type _zz_decode_BRANCH_CTRL;
  wire       `BranchCtrlEnum_binary_sequential_type _zz_decode_to_execute_BRANCH_CTRL;
  wire       `BranchCtrlEnum_binary_sequential_type _zz_decode_to_execute_BRANCH_CTRL_1;
  wire       `ShiftCtrlEnum_binary_sequential_type decode_SHIFT_CTRL;
  wire       `ShiftCtrlEnum_binary_sequential_type _zz_decode_SHIFT_CTRL;
  wire       `ShiftCtrlEnum_binary_sequential_type _zz_decode_to_execute_SHIFT_CTRL;
  wire       `ShiftCtrlEnum_binary_sequential_type _zz_decode_to_execute_SHIFT_CTRL_1;
  wire       `AluBitwiseCtrlEnum_binary_sequential_type decode_ALU_BITWISE_CTRL;
  wire       `AluBitwiseCtrlEnum_binary_sequential_type _zz_decode_ALU_BITWISE_CTRL;
  wire       `AluBitwiseCtrlEnum_binary_sequential_type _zz_decode_to_execute_ALU_BITWISE_CTRL;
  wire       `AluBitwiseCtrlEnum_binary_sequential_type _zz_decode_to_execute_ALU_BITWISE_CTRL_1;
  wire                decode_SRC_LESS_UNSIGNED;
  wire                decode_MEMORY_STORE;
  wire                execute_BYPASSABLE_MEMORY_STAGE;
  wire                decode_BYPASSABLE_MEMORY_STAGE;
  wire                decode_BYPASSABLE_EXECUTE_STAGE;
  wire       `Src2CtrlEnum_binary_sequential_type decode_SRC2_CTRL;
  wire       `Src2CtrlEnum_binary_sequential_type _zz_decode_SRC2_CTRL;
  wire       `Src2CtrlEnum_binary_sequential_type _zz_decode_to_execute_SRC2_CTRL;
  wire       `Src2CtrlEnum_binary_sequential_type _zz_decode_to_execute_SRC2_CTRL_1;
  wire       `AluCtrlEnum_binary_sequential_type decode_ALU_CTRL;
  wire       `AluCtrlEnum_binary_sequential_type _zz_decode_ALU_CTRL;
  wire       `AluCtrlEnum_binary_sequential_type _zz_decode_to_execute_ALU_CTRL;
  wire       `AluCtrlEnum_binary_sequential_type _zz_decode_to_execute_ALU_CTRL_1;
  wire                decode_MEMORY_ENABLE;
  wire       `Src1CtrlEnum_binary_sequential_type decode_SRC1_CTRL;
  wire       `Src1CtrlEnum_binary_sequential_type _zz_decode_SRC1_CTRL;
  wire       `Src1CtrlEnum_binary_sequential_type _zz_decode_to_execute_SRC1_CTRL;
  wire       `Src1CtrlEnum_binary_sequential_type _zz_decode_to_execute_SRC1_CTRL_1;
  wire       [31:0]   writeBack_FORMAL_PC_NEXT;
  wire       [31:0]   memory_FORMAL_PC_NEXT;
  wire       [31:0]   execute_FORMAL_PC_NEXT;
  wire       [31:0]   decode_FORMAL_PC_NEXT;
  wire       [31:0]   memory_PC;
  wire                execute_DO_EBREAK;
  wire                decode_IS_EBREAK;
  wire                execute_CSR_READ_OPCODE;
  wire                execute_CSR_WRITE_OPCODE;
  wire                execute_IS_CSR;
  wire       `EnvCtrlEnum_binary_sequential_type memory_ENV_CTRL;
  wire       `EnvCtrlEnum_binary_sequential_type _zz_memory_ENV_CTRL;
  wire       `EnvCtrlEnum_binary_sequential_type execute_ENV_CTRL;
  wire       `EnvCtrlEnum_binary_sequential_type _zz_execute_ENV_CTRL;
  wire       `EnvCtrlEnum_binary_sequential_type writeBack_ENV_CTRL;
  wire       `EnvCtrlEnum_binary_sequential_type _zz_writeBack_ENV_CTRL;
  wire       [31:0]   memory_BRANCH_CALC;
  wire                memory_BRANCH_DO;
  wire       [31:0]   execute_PC;
  wire       [31:0]   execute_RS1;
  wire       `BranchCtrlEnum_binary_sequential_type execute_BRANCH_CTRL;
  wire       `BranchCtrlEnum_binary_sequential_type _zz_execute_BRANCH_CTRL;
  wire                decode_RS2_USE;
  wire                decode_RS1_USE;
  wire                execute_REGFILE_WRITE_VALID;
  wire                execute_BYPASSABLE_EXECUTE_STAGE;
  wire                memory_REGFILE_WRITE_VALID;
  wire       [31:0]   memory_INSTRUCTION;
  wire                memory_BYPASSABLE_MEMORY_STAGE;
  wire                writeBack_REGFILE_WRITE_VALID;
  reg        [31:0]   _zz_execute_to_memory_REGFILE_WRITE_DATA;
  wire       `ShiftCtrlEnum_binary_sequential_type execute_SHIFT_CTRL;
  wire       `ShiftCtrlEnum_binary_sequential_type _zz_execute_SHIFT_CTRL;
  wire                execute_SRC_LESS_UNSIGNED;
  wire                execute_SRC2_FORCE_ZERO;
  wire                execute_SRC_USE_SUB_LESS;
  wire       [31:0]   _zz_execute_SRC2;
  wire       `Src2CtrlEnum_binary_sequential_type execute_SRC2_CTRL;
  wire       `Src2CtrlEnum_binary_sequential_type _zz_execute_SRC2_CTRL;
  wire       `Src1CtrlEnum_binary_sequential_type execute_SRC1_CTRL;
  wire       `Src1CtrlEnum_binary_sequential_type _zz_execute_SRC1_CTRL;
  wire                decode_SRC_USE_SUB_LESS;
  wire                decode_SRC_ADD_ZERO;
  wire       [31:0]   execute_SRC_ADD_SUB;
  wire                execute_SRC_LESS;
  wire       `AluCtrlEnum_binary_sequential_type execute_ALU_CTRL;
  wire       `AluCtrlEnum_binary_sequential_type _zz_execute_ALU_CTRL;
  wire       [31:0]   execute_SRC2;
  wire       [31:0]   execute_SRC1;
  wire       `AluBitwiseCtrlEnum_binary_sequential_type execute_ALU_BITWISE_CTRL;
  wire       `AluBitwiseCtrlEnum_binary_sequential_type _zz_execute_ALU_BITWISE_CTRL;
  wire       [31:0]   _zz_lastStageRegFileWrite_payload_address;
  wire                _zz_lastStageRegFileWrite_valid;
  reg                 _zz_1;
  wire       [31:0]   decode_INSTRUCTION_ANTICIPATED;
  reg                 decode_REGFILE_WRITE_VALID;
  wire                decode_LEGAL_INSTRUCTION;
  wire       `EnvCtrlEnum_binary_sequential_type _zz_decode_ENV_CTRL_1;
  wire       `BranchCtrlEnum_binary_sequential_type _zz_decode_BRANCH_CTRL_1;
  wire       `ShiftCtrlEnum_binary_sequential_type _zz_decode_SHIFT_CTRL_1;
  wire       `AluBitwiseCtrlEnum_binary_sequential_type _zz_decode_ALU_BITWISE_CTRL_1;
  wire       `Src2CtrlEnum_binary_sequential_type _zz_decode_SRC2_CTRL_1;
  wire       `AluCtrlEnum_binary_sequential_type _zz_decode_ALU_CTRL_1;
  wire       `Src1CtrlEnum_binary_sequential_type _zz_decode_SRC1_CTRL_1;
  wire                writeBack_MEMORY_STORE;
  reg        [31:0]   _zz_lastStageRegFileWrite_payload_data;
  wire                writeBack_MEMORY_ENABLE;
  wire       [1:0]    writeBack_MEMORY_ADDRESS_LOW;
  wire       [31:0]   writeBack_MEMORY_READ_DATA;
  wire                memory_ALIGNEMENT_FAULT;
  wire       [31:0]   memory_REGFILE_WRITE_DATA;
  wire                memory_MEMORY_STORE;
  wire                memory_MEMORY_ENABLE;
  wire       [31:0]   execute_SRC_ADD;
  wire       [31:0]   execute_RS2;
  wire       [31:0]   execute_INSTRUCTION;
  wire                execute_MEMORY_STORE;
  wire                execute_MEMORY_ENABLE;
  wire                execute_ALIGNEMENT_FAULT;
  wire                decode_FLUSH_ALL;
  reg                 IBusCachedPlugin_rsp_issueDetected_4;
  reg                 IBusCachedPlugin_rsp_issueDetected_3;
  reg                 IBusCachedPlugin_rsp_issueDetected_2;
  reg                 IBusCachedPlugin_rsp_issueDetected_1;
  wire       [31:0]   decode_INSTRUCTION;
  reg        [31:0]   _zz_memory_to_writeBack_FORMAL_PC_NEXT;
  wire       [31:0]   decode_PC;
  wire       [31:0]   writeBack_PC;
  wire       [31:0]   writeBack_INSTRUCTION;
  reg                 decode_arbitration_haltItself;
  reg                 decode_arbitration_haltByOther;
  reg                 decode_arbitration_removeIt;
  wire                decode_arbitration_flushIt;
  reg                 decode_arbitration_flushNext;
  reg                 decode_arbitration_isValid;
  wire                decode_arbitration_isStuck;
  wire                decode_arbitration_isStuckByOthers;
  wire                decode_arbitration_isFlushed;
  wire                decode_arbitration_isMoving;
  wire                decode_arbitration_isFiring;
  reg                 execute_arbitration_haltItself;
  reg                 execute_arbitration_haltByOther;
  reg                 execute_arbitration_removeIt;
  reg                 execute_arbitration_flushIt;
  reg                 execute_arbitration_flushNext;
  reg                 execute_arbitration_isValid;
  wire                execute_arbitration_isStuck;
  wire                execute_arbitration_isStuckByOthers;
  wire                execute_arbitration_isFlushed;
  wire                execute_arbitration_isMoving;
  wire                execute_arbitration_isFiring;
  reg                 memory_arbitration_haltItself;
  wire                memory_arbitration_haltByOther;
  reg                 memory_arbitration_removeIt;
  wire                memory_arbitration_flushIt;
  reg                 memory_arbitration_flushNext;
  reg                 memory_arbitration_isValid;
  wire                memory_arbitration_isStuck;
  wire                memory_arbitration_isStuckByOthers;
  wire                memory_arbitration_isFlushed;
  wire                memory_arbitration_isMoving;
  wire                memory_arbitration_isFiring;
  wire                writeBack_arbitration_haltItself;
  wire                writeBack_arbitration_haltByOther;
  reg                 writeBack_arbitration_removeIt;
  wire                writeBack_arbitration_flushIt;
  reg                 writeBack_arbitration_flushNext;
  reg                 writeBack_arbitration_isValid;
  wire                writeBack_arbitration_isStuck;
  wire                writeBack_arbitration_isStuckByOthers;
  wire                writeBack_arbitration_isFlushed;
  wire                writeBack_arbitration_isMoving;
  wire                writeBack_arbitration_isFiring;
  wire       [31:0]   lastStageInstruction /* verilator public */ ;
  wire       [31:0]   lastStagePc /* verilator public */ ;
  wire                lastStageIsValid /* verilator public */ ;
  wire                lastStageIsFiring /* verilator public */ ;
  reg                 IBusCachedPlugin_fetcherHalt;
  reg                 IBusCachedPlugin_incomingInstruction;
  wire                IBusCachedPlugin_pcValids_0;
  wire                IBusCachedPlugin_pcValids_1;
  wire                IBusCachedPlugin_pcValids_2;
  wire                IBusCachedPlugin_pcValids_3;
  reg                 IBusCachedPlugin_decodeExceptionPort_valid;
  reg        [3:0]    IBusCachedPlugin_decodeExceptionPort_payload_code;
  wire       [31:0]   IBusCachedPlugin_decodeExceptionPort_payload_badAddr;
  wire                IBusCachedPlugin_mmuBus_cmd_0_isValid;
  wire                IBusCachedPlugin_mmuBus_cmd_0_isStuck;
  wire       [31:0]   IBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  wire                IBusCachedPlugin_mmuBus_cmd_0_bypassTranslation;
  wire       [31:0]   IBusCachedPlugin_mmuBus_rsp_physicalAddress;
  wire                IBusCachedPlugin_mmuBus_rsp_isIoAccess;
  wire                IBusCachedPlugin_mmuBus_rsp_isPaging;
  wire                IBusCachedPlugin_mmuBus_rsp_allowRead;
  wire                IBusCachedPlugin_mmuBus_rsp_allowWrite;
  wire                IBusCachedPlugin_mmuBus_rsp_allowExecute;
  wire                IBusCachedPlugin_mmuBus_rsp_exception;
  wire                IBusCachedPlugin_mmuBus_rsp_refilling;
  wire                IBusCachedPlugin_mmuBus_rsp_bypassTranslation;
  wire                IBusCachedPlugin_mmuBus_end;
  wire                IBusCachedPlugin_mmuBus_busy;
  reg                 DBusSimplePlugin_memoryExceptionPort_valid;
  reg        [3:0]    DBusSimplePlugin_memoryExceptionPort_payload_code;
  wire       [31:0]   DBusSimplePlugin_memoryExceptionPort_payload_badAddr;
  wire                decodeExceptionPort_valid;
  wire       [3:0]    decodeExceptionPort_payload_code;
  wire       [31:0]   decodeExceptionPort_payload_badAddr;
  wire                BranchPlugin_jumpInterface_valid;
  wire       [31:0]   BranchPlugin_jumpInterface_payload;
  wire                BranchPlugin_branchExceptionPort_valid;
  wire       [3:0]    BranchPlugin_branchExceptionPort_payload_code;
  wire       [31:0]   BranchPlugin_branchExceptionPort_payload_badAddr;
  wire       [31:0]   CsrPlugin_csrMapping_readDataSignal;
  wire       [31:0]   CsrPlugin_csrMapping_readDataInit;
  wire       [31:0]   CsrPlugin_csrMapping_writeDataSignal;
  wire                CsrPlugin_csrMapping_allowCsrSignal;
  wire                CsrPlugin_csrMapping_hazardFree;
  wire                CsrPlugin_inWfi /* verilator public */ ;
  reg                 CsrPlugin_thirdPartyWake;
  reg                 CsrPlugin_jumpInterface_valid;
  reg        [31:0]   CsrPlugin_jumpInterface_payload;
  wire                CsrPlugin_exceptionPendings_0;
  wire                CsrPlugin_exceptionPendings_1;
  wire                CsrPlugin_exceptionPendings_2;
  wire                CsrPlugin_exceptionPendings_3;
  wire                externalInterrupt;
  wire                contextSwitching;
  reg        [1:0]    CsrPlugin_privilege;
  reg                 CsrPlugin_forceMachineWire;
  reg                 CsrPlugin_selfException_valid;
  reg        [3:0]    CsrPlugin_selfException_payload_code;
  wire       [31:0]   CsrPlugin_selfException_payload_badAddr;
  reg                 CsrPlugin_allowInterrupts;
  reg                 CsrPlugin_allowException;
  reg                 CsrPlugin_allowEbreakException;
  reg                 IBusCachedPlugin_injectionPort_valid;
  reg                 IBusCachedPlugin_injectionPort_ready;
  wire       [31:0]   IBusCachedPlugin_injectionPort_payload;
  wire                IBusCachedPlugin_externalFlush;
  wire                IBusCachedPlugin_jump_pcLoad_valid;
  wire       [31:0]   IBusCachedPlugin_jump_pcLoad_payload;
  wire       [1:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload;
  wire                IBusCachedPlugin_fetchPc_output_valid;
  wire                IBusCachedPlugin_fetchPc_output_ready;
  wire       [31:0]   IBusCachedPlugin_fetchPc_output_payload;
  reg        [31:0]   IBusCachedPlugin_fetchPc_pcReg /* verilator public */ ;
  reg                 IBusCachedPlugin_fetchPc_correction;
  reg                 IBusCachedPlugin_fetchPc_correctionReg;
  wire                IBusCachedPlugin_fetchPc_output_fire;
  wire                IBusCachedPlugin_fetchPc_corrected;
  reg                 IBusCachedPlugin_fetchPc_pcRegPropagate;
  reg                 IBusCachedPlugin_fetchPc_booted;
  reg                 IBusCachedPlugin_fetchPc_inc;
  wire                when_Fetcher_l131;
  wire                IBusCachedPlugin_fetchPc_output_fire_1;
  wire                when_Fetcher_l131_1;
  reg        [31:0]   IBusCachedPlugin_fetchPc_pc;
  wire                IBusCachedPlugin_fetchPc_redo_valid;
  wire       [31:0]   IBusCachedPlugin_fetchPc_redo_payload;
  reg                 IBusCachedPlugin_fetchPc_flushed;
  wire                when_Fetcher_l158;
  reg                 IBusCachedPlugin_iBusRsp_redoFetch;
  wire                IBusCachedPlugin_iBusRsp_stages_0_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_0_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_0_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_0_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_0_halt;
  wire                IBusCachedPlugin_iBusRsp_stages_1_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_1_halt;
  wire                IBusCachedPlugin_iBusRsp_stages_2_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_2_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_2_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_2_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_2_halt;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  wire                IBusCachedPlugin_iBusRsp_flush;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1;
  reg                 _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  reg                 _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  reg        [31:0]   _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  reg                 IBusCachedPlugin_iBusRsp_readyForError;
  wire                IBusCachedPlugin_iBusRsp_output_valid;
  wire                IBusCachedPlugin_iBusRsp_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_output_payload_pc;
  wire                IBusCachedPlugin_iBusRsp_output_payload_rsp_error;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_output_payload_rsp_inst;
  wire                IBusCachedPlugin_iBusRsp_output_payload_isRvc;
  wire                when_Fetcher_l240;
  wire                when_Fetcher_l320;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_0;
  wire                when_Fetcher_l329;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_1;
  wire                when_Fetcher_l329_1;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_2;
  wire                when_Fetcher_l329_2;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_3;
  wire                when_Fetcher_l329_3;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_4;
  wire                when_Fetcher_l329_4;
  wire                iBus_cmd_valid;
  wire                iBus_cmd_ready;
  reg        [31:0]   iBus_cmd_payload_address;
  wire       [2:0]    iBus_cmd_payload_size;
  wire                iBus_rsp_valid;
  wire       [31:0]   iBus_rsp_payload_data;
  wire                iBus_rsp_payload_error;
  wire       [31:0]   _zz_IBusCachedPlugin_rspCounter;
  reg        [31:0]   IBusCachedPlugin_rspCounter;
  wire                IBusCachedPlugin_s0_tightlyCoupledHit;
  reg                 IBusCachedPlugin_s1_tightlyCoupledHit;
  reg                 IBusCachedPlugin_s2_tightlyCoupledHit;
  wire                IBusCachedPlugin_rsp_iBusRspOutputHalt;
  wire                IBusCachedPlugin_rsp_issueDetected;
  reg                 IBusCachedPlugin_rsp_redoFetch;
  wire                when_IBusCachedPlugin_l239;
  wire                when_IBusCachedPlugin_l244;
  wire                when_IBusCachedPlugin_l250;
  wire                when_IBusCachedPlugin_l256;
  wire                when_IBusCachedPlugin_l267;
  wire                dBus_cmd_valid;
  wire                dBus_cmd_ready;
  wire                dBus_cmd_payload_wr;
  wire       [31:0]   dBus_cmd_payload_address;
  wire       [31:0]   dBus_cmd_payload_data;
  wire       [1:0]    dBus_cmd_payload_size;
  wire                dBus_rsp_ready;
  wire                dBus_rsp_error;
  wire       [31:0]   dBus_rsp_data;
  wire                _zz_dBus_cmd_valid;
  reg                 execute_DBusSimplePlugin_skipCmd;
  reg        [31:0]   _zz_dBus_cmd_payload_data;
  wire                when_DBusSimplePlugin_l426;
  reg        [3:0]    _zz_execute_DBusSimplePlugin_formalMask;
  wire       [3:0]    execute_DBusSimplePlugin_formalMask;
  wire                when_DBusSimplePlugin_l479;
  wire                when_DBusSimplePlugin_l486;
  wire                when_DBusSimplePlugin_l512;
  reg        [31:0]   writeBack_DBusSimplePlugin_rspShifted;
  wire       [1:0]    switch_Misc_l200;
  wire                _zz_writeBack_DBusSimplePlugin_rspFormated;
  reg        [31:0]   _zz_writeBack_DBusSimplePlugin_rspFormated_1;
  wire                _zz_writeBack_DBusSimplePlugin_rspFormated_2;
  reg        [31:0]   _zz_writeBack_DBusSimplePlugin_rspFormated_3;
  reg        [31:0]   writeBack_DBusSimplePlugin_rspFormated;
  wire                when_DBusSimplePlugin_l558;
  wire       [27:0]   _zz_decode_ENV_CTRL_2;
  wire                _zz_decode_ENV_CTRL_3;
  wire                _zz_decode_ENV_CTRL_4;
  wire                _zz_decode_ENV_CTRL_5;
  wire                _zz_decode_ENV_CTRL_6;
  wire       `Src1CtrlEnum_binary_sequential_type _zz_decode_SRC1_CTRL_2;
  wire       `AluCtrlEnum_binary_sequential_type _zz_decode_ALU_CTRL_2;
  wire       `Src2CtrlEnum_binary_sequential_type _zz_decode_SRC2_CTRL_2;
  wire       `AluBitwiseCtrlEnum_binary_sequential_type _zz_decode_ALU_BITWISE_CTRL_2;
  wire       `ShiftCtrlEnum_binary_sequential_type _zz_decode_SHIFT_CTRL_2;
  wire       `BranchCtrlEnum_binary_sequential_type _zz_decode_BRANCH_CTRL_2;
  wire       `EnvCtrlEnum_binary_sequential_type _zz_decode_ENV_CTRL_7;
  wire                when_RegFilePlugin_l63;
  wire       [4:0]    decode_RegFilePlugin_regFileReadAddress1;
  wire       [4:0]    decode_RegFilePlugin_regFileReadAddress2;
  wire       [31:0]   decode_RegFilePlugin_rs1Data;
  wire       [31:0]   decode_RegFilePlugin_rs2Data;
  reg                 lastStageRegFileWrite_valid /* verilator public */ ;
  reg        [4:0]    lastStageRegFileWrite_payload_address /* verilator public */ ;
  reg        [31:0]   lastStageRegFileWrite_payload_data /* verilator public */ ;
  reg                 _zz_2;
  reg        [31:0]   execute_IntAluPlugin_bitwise;
  reg        [31:0]   _zz_execute_REGFILE_WRITE_DATA;
  reg        [31:0]   _zz_execute_SRC1;
  wire                _zz_execute_SRC2_1;
  reg        [19:0]   _zz_execute_SRC2_2;
  wire                _zz_execute_SRC2_3;
  reg        [19:0]   _zz_execute_SRC2_4;
  reg        [31:0]   _zz_execute_SRC2_5;
  reg        [31:0]   execute_SrcPlugin_addSub;
  wire                execute_SrcPlugin_less;
  reg                 execute_LightShifterPlugin_isActive;
  wire                execute_LightShifterPlugin_isShift;
  reg        [4:0]    execute_LightShifterPlugin_amplitudeReg;
  wire       [4:0]    execute_LightShifterPlugin_amplitude;
  wire       [31:0]   execute_LightShifterPlugin_shiftInput;
  wire                execute_LightShifterPlugin_done;
  wire                when_ShiftPlugins_l169;
  reg        [31:0]   _zz_execute_to_memory_REGFILE_WRITE_DATA_1;
  wire                when_ShiftPlugins_l175;
  wire                when_ShiftPlugins_l184;
  reg                 HazardSimplePlugin_src0Hazard;
  reg                 HazardSimplePlugin_src1Hazard;
  wire                HazardSimplePlugin_writeBackWrites_valid;
  wire       [4:0]    HazardSimplePlugin_writeBackWrites_payload_address;
  wire       [31:0]   HazardSimplePlugin_writeBackWrites_payload_data;
  reg                 HazardSimplePlugin_writeBackBuffer_valid;
  reg        [4:0]    HazardSimplePlugin_writeBackBuffer_payload_address;
  reg        [31:0]   HazardSimplePlugin_writeBackBuffer_payload_data;
  wire                HazardSimplePlugin_addr0Match;
  wire                HazardSimplePlugin_addr1Match;
  wire                when_HazardSimplePlugin_l59;
  wire                when_HazardSimplePlugin_l62;
  wire                when_HazardSimplePlugin_l57;
  wire                when_HazardSimplePlugin_l58;
  wire                when_HazardSimplePlugin_l59_1;
  wire                when_HazardSimplePlugin_l62_1;
  wire                when_HazardSimplePlugin_l57_1;
  wire                when_HazardSimplePlugin_l58_1;
  wire                when_HazardSimplePlugin_l59_2;
  wire                when_HazardSimplePlugin_l62_2;
  wire                when_HazardSimplePlugin_l57_2;
  wire                when_HazardSimplePlugin_l58_2;
  wire                when_HazardSimplePlugin_l105;
  wire                when_HazardSimplePlugin_l108;
  wire                when_HazardSimplePlugin_l113;
  wire                execute_BranchPlugin_eq;
  wire       [2:0]    switch_Misc_l200_1;
  reg                 _zz_execute_BRANCH_DO;
  reg                 _zz_execute_BRANCH_DO_1;
  wire       [31:0]   execute_BranchPlugin_branch_src1;
  wire                _zz_execute_BranchPlugin_branch_src2;
  reg        [10:0]   _zz_execute_BranchPlugin_branch_src2_1;
  wire                _zz_execute_BranchPlugin_branch_src2_2;
  reg        [19:0]   _zz_execute_BranchPlugin_branch_src2_3;
  wire                _zz_execute_BranchPlugin_branch_src2_4;
  reg        [18:0]   _zz_execute_BranchPlugin_branch_src2_5;
  reg        [31:0]   _zz_execute_BranchPlugin_branch_src2_6;
  wire       [31:0]   execute_BranchPlugin_branch_src2;
  wire       [31:0]   execute_BranchPlugin_branchAdder;
  wire       [1:0]    CsrPlugin_misa_base;
  wire       [25:0]   CsrPlugin_misa_extensions;
  reg        [1:0]    CsrPlugin_mtvec_mode;
  reg        [29:0]   CsrPlugin_mtvec_base;
  reg        [31:0]   CsrPlugin_mepc;
  reg                 CsrPlugin_mstatus_MIE;
  reg                 CsrPlugin_mstatus_MPIE;
  reg        [1:0]    CsrPlugin_mstatus_MPP;
  reg                 CsrPlugin_mip_MEIP;
  reg                 CsrPlugin_mip_MTIP;
  reg                 CsrPlugin_mip_MSIP;
  reg                 CsrPlugin_mie_MEIE;
  reg                 CsrPlugin_mie_MTIE;
  reg                 CsrPlugin_mie_MSIE;
  reg                 CsrPlugin_mcause_interrupt;
  reg        [3:0]    CsrPlugin_mcause_exceptionCode;
  reg        [31:0]   CsrPlugin_mtval;
  reg        [63:0]   CsrPlugin_mcycle = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  reg        [63:0]   CsrPlugin_minstret = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire                _zz_when_CsrPlugin_l952;
  wire                _zz_when_CsrPlugin_l952_1;
  wire                _zz_when_CsrPlugin_l952_2;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_decode;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_execute;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_memory;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
  reg        [3:0]    CsrPlugin_exceptionPortCtrl_exceptionContext_code;
  reg        [31:0]   CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr;
  wire       [1:0]    CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped;
  wire       [1:0]    CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege;
  wire       [1:0]    _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code;
  wire                _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1;
  wire       [1:0]    _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_2;
  wire                _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3;
  wire                when_CsrPlugin_l909;
  wire                when_CsrPlugin_l909_1;
  wire                when_CsrPlugin_l909_2;
  wire                when_CsrPlugin_l909_3;
  wire                when_CsrPlugin_l922;
  reg                 CsrPlugin_interrupt_valid;
  reg        [3:0]    CsrPlugin_interrupt_code /* verilator public */ ;
  reg        [1:0]    CsrPlugin_interrupt_targetPrivilege;
  wire                when_CsrPlugin_l946;
  wire                when_CsrPlugin_l952;
  wire                when_CsrPlugin_l952_1;
  wire                when_CsrPlugin_l952_2;
  wire                CsrPlugin_exception;
  wire                CsrPlugin_lastStageWasWfi;
  reg                 CsrPlugin_pipelineLiberator_pcValids_0;
  reg                 CsrPlugin_pipelineLiberator_pcValids_1;
  reg                 CsrPlugin_pipelineLiberator_pcValids_2;
  wire                CsrPlugin_pipelineLiberator_active;
  wire                when_CsrPlugin_l980;
  wire                when_CsrPlugin_l980_1;
  wire                when_CsrPlugin_l980_2;
  wire                when_CsrPlugin_l985;
  reg                 CsrPlugin_pipelineLiberator_done;
  wire                when_CsrPlugin_l991;
  wire                CsrPlugin_interruptJump /* verilator public */ ;
  reg                 CsrPlugin_hadException /* verilator public */ ;
  reg        [1:0]    CsrPlugin_targetPrivilege;
  reg        [3:0]    CsrPlugin_trapCause;
  reg        [1:0]    CsrPlugin_xtvec_mode;
  reg        [29:0]   CsrPlugin_xtvec_base;
  wire                when_CsrPlugin_l1019;
  wire                when_CsrPlugin_l1064;
  wire       [1:0]    switch_CsrPlugin_l1068;
  reg                 execute_CsrPlugin_wfiWake;
  wire                when_CsrPlugin_l1116;
  wire                execute_CsrPlugin_blockedBySideEffects;
  reg                 execute_CsrPlugin_illegalAccess;
  reg                 execute_CsrPlugin_illegalInstruction;
  wire                when_CsrPlugin_l1136;
  wire                when_CsrPlugin_l1137;
  wire                when_CsrPlugin_l1144;
  reg                 execute_CsrPlugin_writeInstruction;
  reg                 execute_CsrPlugin_readInstruction;
  wire                execute_CsrPlugin_writeEnable;
  wire                execute_CsrPlugin_readEnable;
  wire       [31:0]   execute_CsrPlugin_readToWriteData;
  wire                switch_Misc_l200_2;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_writeDataSignal;
  wire                when_CsrPlugin_l1176;
  wire                when_CsrPlugin_l1180;
  wire       [11:0]   execute_CsrPlugin_csrAddress;
  reg        [31:0]   externalInterruptArray_regNext;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit;
  wire       [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_1;
  reg                 DebugPlugin_firstCycle;
  reg                 DebugPlugin_secondCycle;
  reg                 DebugPlugin_resetIt;
  reg                 DebugPlugin_haltIt;
  reg                 DebugPlugin_stepIt;
  reg                 DebugPlugin_isPipBusy;
  reg                 DebugPlugin_godmode;
  wire                when_DebugPlugin_l225;
  reg                 DebugPlugin_haltedByBreak;
  reg                 DebugPlugin_debugUsed /* verilator public */ ;
  reg                 DebugPlugin_disableEbreak;
  wire                DebugPlugin_allowEBreak;
  reg        [31:0]   DebugPlugin_busReadDataReg;
  reg                 _zz_when_DebugPlugin_l244;
  wire                when_DebugPlugin_l244;
  wire       [5:0]    switch_DebugPlugin_l256;
  wire                when_DebugPlugin_l260;
  wire                when_DebugPlugin_l260_1;
  wire                when_DebugPlugin_l261;
  wire                when_DebugPlugin_l261_1;
  wire                when_DebugPlugin_l262;
  wire                when_DebugPlugin_l263;
  wire                when_DebugPlugin_l264;
  wire                when_DebugPlugin_l264_1;
  wire                when_DebugPlugin_l284;
  wire                when_DebugPlugin_l287;
  wire                when_DebugPlugin_l300;
  reg                 DebugPlugin_resetIt_regNext;
  wire                when_DebugPlugin_l316;
  wire                when_Pipeline_l124;
  reg        [31:0]   decode_to_execute_PC;
  wire                when_Pipeline_l124_1;
  reg        [31:0]   execute_to_memory_PC;
  wire                when_Pipeline_l124_2;
  reg        [31:0]   memory_to_writeBack_PC;
  wire                when_Pipeline_l124_3;
  reg        [31:0]   decode_to_execute_INSTRUCTION;
  wire                when_Pipeline_l124_4;
  reg        [31:0]   execute_to_memory_INSTRUCTION;
  wire                when_Pipeline_l124_5;
  reg        [31:0]   memory_to_writeBack_INSTRUCTION;
  wire                when_Pipeline_l124_6;
  reg        [31:0]   decode_to_execute_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_7;
  reg        [31:0]   execute_to_memory_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_8;
  reg        [31:0]   memory_to_writeBack_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_9;
  reg        `Src1CtrlEnum_binary_sequential_type decode_to_execute_SRC1_CTRL;
  wire                when_Pipeline_l124_10;
  reg                 decode_to_execute_SRC_USE_SUB_LESS;
  wire                when_Pipeline_l124_11;
  reg                 decode_to_execute_MEMORY_ENABLE;
  wire                when_Pipeline_l124_12;
  reg                 execute_to_memory_MEMORY_ENABLE;
  wire                when_Pipeline_l124_13;
  reg                 memory_to_writeBack_MEMORY_ENABLE;
  wire                when_Pipeline_l124_14;
  reg        `AluCtrlEnum_binary_sequential_type decode_to_execute_ALU_CTRL;
  wire                when_Pipeline_l124_15;
  reg        `Src2CtrlEnum_binary_sequential_type decode_to_execute_SRC2_CTRL;
  wire                when_Pipeline_l124_16;
  reg                 decode_to_execute_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_17;
  reg                 execute_to_memory_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_18;
  reg                 memory_to_writeBack_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_19;
  reg                 decode_to_execute_BYPASSABLE_EXECUTE_STAGE;
  wire                when_Pipeline_l124_20;
  reg                 decode_to_execute_BYPASSABLE_MEMORY_STAGE;
  wire                when_Pipeline_l124_21;
  reg                 execute_to_memory_BYPASSABLE_MEMORY_STAGE;
  wire                when_Pipeline_l124_22;
  reg                 decode_to_execute_MEMORY_STORE;
  wire                when_Pipeline_l124_23;
  reg                 execute_to_memory_MEMORY_STORE;
  wire                when_Pipeline_l124_24;
  reg                 memory_to_writeBack_MEMORY_STORE;
  wire                when_Pipeline_l124_25;
  reg                 decode_to_execute_SRC_LESS_UNSIGNED;
  wire                when_Pipeline_l124_26;
  reg        `AluBitwiseCtrlEnum_binary_sequential_type decode_to_execute_ALU_BITWISE_CTRL;
  wire                when_Pipeline_l124_27;
  reg        `ShiftCtrlEnum_binary_sequential_type decode_to_execute_SHIFT_CTRL;
  wire                when_Pipeline_l124_28;
  reg        `BranchCtrlEnum_binary_sequential_type decode_to_execute_BRANCH_CTRL;
  wire                when_Pipeline_l124_29;
  reg                 decode_to_execute_IS_CSR;
  wire                when_Pipeline_l124_30;
  reg        `EnvCtrlEnum_binary_sequential_type decode_to_execute_ENV_CTRL;
  wire                when_Pipeline_l124_31;
  reg        `EnvCtrlEnum_binary_sequential_type execute_to_memory_ENV_CTRL;
  wire                when_Pipeline_l124_32;
  reg        `EnvCtrlEnum_binary_sequential_type memory_to_writeBack_ENV_CTRL;
  wire                when_Pipeline_l124_33;
  reg        [31:0]   decode_to_execute_RS1;
  wire                when_Pipeline_l124_34;
  reg        [31:0]   decode_to_execute_RS2;
  wire                when_Pipeline_l124_35;
  reg                 decode_to_execute_SRC2_FORCE_ZERO;
  wire                when_Pipeline_l124_36;
  reg                 decode_to_execute_CSR_WRITE_OPCODE;
  wire                when_Pipeline_l124_37;
  reg                 decode_to_execute_CSR_READ_OPCODE;
  wire                when_Pipeline_l124_38;
  reg                 decode_to_execute_DO_EBREAK;
  wire                when_Pipeline_l124_39;
  reg                 execute_to_memory_ALIGNEMENT_FAULT;
  wire                when_Pipeline_l124_40;
  reg        [1:0]    execute_to_memory_MEMORY_ADDRESS_LOW;
  wire                when_Pipeline_l124_41;
  reg        [1:0]    memory_to_writeBack_MEMORY_ADDRESS_LOW;
  wire                when_Pipeline_l124_42;
  reg        [31:0]   execute_to_memory_REGFILE_WRITE_DATA;
  wire                when_Pipeline_l124_43;
  reg        [31:0]   memory_to_writeBack_REGFILE_WRITE_DATA;
  wire                when_Pipeline_l124_44;
  reg                 execute_to_memory_BRANCH_DO;
  wire                when_Pipeline_l124_45;
  reg        [31:0]   execute_to_memory_BRANCH_CALC;
  wire                when_Pipeline_l124_46;
  reg        [31:0]   memory_to_writeBack_MEMORY_READ_DATA;
  wire                when_Pipeline_l151;
  wire                when_Pipeline_l154;
  wire                when_Pipeline_l151_1;
  wire                when_Pipeline_l154_1;
  wire                when_Pipeline_l151_2;
  wire                when_Pipeline_l154_2;
  reg        [2:0]    switch_Fetcher_l362;
  wire                when_Fetcher_l378;
  wire                when_CsrPlugin_l1264;
  reg                 execute_CsrPlugin_csr_768;
  wire                when_CsrPlugin_l1264_1;
  reg                 execute_CsrPlugin_csr_836;
  wire                when_CsrPlugin_l1264_2;
  reg                 execute_CsrPlugin_csr_772;
  wire                when_CsrPlugin_l1264_3;
  reg                 execute_CsrPlugin_csr_773;
  wire                when_CsrPlugin_l1264_4;
  reg                 execute_CsrPlugin_csr_833;
  wire                when_CsrPlugin_l1264_5;
  reg                 execute_CsrPlugin_csr_834;
  wire                when_CsrPlugin_l1264_6;
  reg                 execute_CsrPlugin_csr_835;
  wire                when_CsrPlugin_l1264_7;
  reg                 execute_CsrPlugin_csr_3008;
  wire                when_CsrPlugin_l1264_8;
  reg                 execute_CsrPlugin_csr_4032;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_2;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_3;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_4;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_5;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_6;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_7;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_8;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_9;
  wire                when_CsrPlugin_l1297;
  wire                when_CsrPlugin_l1302;
  reg        [2:0]    _zz_iBusWishbone_ADR;
  wire                when_InstructionCache_l239;
  reg                 _zz_iBus_rsp_valid;
  reg        [31:0]   iBusWishbone_DAT_MISO_regNext;
  wire                dBus_cmd_halfPipe_valid;
  wire                dBus_cmd_halfPipe_ready;
  wire                dBus_cmd_halfPipe_payload_wr;
  wire       [31:0]   dBus_cmd_halfPipe_payload_address;
  wire       [31:0]   dBus_cmd_halfPipe_payload_data;
  wire       [1:0]    dBus_cmd_halfPipe_payload_size;
  reg                 dBus_cmd_rValid;
  wire                dBus_cmd_halfPipe_fire;
  reg                 dBus_cmd_rData_wr;
  reg        [31:0]   dBus_cmd_rData_address;
  reg        [31:0]   dBus_cmd_rData_data;
  reg        [1:0]    dBus_cmd_rData_size;
  reg        [3:0]    _zz_dBusWishbone_SEL;
  wire                when_DBusSimplePlugin_l189;

  reg [39:0] _zz_memory_to_writeBack_ENV_CTRL_string;
  reg [39:0] _zz_memory_to_writeBack_ENV_CTRL_1_string;
  reg [39:0] _zz_execute_to_memory_ENV_CTRL_string;
  reg [39:0] _zz_execute_to_memory_ENV_CTRL_1_string;
  reg [39:0] decode_ENV_CTRL_string;
  reg [39:0] _zz_decode_ENV_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ENV_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ENV_CTRL_1_string;
  reg [31:0] decode_BRANCH_CTRL_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_string;
  reg [31:0] _zz_decode_to_execute_BRANCH_CTRL_string;
  reg [31:0] _zz_decode_to_execute_BRANCH_CTRL_1_string;
  reg [71:0] decode_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_to_execute_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_to_execute_SHIFT_CTRL_1_string;
  reg [39:0] decode_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string;
  reg [23:0] decode_SRC2_CTRL_string;
  reg [23:0] _zz_decode_SRC2_CTRL_string;
  reg [23:0] _zz_decode_to_execute_SRC2_CTRL_string;
  reg [23:0] _zz_decode_to_execute_SRC2_CTRL_1_string;
  reg [63:0] decode_ALU_CTRL_string;
  reg [63:0] _zz_decode_ALU_CTRL_string;
  reg [63:0] _zz_decode_to_execute_ALU_CTRL_string;
  reg [63:0] _zz_decode_to_execute_ALU_CTRL_1_string;
  reg [95:0] decode_SRC1_CTRL_string;
  reg [95:0] _zz_decode_SRC1_CTRL_string;
  reg [95:0] _zz_decode_to_execute_SRC1_CTRL_string;
  reg [95:0] _zz_decode_to_execute_SRC1_CTRL_1_string;
  reg [39:0] memory_ENV_CTRL_string;
  reg [39:0] _zz_memory_ENV_CTRL_string;
  reg [39:0] execute_ENV_CTRL_string;
  reg [39:0] _zz_execute_ENV_CTRL_string;
  reg [39:0] writeBack_ENV_CTRL_string;
  reg [39:0] _zz_writeBack_ENV_CTRL_string;
  reg [31:0] execute_BRANCH_CTRL_string;
  reg [31:0] _zz_execute_BRANCH_CTRL_string;
  reg [71:0] execute_SHIFT_CTRL_string;
  reg [71:0] _zz_execute_SHIFT_CTRL_string;
  reg [23:0] execute_SRC2_CTRL_string;
  reg [23:0] _zz_execute_SRC2_CTRL_string;
  reg [95:0] execute_SRC1_CTRL_string;
  reg [95:0] _zz_execute_SRC1_CTRL_string;
  reg [63:0] execute_ALU_CTRL_string;
  reg [63:0] _zz_execute_ALU_CTRL_string;
  reg [39:0] execute_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_execute_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_ENV_CTRL_1_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_1_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_1_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_1_string;
  reg [23:0] _zz_decode_SRC2_CTRL_1_string;
  reg [63:0] _zz_decode_ALU_CTRL_1_string;
  reg [95:0] _zz_decode_SRC1_CTRL_1_string;
  reg [95:0] _zz_decode_SRC1_CTRL_2_string;
  reg [63:0] _zz_decode_ALU_CTRL_2_string;
  reg [23:0] _zz_decode_SRC2_CTRL_2_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_2_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_2_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_2_string;
  reg [39:0] _zz_decode_ENV_CTRL_7_string;
  reg [95:0] decode_to_execute_SRC1_CTRL_string;
  reg [63:0] decode_to_execute_ALU_CTRL_string;
  reg [23:0] decode_to_execute_SRC2_CTRL_string;
  reg [39:0] decode_to_execute_ALU_BITWISE_CTRL_string;
  reg [71:0] decode_to_execute_SHIFT_CTRL_string;
  reg [31:0] decode_to_execute_BRANCH_CTRL_string;
  reg [39:0] decode_to_execute_ENV_CTRL_string;
  reg [39:0] execute_to_memory_ENV_CTRL_string;
  reg [39:0] memory_to_writeBack_ENV_CTRL_string;


  (* ram_style = "block" *) reg [31:0] RegFilePlugin_regFile [0:31] /* verilator public */ ;

  assign _zz_when = ({decodeExceptionPort_valid,IBusCachedPlugin_decodeExceptionPort_valid} != 2'b00);
  assign _zz_when_1 = ({BranchPlugin_branchExceptionPort_valid,DBusSimplePlugin_memoryExceptionPort_valid} != 2'b00);
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_1 = (_zz_IBusCachedPlugin_jump_pcLoad_payload & (~ _zz_IBusCachedPlugin_jump_pcLoad_payload_2));
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_2 = (_zz_IBusCachedPlugin_jump_pcLoad_payload - 2'b01);
  assign _zz_IBusCachedPlugin_fetchPc_pc_1 = {IBusCachedPlugin_fetchPc_inc,2'b00};
  assign _zz_IBusCachedPlugin_fetchPc_pc = {29'd0, _zz_IBusCachedPlugin_fetchPc_pc_1};
  assign _zz_DBusSimplePlugin_memoryExceptionPort_payload_code = (memory_MEMORY_STORE ? 3'b110 : 3'b100);
  assign _zz__zz_execute_REGFILE_WRITE_DATA = execute_SRC_LESS;
  assign _zz__zz_execute_SRC1 = 3'b100;
  assign _zz__zz_execute_SRC1_1 = execute_INSTRUCTION[19 : 15];
  assign _zz__zz_execute_SRC2_3 = {execute_INSTRUCTION[31 : 25],execute_INSTRUCTION[11 : 7]};
  assign _zz_execute_SrcPlugin_addSub = ($signed(_zz_execute_SrcPlugin_addSub_1) + $signed(_zz_execute_SrcPlugin_addSub_4));
  assign _zz_execute_SrcPlugin_addSub_1 = ($signed(_zz_execute_SrcPlugin_addSub_2) + $signed(_zz_execute_SrcPlugin_addSub_3));
  assign _zz_execute_SrcPlugin_addSub_2 = execute_SRC1;
  assign _zz_execute_SrcPlugin_addSub_3 = (execute_SRC_USE_SUB_LESS ? (~ execute_SRC2) : execute_SRC2);
  assign _zz_execute_SrcPlugin_addSub_4 = (execute_SRC_USE_SUB_LESS ? _zz_execute_SrcPlugin_addSub_5 : _zz_execute_SrcPlugin_addSub_6);
  assign _zz_execute_SrcPlugin_addSub_5 = 32'h00000001;
  assign _zz_execute_SrcPlugin_addSub_6 = 32'h0;
  assign _zz__zz_execute_to_memory_REGFILE_WRITE_DATA_1 = (_zz__zz_execute_to_memory_REGFILE_WRITE_DATA_1_1 >>> 1);
  assign _zz__zz_execute_to_memory_REGFILE_WRITE_DATA_1_1 = {((execute_SHIFT_CTRL == `ShiftCtrlEnum_binary_sequential_SRA_1) && execute_LightShifterPlugin_shiftInput[31]),execute_LightShifterPlugin_shiftInput};
  assign _zz__zz_execute_BranchPlugin_branch_src2 = {{{execute_INSTRUCTION[31],execute_INSTRUCTION[19 : 12]},execute_INSTRUCTION[20]},execute_INSTRUCTION[30 : 21]};
  assign _zz__zz_execute_BranchPlugin_branch_src2_4 = {{{execute_INSTRUCTION[31],execute_INSTRUCTION[7]},execute_INSTRUCTION[30 : 25]},execute_INSTRUCTION[11 : 8]};
  assign _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 = (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code & (~ _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1));
  assign _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1 = (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code - 2'b01);
  assign _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3 = (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_2 & (~ _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3_1));
  assign _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3_1 = (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_2 - 2'b01);
  assign _zz_iBusWishbone_ADR_1 = (iBus_cmd_payload_address >>> 5);
  assign _zz_decode_RegFilePlugin_rs1Data = 1'b1;
  assign _zz_decode_RegFilePlugin_rs2Data = 1'b1;
  assign _zz_decode_LEGAL_INSTRUCTION = 32'h0000107f;
  assign _zz_decode_LEGAL_INSTRUCTION_1 = (decode_INSTRUCTION & 32'h0000207f);
  assign _zz_decode_LEGAL_INSTRUCTION_2 = 32'h00002073;
  assign _zz_decode_LEGAL_INSTRUCTION_3 = ((decode_INSTRUCTION & 32'h0000407f) == 32'h00004063);
  assign _zz_decode_LEGAL_INSTRUCTION_4 = ((decode_INSTRUCTION & 32'h0000207f) == 32'h00002013);
  assign _zz_decode_LEGAL_INSTRUCTION_5 = {((decode_INSTRUCTION & 32'h0000603f) == 32'h00000023),{((decode_INSTRUCTION & 32'h0000207f) == 32'h00000003),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_6) == 32'h00000003),{(_zz_decode_LEGAL_INSTRUCTION_7 == _zz_decode_LEGAL_INSTRUCTION_8),{_zz_decode_LEGAL_INSTRUCTION_9,{_zz_decode_LEGAL_INSTRUCTION_10,_zz_decode_LEGAL_INSTRUCTION_11}}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_6 = 32'h0000505f;
  assign _zz_decode_LEGAL_INSTRUCTION_7 = (decode_INSTRUCTION & 32'h0000707b);
  assign _zz_decode_LEGAL_INSTRUCTION_8 = 32'h00000063;
  assign _zz_decode_LEGAL_INSTRUCTION_9 = ((decode_INSTRUCTION & 32'h0000607f) == 32'h0000000f);
  assign _zz_decode_LEGAL_INSTRUCTION_10 = ((decode_INSTRUCTION & 32'hfe00007f) == 32'h00000033);
  assign _zz_decode_LEGAL_INSTRUCTION_11 = {((decode_INSTRUCTION & 32'hbc00707f) == 32'h00005013),{((decode_INSTRUCTION & 32'hfc00307f) == 32'h00001013),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_12) == 32'h00005033),{(_zz_decode_LEGAL_INSTRUCTION_13 == _zz_decode_LEGAL_INSTRUCTION_14),{_zz_decode_LEGAL_INSTRUCTION_15,{_zz_decode_LEGAL_INSTRUCTION_16,_zz_decode_LEGAL_INSTRUCTION_17}}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_12 = 32'hbe00707f;
  assign _zz_decode_LEGAL_INSTRUCTION_13 = (decode_INSTRUCTION & 32'hbe00707f);
  assign _zz_decode_LEGAL_INSTRUCTION_14 = 32'h00000033;
  assign _zz_decode_LEGAL_INSTRUCTION_15 = ((decode_INSTRUCTION & 32'hdfffffff) == 32'h10200073);
  assign _zz_decode_LEGAL_INSTRUCTION_16 = ((decode_INSTRUCTION & 32'hffefffff) == 32'h00000073);
  assign _zz_decode_LEGAL_INSTRUCTION_17 = ((decode_INSTRUCTION & 32'hffffffff) == 32'h10500073);
  assign _zz__zz_decode_ENV_CTRL_2 = 32'h10103050;
  assign _zz__zz_decode_ENV_CTRL_2_1 = (decode_INSTRUCTION & 32'h10103050);
  assign _zz__zz_decode_ENV_CTRL_2_2 = 32'h00000050;
  assign _zz__zz_decode_ENV_CTRL_2_3 = ((decode_INSTRUCTION & 32'h10403050) == 32'h10000050);
  assign _zz__zz_decode_ENV_CTRL_2_4 = {(_zz__zz_decode_ENV_CTRL_2_5 == _zz__zz_decode_ENV_CTRL_2_6),(_zz__zz_decode_ENV_CTRL_2_7 == _zz__zz_decode_ENV_CTRL_2_8)};
  assign _zz__zz_decode_ENV_CTRL_2_9 = 2'b00;
  assign _zz__zz_decode_ENV_CTRL_2_10 = ({_zz_decode_ENV_CTRL_6,_zz__zz_decode_ENV_CTRL_2_11} != 2'b00);
  assign _zz__zz_decode_ENV_CTRL_2_12 = (_zz__zz_decode_ENV_CTRL_2_13 != 1'b0);
  assign _zz__zz_decode_ENV_CTRL_2_14 = {(_zz__zz_decode_ENV_CTRL_2_15 != _zz__zz_decode_ENV_CTRL_2_17),{_zz__zz_decode_ENV_CTRL_2_18,{_zz__zz_decode_ENV_CTRL_2_21,_zz__zz_decode_ENV_CTRL_2_26}}};
  assign _zz__zz_decode_ENV_CTRL_2_5 = (decode_INSTRUCTION & 32'h00001050);
  assign _zz__zz_decode_ENV_CTRL_2_6 = 32'h00001050;
  assign _zz__zz_decode_ENV_CTRL_2_7 = (decode_INSTRUCTION & 32'h00002050);
  assign _zz__zz_decode_ENV_CTRL_2_8 = 32'h00002050;
  assign _zz__zz_decode_ENV_CTRL_2_11 = ((decode_INSTRUCTION & 32'h0000001c) == 32'h00000004);
  assign _zz__zz_decode_ENV_CTRL_2_13 = ((decode_INSTRUCTION & 32'h00000058) == 32'h00000040);
  assign _zz__zz_decode_ENV_CTRL_2_15 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_16) == 32'h00005010);
  assign _zz__zz_decode_ENV_CTRL_2_17 = 1'b0;
  assign _zz__zz_decode_ENV_CTRL_2_18 = ({_zz__zz_decode_ENV_CTRL_2_19,_zz__zz_decode_ENV_CTRL_2_20} != 2'b00);
  assign _zz__zz_decode_ENV_CTRL_2_21 = ({_zz__zz_decode_ENV_CTRL_2_22,_zz__zz_decode_ENV_CTRL_2_24} != 2'b00);
  assign _zz__zz_decode_ENV_CTRL_2_26 = {(_zz__zz_decode_ENV_CTRL_2_27 != _zz__zz_decode_ENV_CTRL_2_29),{_zz__zz_decode_ENV_CTRL_2_30,{_zz__zz_decode_ENV_CTRL_2_33,_zz__zz_decode_ENV_CTRL_2_38}}};
  assign _zz__zz_decode_ENV_CTRL_2_16 = 32'h00007054;
  assign _zz__zz_decode_ENV_CTRL_2_19 = ((decode_INSTRUCTION & 32'h40003054) == 32'h40001010);
  assign _zz__zz_decode_ENV_CTRL_2_20 = ((decode_INSTRUCTION & 32'h00007054) == 32'h00001010);
  assign _zz__zz_decode_ENV_CTRL_2_22 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_23) == 32'h00000024);
  assign _zz__zz_decode_ENV_CTRL_2_24 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_25) == 32'h00001010);
  assign _zz__zz_decode_ENV_CTRL_2_27 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_28) == 32'h00001000);
  assign _zz__zz_decode_ENV_CTRL_2_29 = 1'b0;
  assign _zz__zz_decode_ENV_CTRL_2_30 = ((_zz__zz_decode_ENV_CTRL_2_31 == _zz__zz_decode_ENV_CTRL_2_32) != 1'b0);
  assign _zz__zz_decode_ENV_CTRL_2_33 = ({_zz__zz_decode_ENV_CTRL_2_34,_zz__zz_decode_ENV_CTRL_2_36} != 2'b00);
  assign _zz__zz_decode_ENV_CTRL_2_38 = {(_zz__zz_decode_ENV_CTRL_2_39 != _zz__zz_decode_ENV_CTRL_2_44),{_zz__zz_decode_ENV_CTRL_2_45,{_zz__zz_decode_ENV_CTRL_2_51,_zz__zz_decode_ENV_CTRL_2_53}}};
  assign _zz__zz_decode_ENV_CTRL_2_23 = 32'h00000064;
  assign _zz__zz_decode_ENV_CTRL_2_25 = 32'h00003054;
  assign _zz__zz_decode_ENV_CTRL_2_28 = 32'h00001000;
  assign _zz__zz_decode_ENV_CTRL_2_31 = (decode_INSTRUCTION & 32'h00003000);
  assign _zz__zz_decode_ENV_CTRL_2_32 = 32'h00002000;
  assign _zz__zz_decode_ENV_CTRL_2_34 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_35) == 32'h00002000);
  assign _zz__zz_decode_ENV_CTRL_2_36 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_37) == 32'h00001000);
  assign _zz__zz_decode_ENV_CTRL_2_39 = {(_zz__zz_decode_ENV_CTRL_2_40 == _zz__zz_decode_ENV_CTRL_2_41),(_zz__zz_decode_ENV_CTRL_2_42 == _zz__zz_decode_ENV_CTRL_2_43)};
  assign _zz__zz_decode_ENV_CTRL_2_44 = 2'b00;
  assign _zz__zz_decode_ENV_CTRL_2_45 = ({_zz__zz_decode_ENV_CTRL_2_46,{_zz__zz_decode_ENV_CTRL_2_47,_zz__zz_decode_ENV_CTRL_2_49}} != 3'b000);
  assign _zz__zz_decode_ENV_CTRL_2_51 = (_zz__zz_decode_ENV_CTRL_2_52 != 1'b0);
  assign _zz__zz_decode_ENV_CTRL_2_53 = {(_zz__zz_decode_ENV_CTRL_2_54 != _zz__zz_decode_ENV_CTRL_2_56),{_zz__zz_decode_ENV_CTRL_2_57,{_zz__zz_decode_ENV_CTRL_2_58,_zz__zz_decode_ENV_CTRL_2_69}}};
  assign _zz__zz_decode_ENV_CTRL_2_35 = 32'h00002010;
  assign _zz__zz_decode_ENV_CTRL_2_37 = 32'h00005000;
  assign _zz__zz_decode_ENV_CTRL_2_40 = (decode_INSTRUCTION & 32'h00000034);
  assign _zz__zz_decode_ENV_CTRL_2_41 = 32'h00000020;
  assign _zz__zz_decode_ENV_CTRL_2_42 = (decode_INSTRUCTION & 32'h00000064);
  assign _zz__zz_decode_ENV_CTRL_2_43 = 32'h00000020;
  assign _zz__zz_decode_ENV_CTRL_2_46 = ((decode_INSTRUCTION & 32'h00000050) == 32'h00000040);
  assign _zz__zz_decode_ENV_CTRL_2_47 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_48) == 32'h0);
  assign _zz__zz_decode_ENV_CTRL_2_49 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_50) == 32'h00000040);
  assign _zz__zz_decode_ENV_CTRL_2_52 = ((decode_INSTRUCTION & 32'h00000020) == 32'h00000020);
  assign _zz__zz_decode_ENV_CTRL_2_54 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_55) == 32'h00000010);
  assign _zz__zz_decode_ENV_CTRL_2_56 = 1'b0;
  assign _zz__zz_decode_ENV_CTRL_2_57 = (_zz_decode_ENV_CTRL_5 != 1'b0);
  assign _zz__zz_decode_ENV_CTRL_2_58 = ({_zz__zz_decode_ENV_CTRL_2_59,_zz__zz_decode_ENV_CTRL_2_60} != 6'h0);
  assign _zz__zz_decode_ENV_CTRL_2_69 = {(_zz__zz_decode_ENV_CTRL_2_70 != _zz__zz_decode_ENV_CTRL_2_73),{_zz__zz_decode_ENV_CTRL_2_74,{_zz__zz_decode_ENV_CTRL_2_77,_zz__zz_decode_ENV_CTRL_2_84}}};
  assign _zz__zz_decode_ENV_CTRL_2_48 = 32'h00000038;
  assign _zz__zz_decode_ENV_CTRL_2_50 = 32'h00103040;
  assign _zz__zz_decode_ENV_CTRL_2_55 = 32'h00000010;
  assign _zz__zz_decode_ENV_CTRL_2_59 = _zz_decode_ENV_CTRL_6;
  assign _zz__zz_decode_ENV_CTRL_2_60 = {(_zz__zz_decode_ENV_CTRL_2_61 == _zz__zz_decode_ENV_CTRL_2_62),{_zz__zz_decode_ENV_CTRL_2_63,{_zz__zz_decode_ENV_CTRL_2_65,_zz__zz_decode_ENV_CTRL_2_66}}};
  assign _zz__zz_decode_ENV_CTRL_2_70 = {_zz_decode_ENV_CTRL_4,(_zz__zz_decode_ENV_CTRL_2_71 == _zz__zz_decode_ENV_CTRL_2_72)};
  assign _zz__zz_decode_ENV_CTRL_2_73 = 2'b00;
  assign _zz__zz_decode_ENV_CTRL_2_74 = ({_zz_decode_ENV_CTRL_4,_zz__zz_decode_ENV_CTRL_2_75} != 2'b00);
  assign _zz__zz_decode_ENV_CTRL_2_77 = ({_zz__zz_decode_ENV_CTRL_2_78,_zz__zz_decode_ENV_CTRL_2_81} != 2'b00);
  assign _zz__zz_decode_ENV_CTRL_2_84 = {(_zz__zz_decode_ENV_CTRL_2_85 != _zz__zz_decode_ENV_CTRL_2_88),{_zz__zz_decode_ENV_CTRL_2_89,{_zz__zz_decode_ENV_CTRL_2_97,_zz__zz_decode_ENV_CTRL_2_101}}};
  assign _zz__zz_decode_ENV_CTRL_2_61 = (decode_INSTRUCTION & 32'h00001010);
  assign _zz__zz_decode_ENV_CTRL_2_62 = 32'h00001010;
  assign _zz__zz_decode_ENV_CTRL_2_63 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_64) == 32'h00002010);
  assign _zz__zz_decode_ENV_CTRL_2_65 = _zz_decode_ENV_CTRL_5;
  assign _zz__zz_decode_ENV_CTRL_2_66 = {_zz__zz_decode_ENV_CTRL_2_67,_zz__zz_decode_ENV_CTRL_2_68};
  assign _zz__zz_decode_ENV_CTRL_2_71 = (decode_INSTRUCTION & 32'h00000070);
  assign _zz__zz_decode_ENV_CTRL_2_72 = 32'h00000020;
  assign _zz__zz_decode_ENV_CTRL_2_75 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_76) == 32'h0);
  assign _zz__zz_decode_ENV_CTRL_2_78 = (_zz__zz_decode_ENV_CTRL_2_79 == _zz__zz_decode_ENV_CTRL_2_80);
  assign _zz__zz_decode_ENV_CTRL_2_81 = (_zz__zz_decode_ENV_CTRL_2_82 == _zz__zz_decode_ENV_CTRL_2_83);
  assign _zz__zz_decode_ENV_CTRL_2_85 = (_zz__zz_decode_ENV_CTRL_2_86 == _zz__zz_decode_ENV_CTRL_2_87);
  assign _zz__zz_decode_ENV_CTRL_2_88 = 1'b0;
  assign _zz__zz_decode_ENV_CTRL_2_89 = ({_zz__zz_decode_ENV_CTRL_2_90,_zz__zz_decode_ENV_CTRL_2_92} != 4'b0000);
  assign _zz__zz_decode_ENV_CTRL_2_97 = (_zz__zz_decode_ENV_CTRL_2_98 != _zz__zz_decode_ENV_CTRL_2_100);
  assign _zz__zz_decode_ENV_CTRL_2_101 = {_zz__zz_decode_ENV_CTRL_2_102,{_zz__zz_decode_ENV_CTRL_2_108,_zz__zz_decode_ENV_CTRL_2_112}};
  assign _zz__zz_decode_ENV_CTRL_2_64 = 32'h00002010;
  assign _zz__zz_decode_ENV_CTRL_2_67 = ((decode_INSTRUCTION & 32'h0000000c) == 32'h00000004);
  assign _zz__zz_decode_ENV_CTRL_2_68 = ((decode_INSTRUCTION & 32'h00000028) == 32'h0);
  assign _zz__zz_decode_ENV_CTRL_2_76 = 32'h00000020;
  assign _zz__zz_decode_ENV_CTRL_2_79 = (decode_INSTRUCTION & 32'h00006014);
  assign _zz__zz_decode_ENV_CTRL_2_80 = 32'h00006010;
  assign _zz__zz_decode_ENV_CTRL_2_82 = (decode_INSTRUCTION & 32'h00005014);
  assign _zz__zz_decode_ENV_CTRL_2_83 = 32'h00004010;
  assign _zz__zz_decode_ENV_CTRL_2_86 = (decode_INSTRUCTION & 32'h00006014);
  assign _zz__zz_decode_ENV_CTRL_2_87 = 32'h00002010;
  assign _zz__zz_decode_ENV_CTRL_2_90 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_91) == 32'h0);
  assign _zz__zz_decode_ENV_CTRL_2_92 = {(_zz__zz_decode_ENV_CTRL_2_93 == _zz__zz_decode_ENV_CTRL_2_94),{_zz__zz_decode_ENV_CTRL_2_95,_zz__zz_decode_ENV_CTRL_2_96}};
  assign _zz__zz_decode_ENV_CTRL_2_98 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_99) == 32'h0);
  assign _zz__zz_decode_ENV_CTRL_2_100 = 1'b0;
  assign _zz__zz_decode_ENV_CTRL_2_102 = ({_zz__zz_decode_ENV_CTRL_2_103,{_zz__zz_decode_ENV_CTRL_2_104,_zz__zz_decode_ENV_CTRL_2_106}} != 3'b000);
  assign _zz__zz_decode_ENV_CTRL_2_108 = ({_zz__zz_decode_ENV_CTRL_2_109,_zz__zz_decode_ENV_CTRL_2_111} != 2'b00);
  assign _zz__zz_decode_ENV_CTRL_2_112 = {(_zz__zz_decode_ENV_CTRL_2_113 != _zz__zz_decode_ENV_CTRL_2_116),(_zz__zz_decode_ENV_CTRL_2_117 != _zz__zz_decode_ENV_CTRL_2_119)};
  assign _zz__zz_decode_ENV_CTRL_2_91 = 32'h00000044;
  assign _zz__zz_decode_ENV_CTRL_2_93 = (decode_INSTRUCTION & 32'h00000018);
  assign _zz__zz_decode_ENV_CTRL_2_94 = 32'h0;
  assign _zz__zz_decode_ENV_CTRL_2_95 = ((decode_INSTRUCTION & 32'h00006004) == 32'h00002000);
  assign _zz__zz_decode_ENV_CTRL_2_96 = ((decode_INSTRUCTION & 32'h00005004) == 32'h00001000);
  assign _zz__zz_decode_ENV_CTRL_2_99 = 32'h00000058;
  assign _zz__zz_decode_ENV_CTRL_2_103 = ((decode_INSTRUCTION & 32'h00000044) == 32'h00000040);
  assign _zz__zz_decode_ENV_CTRL_2_104 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_105) == 32'h00002010);
  assign _zz__zz_decode_ENV_CTRL_2_106 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_107) == 32'h40000030);
  assign _zz__zz_decode_ENV_CTRL_2_109 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_110) == 32'h00000004);
  assign _zz__zz_decode_ENV_CTRL_2_111 = _zz_decode_ENV_CTRL_3;
  assign _zz__zz_decode_ENV_CTRL_2_113 = {(_zz__zz_decode_ENV_CTRL_2_114 == _zz__zz_decode_ENV_CTRL_2_115),_zz_decode_ENV_CTRL_3};
  assign _zz__zz_decode_ENV_CTRL_2_116 = 2'b00;
  assign _zz__zz_decode_ENV_CTRL_2_117 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_118) == 32'h00001008);
  assign _zz__zz_decode_ENV_CTRL_2_119 = 1'b0;
  assign _zz__zz_decode_ENV_CTRL_2_105 = 32'h00002014;
  assign _zz__zz_decode_ENV_CTRL_2_107 = 32'h40004034;
  assign _zz__zz_decode_ENV_CTRL_2_110 = 32'h00000014;
  assign _zz__zz_decode_ENV_CTRL_2_114 = (decode_INSTRUCTION & 32'h00000044);
  assign _zz__zz_decode_ENV_CTRL_2_115 = 32'h00000004;
  assign _zz__zz_decode_ENV_CTRL_2_118 = 32'h00001048;
  always @(posedge clk) begin
    if(_zz_decode_RegFilePlugin_rs1Data) begin
      _zz_RegFilePlugin_regFile_port0 <= RegFilePlugin_regFile[decode_RegFilePlugin_regFileReadAddress1];
    end
  end

  always @(posedge clk) begin
    if(_zz_decode_RegFilePlugin_rs2Data) begin
      _zz_RegFilePlugin_regFile_port1 <= RegFilePlugin_regFile[decode_RegFilePlugin_regFileReadAddress2];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      RegFilePlugin_regFile[lastStageRegFileWrite_payload_address] <= lastStageRegFileWrite_payload_data;
    end
  end

  InstructionCache IBusCachedPlugin_cache (
    .io_flush                                 (IBusCachedPlugin_cache_io_flush                       ), //i
    .io_cpu_prefetch_isValid                  (IBusCachedPlugin_cache_io_cpu_prefetch_isValid        ), //i
    .io_cpu_prefetch_haltIt                   (IBusCachedPlugin_cache_io_cpu_prefetch_haltIt         ), //o
    .io_cpu_prefetch_pc                       (IBusCachedPlugin_iBusRsp_stages_0_input_payload       ), //i
    .io_cpu_fetch_isValid                     (IBusCachedPlugin_cache_io_cpu_fetch_isValid           ), //i
    .io_cpu_fetch_isStuck                     (IBusCachedPlugin_cache_io_cpu_fetch_isStuck           ), //i
    .io_cpu_fetch_isRemoved                   (IBusCachedPlugin_cache_io_cpu_fetch_isRemoved         ), //i
    .io_cpu_fetch_pc                          (IBusCachedPlugin_iBusRsp_stages_1_input_payload       ), //i
    .io_cpu_fetch_data                        (IBusCachedPlugin_cache_io_cpu_fetch_data              ), //o
    .io_cpu_fetch_mmuRsp_physicalAddress      (IBusCachedPlugin_mmuBus_rsp_physicalAddress           ), //i
    .io_cpu_fetch_mmuRsp_isIoAccess           (IBusCachedPlugin_mmuBus_rsp_isIoAccess                ), //i
    .io_cpu_fetch_mmuRsp_isPaging             (IBusCachedPlugin_mmuBus_rsp_isPaging                  ), //i
    .io_cpu_fetch_mmuRsp_allowRead            (IBusCachedPlugin_mmuBus_rsp_allowRead                 ), //i
    .io_cpu_fetch_mmuRsp_allowWrite           (IBusCachedPlugin_mmuBus_rsp_allowWrite                ), //i
    .io_cpu_fetch_mmuRsp_allowExecute         (IBusCachedPlugin_mmuBus_rsp_allowExecute              ), //i
    .io_cpu_fetch_mmuRsp_exception            (IBusCachedPlugin_mmuBus_rsp_exception                 ), //i
    .io_cpu_fetch_mmuRsp_refilling            (IBusCachedPlugin_mmuBus_rsp_refilling                 ), //i
    .io_cpu_fetch_mmuRsp_bypassTranslation    (IBusCachedPlugin_mmuBus_rsp_bypassTranslation         ), //i
    .io_cpu_fetch_physicalAddress             (IBusCachedPlugin_cache_io_cpu_fetch_physicalAddress   ), //o
    .io_cpu_decode_isValid                    (IBusCachedPlugin_cache_io_cpu_decode_isValid          ), //i
    .io_cpu_decode_isStuck                    (IBusCachedPlugin_cache_io_cpu_decode_isStuck          ), //i
    .io_cpu_decode_pc                         (IBusCachedPlugin_iBusRsp_stages_2_input_payload       ), //i
    .io_cpu_decode_physicalAddress            (IBusCachedPlugin_cache_io_cpu_decode_physicalAddress  ), //o
    .io_cpu_decode_data                       (IBusCachedPlugin_cache_io_cpu_decode_data             ), //o
    .io_cpu_decode_cacheMiss                  (IBusCachedPlugin_cache_io_cpu_decode_cacheMiss        ), //o
    .io_cpu_decode_error                      (IBusCachedPlugin_cache_io_cpu_decode_error            ), //o
    .io_cpu_decode_mmuRefilling               (IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling     ), //o
    .io_cpu_decode_mmuException               (IBusCachedPlugin_cache_io_cpu_decode_mmuException     ), //o
    .io_cpu_decode_isUser                     (IBusCachedPlugin_cache_io_cpu_decode_isUser           ), //i
    .io_cpu_fill_valid                        (IBusCachedPlugin_cache_io_cpu_fill_valid              ), //i
    .io_cpu_fill_payload                      (IBusCachedPlugin_cache_io_cpu_decode_physicalAddress  ), //i
    .io_mem_cmd_valid                         (IBusCachedPlugin_cache_io_mem_cmd_valid               ), //o
    .io_mem_cmd_ready                         (iBus_cmd_ready                                        ), //i
    .io_mem_cmd_payload_address               (IBusCachedPlugin_cache_io_mem_cmd_payload_address     ), //o
    .io_mem_cmd_payload_size                  (IBusCachedPlugin_cache_io_mem_cmd_payload_size        ), //o
    .io_mem_rsp_valid                         (iBus_rsp_valid                                        ), //i
    .io_mem_rsp_payload_data                  (iBus_rsp_payload_data                                 ), //i
    .io_mem_rsp_payload_error                 (iBus_rsp_payload_error                                ), //i
    ._zz_when_Fetcher_l398                    (switch_Fetcher_l362                                   ), //i
    ._zz_io_cpu_fetch_data_regNextWhen        (IBusCachedPlugin_injectionPort_payload                ), //i
    .clk                                      (clk                                                   ), //i
    .reset                                    (reset                                                 )  //i
  );
  

  assign memory_MEMORY_READ_DATA = dBus_rsp_data;
  assign execute_BRANCH_CALC = {execute_BranchPlugin_branchAdder[31 : 1],1'b0};
  assign execute_BRANCH_DO = _zz_execute_BRANCH_DO_1;
  assign writeBack_REGFILE_WRITE_DATA = memory_to_writeBack_REGFILE_WRITE_DATA;
  assign execute_REGFILE_WRITE_DATA = _zz_execute_REGFILE_WRITE_DATA;
  assign memory_MEMORY_ADDRESS_LOW = execute_to_memory_MEMORY_ADDRESS_LOW;
  assign execute_MEMORY_ADDRESS_LOW = dBus_cmd_payload_address[1 : 0];
  assign decode_DO_EBREAK = (((! DebugPlugin_haltIt) && (decode_IS_EBREAK || 1'b0)) && DebugPlugin_allowEBreak);
  assign decode_CSR_READ_OPCODE = (decode_INSTRUCTION[13 : 7] != 7'h20);
  assign decode_CSR_WRITE_OPCODE = (! (((decode_INSTRUCTION[14 : 13] == 2'b01) && (decode_INSTRUCTION[19 : 15] == 5'h0)) || ((decode_INSTRUCTION[14 : 13] == 2'b11) && (decode_INSTRUCTION[19 : 15] == 5'h0))));
  assign decode_SRC2_FORCE_ZERO = (decode_SRC_ADD_ZERO && (! decode_SRC_USE_SUB_LESS));
  assign decode_RS2 = decode_RegFilePlugin_rs2Data;
  assign decode_RS1 = decode_RegFilePlugin_rs1Data;
  assign _zz_memory_to_writeBack_ENV_CTRL = _zz_memory_to_writeBack_ENV_CTRL_1;
  assign _zz_execute_to_memory_ENV_CTRL = _zz_execute_to_memory_ENV_CTRL_1;
  assign decode_ENV_CTRL = _zz_decode_ENV_CTRL;
  assign _zz_decode_to_execute_ENV_CTRL = _zz_decode_to_execute_ENV_CTRL_1;
  assign decode_IS_CSR = _zz_decode_ENV_CTRL_2[24];
  assign decode_BRANCH_CTRL = _zz_decode_BRANCH_CTRL;
  assign _zz_decode_to_execute_BRANCH_CTRL = _zz_decode_to_execute_BRANCH_CTRL_1;
  assign decode_SHIFT_CTRL = _zz_decode_SHIFT_CTRL;
  assign _zz_decode_to_execute_SHIFT_CTRL = _zz_decode_to_execute_SHIFT_CTRL_1;
  assign decode_ALU_BITWISE_CTRL = _zz_decode_ALU_BITWISE_CTRL;
  assign _zz_decode_to_execute_ALU_BITWISE_CTRL = _zz_decode_to_execute_ALU_BITWISE_CTRL_1;
  assign decode_SRC_LESS_UNSIGNED = _zz_decode_ENV_CTRL_2[16];
  assign decode_MEMORY_STORE = _zz_decode_ENV_CTRL_2[13];
  assign execute_BYPASSABLE_MEMORY_STAGE = decode_to_execute_BYPASSABLE_MEMORY_STAGE;
  assign decode_BYPASSABLE_MEMORY_STAGE = _zz_decode_ENV_CTRL_2[12];
  assign decode_BYPASSABLE_EXECUTE_STAGE = _zz_decode_ENV_CTRL_2[11];
  assign decode_SRC2_CTRL = _zz_decode_SRC2_CTRL;
  assign _zz_decode_to_execute_SRC2_CTRL = _zz_decode_to_execute_SRC2_CTRL_1;
  assign decode_ALU_CTRL = _zz_decode_ALU_CTRL;
  assign _zz_decode_to_execute_ALU_CTRL = _zz_decode_to_execute_ALU_CTRL_1;
  assign decode_MEMORY_ENABLE = _zz_decode_ENV_CTRL_2[4];
  assign decode_SRC1_CTRL = _zz_decode_SRC1_CTRL;
  assign _zz_decode_to_execute_SRC1_CTRL = _zz_decode_to_execute_SRC1_CTRL_1;
  assign writeBack_FORMAL_PC_NEXT = memory_to_writeBack_FORMAL_PC_NEXT;
  assign memory_FORMAL_PC_NEXT = execute_to_memory_FORMAL_PC_NEXT;
  assign execute_FORMAL_PC_NEXT = decode_to_execute_FORMAL_PC_NEXT;
  assign decode_FORMAL_PC_NEXT = (decode_PC + 32'h00000004);
  assign memory_PC = execute_to_memory_PC;
  assign execute_DO_EBREAK = decode_to_execute_DO_EBREAK;
  assign decode_IS_EBREAK = _zz_decode_ENV_CTRL_2[27];
  assign execute_CSR_READ_OPCODE = decode_to_execute_CSR_READ_OPCODE;
  assign execute_CSR_WRITE_OPCODE = decode_to_execute_CSR_WRITE_OPCODE;
  assign execute_IS_CSR = decode_to_execute_IS_CSR;
  assign memory_ENV_CTRL = _zz_memory_ENV_CTRL;
  assign execute_ENV_CTRL = _zz_execute_ENV_CTRL;
  assign writeBack_ENV_CTRL = _zz_writeBack_ENV_CTRL;
  assign memory_BRANCH_CALC = execute_to_memory_BRANCH_CALC;
  assign memory_BRANCH_DO = execute_to_memory_BRANCH_DO;
  assign execute_PC = decode_to_execute_PC;
  assign execute_RS1 = decode_to_execute_RS1;
  assign execute_BRANCH_CTRL = _zz_execute_BRANCH_CTRL;
  assign decode_RS2_USE = _zz_decode_ENV_CTRL_2[15];
  assign decode_RS1_USE = _zz_decode_ENV_CTRL_2[5];
  assign execute_REGFILE_WRITE_VALID = decode_to_execute_REGFILE_WRITE_VALID;
  assign execute_BYPASSABLE_EXECUTE_STAGE = decode_to_execute_BYPASSABLE_EXECUTE_STAGE;
  assign memory_REGFILE_WRITE_VALID = execute_to_memory_REGFILE_WRITE_VALID;
  assign memory_INSTRUCTION = execute_to_memory_INSTRUCTION;
  assign memory_BYPASSABLE_MEMORY_STAGE = execute_to_memory_BYPASSABLE_MEMORY_STAGE;
  assign writeBack_REGFILE_WRITE_VALID = memory_to_writeBack_REGFILE_WRITE_VALID;
  always @(*) begin
    _zz_execute_to_memory_REGFILE_WRITE_DATA = execute_REGFILE_WRITE_DATA;
    if(when_ShiftPlugins_l169) begin
      _zz_execute_to_memory_REGFILE_WRITE_DATA = _zz_execute_to_memory_REGFILE_WRITE_DATA_1;
    end
    if(when_CsrPlugin_l1176) begin
      _zz_execute_to_memory_REGFILE_WRITE_DATA = CsrPlugin_csrMapping_readDataSignal;
    end
  end

  assign execute_SHIFT_CTRL = _zz_execute_SHIFT_CTRL;
  assign execute_SRC_LESS_UNSIGNED = decode_to_execute_SRC_LESS_UNSIGNED;
  assign execute_SRC2_FORCE_ZERO = decode_to_execute_SRC2_FORCE_ZERO;
  assign execute_SRC_USE_SUB_LESS = decode_to_execute_SRC_USE_SUB_LESS;
  assign _zz_execute_SRC2 = execute_PC;
  assign execute_SRC2_CTRL = _zz_execute_SRC2_CTRL;
  assign execute_SRC1_CTRL = _zz_execute_SRC1_CTRL;
  assign decode_SRC_USE_SUB_LESS = _zz_decode_ENV_CTRL_2[3];
  assign decode_SRC_ADD_ZERO = _zz_decode_ENV_CTRL_2[19];
  assign execute_SRC_ADD_SUB = execute_SrcPlugin_addSub;
  assign execute_SRC_LESS = execute_SrcPlugin_less;
  assign execute_ALU_CTRL = _zz_execute_ALU_CTRL;
  assign execute_SRC2 = _zz_execute_SRC2_5;
  assign execute_SRC1 = _zz_execute_SRC1;
  assign execute_ALU_BITWISE_CTRL = _zz_execute_ALU_BITWISE_CTRL;
  assign _zz_lastStageRegFileWrite_payload_address = writeBack_INSTRUCTION;
  assign _zz_lastStageRegFileWrite_valid = writeBack_REGFILE_WRITE_VALID;
  always @(*) begin
    _zz_1 = 1'b0;
    if(lastStageRegFileWrite_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign decode_INSTRUCTION_ANTICIPATED = (decode_arbitration_isStuck ? decode_INSTRUCTION : IBusCachedPlugin_cache_io_cpu_fetch_data);
  always @(*) begin
    decode_REGFILE_WRITE_VALID = _zz_decode_ENV_CTRL_2[10];
    if(when_RegFilePlugin_l63) begin
      decode_REGFILE_WRITE_VALID = 1'b0;
    end
  end

  assign decode_LEGAL_INSTRUCTION = ({((decode_INSTRUCTION & 32'h0000005f) == 32'h00000017),{((decode_INSTRUCTION & 32'h0000007f) == 32'h0000006f),{((decode_INSTRUCTION & 32'h0000106f) == 32'h00000003),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION) == 32'h00001073),{(_zz_decode_LEGAL_INSTRUCTION_1 == _zz_decode_LEGAL_INSTRUCTION_2),{_zz_decode_LEGAL_INSTRUCTION_3,{_zz_decode_LEGAL_INSTRUCTION_4,_zz_decode_LEGAL_INSTRUCTION_5}}}}}}} != 20'h0);
  assign writeBack_MEMORY_STORE = memory_to_writeBack_MEMORY_STORE;
  always @(*) begin
    _zz_lastStageRegFileWrite_payload_data = writeBack_REGFILE_WRITE_DATA;
    if(when_DBusSimplePlugin_l558) begin
      _zz_lastStageRegFileWrite_payload_data = writeBack_DBusSimplePlugin_rspFormated;
    end
  end

  assign writeBack_MEMORY_ENABLE = memory_to_writeBack_MEMORY_ENABLE;
  assign writeBack_MEMORY_ADDRESS_LOW = memory_to_writeBack_MEMORY_ADDRESS_LOW;
  assign writeBack_MEMORY_READ_DATA = memory_to_writeBack_MEMORY_READ_DATA;
  assign memory_ALIGNEMENT_FAULT = execute_to_memory_ALIGNEMENT_FAULT;
  assign memory_REGFILE_WRITE_DATA = execute_to_memory_REGFILE_WRITE_DATA;
  assign memory_MEMORY_STORE = execute_to_memory_MEMORY_STORE;
  assign memory_MEMORY_ENABLE = execute_to_memory_MEMORY_ENABLE;
  assign execute_SRC_ADD = execute_SrcPlugin_addSub;
  assign execute_RS2 = decode_to_execute_RS2;
  assign execute_INSTRUCTION = decode_to_execute_INSTRUCTION;
  assign execute_MEMORY_STORE = decode_to_execute_MEMORY_STORE;
  assign execute_MEMORY_ENABLE = decode_to_execute_MEMORY_ENABLE;
  assign execute_ALIGNEMENT_FAULT = (((dBus_cmd_payload_size == 2'b10) && (dBus_cmd_payload_address[1 : 0] != 2'b00)) || ((dBus_cmd_payload_size == 2'b01) && (dBus_cmd_payload_address[0 : 0] != 1'b0)));
  assign decode_FLUSH_ALL = _zz_decode_ENV_CTRL_2[0];
  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_4 = IBusCachedPlugin_rsp_issueDetected_3;
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_rsp_issueDetected_4 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_3 = IBusCachedPlugin_rsp_issueDetected_2;
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_rsp_issueDetected_3 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_2 = IBusCachedPlugin_rsp_issueDetected_1;
    if(when_IBusCachedPlugin_l244) begin
      IBusCachedPlugin_rsp_issueDetected_2 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_1 = IBusCachedPlugin_rsp_issueDetected;
    if(when_IBusCachedPlugin_l239) begin
      IBusCachedPlugin_rsp_issueDetected_1 = 1'b1;
    end
  end

  assign decode_INSTRUCTION = IBusCachedPlugin_iBusRsp_output_payload_rsp_inst;
  always @(*) begin
    _zz_memory_to_writeBack_FORMAL_PC_NEXT = memory_FORMAL_PC_NEXT;
    if(BranchPlugin_jumpInterface_valid) begin
      _zz_memory_to_writeBack_FORMAL_PC_NEXT = BranchPlugin_jumpInterface_payload;
    end
  end

  assign decode_PC = IBusCachedPlugin_iBusRsp_output_payload_pc;
  assign writeBack_PC = memory_to_writeBack_PC;
  assign writeBack_INSTRUCTION = memory_to_writeBack_INSTRUCTION;
  always @(*) begin
    decode_arbitration_haltItself = 1'b0;
    case(switch_Fetcher_l362)
      3'b010 : begin
        decode_arbitration_haltItself = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    decode_arbitration_haltByOther = 1'b0;
    if(when_HazardSimplePlugin_l113) begin
      decode_arbitration_haltByOther = 1'b1;
    end
    if(CsrPlugin_pipelineLiberator_active) begin
      decode_arbitration_haltByOther = 1'b1;
    end
    if(when_CsrPlugin_l1116) begin
      decode_arbitration_haltByOther = 1'b1;
    end
  end

  always @(*) begin
    decode_arbitration_removeIt = 1'b0;
    if(_zz_when) begin
      decode_arbitration_removeIt = 1'b1;
    end
    if(decode_arbitration_isFlushed) begin
      decode_arbitration_removeIt = 1'b1;
    end
  end

  assign decode_arbitration_flushIt = 1'b0;
  always @(*) begin
    decode_arbitration_flushNext = 1'b0;
    if(_zz_when) begin
      decode_arbitration_flushNext = 1'b1;
    end
  end

  always @(*) begin
    execute_arbitration_haltItself = 1'b0;
    if(when_DBusSimplePlugin_l426) begin
      execute_arbitration_haltItself = 1'b1;
    end
    if(when_ShiftPlugins_l169) begin
      if(when_ShiftPlugins_l184) begin
        execute_arbitration_haltItself = 1'b1;
      end
    end
    if(when_CsrPlugin_l1180) begin
      if(execute_CsrPlugin_blockedBySideEffects) begin
        execute_arbitration_haltItself = 1'b1;
      end
    end
  end

  always @(*) begin
    execute_arbitration_haltByOther = 1'b0;
    if(when_DebugPlugin_l284) begin
      execute_arbitration_haltByOther = 1'b1;
    end
  end

  always @(*) begin
    execute_arbitration_removeIt = 1'b0;
    if(CsrPlugin_selfException_valid) begin
      execute_arbitration_removeIt = 1'b1;
    end
    if(execute_arbitration_isFlushed) begin
      execute_arbitration_removeIt = 1'b1;
    end
  end

  always @(*) begin
    execute_arbitration_flushIt = 1'b0;
    if(when_DebugPlugin_l284) begin
      if(when_DebugPlugin_l287) begin
        execute_arbitration_flushIt = 1'b1;
      end
    end
  end

  always @(*) begin
    execute_arbitration_flushNext = 1'b0;
    if(CsrPlugin_selfException_valid) begin
      execute_arbitration_flushNext = 1'b1;
    end
    if(when_DebugPlugin_l284) begin
      if(when_DebugPlugin_l287) begin
        execute_arbitration_flushNext = 1'b1;
      end
    end
  end

  always @(*) begin
    memory_arbitration_haltItself = 1'b0;
    if(when_DBusSimplePlugin_l479) begin
      memory_arbitration_haltItself = 1'b1;
    end
  end

  assign memory_arbitration_haltByOther = 1'b0;
  always @(*) begin
    memory_arbitration_removeIt = 1'b0;
    if(_zz_when_1) begin
      memory_arbitration_removeIt = 1'b1;
    end
    if(memory_arbitration_isFlushed) begin
      memory_arbitration_removeIt = 1'b1;
    end
  end

  assign memory_arbitration_flushIt = 1'b0;
  always @(*) begin
    memory_arbitration_flushNext = 1'b0;
    if(BranchPlugin_jumpInterface_valid) begin
      memory_arbitration_flushNext = 1'b1;
    end
    if(_zz_when_1) begin
      memory_arbitration_flushNext = 1'b1;
    end
  end

  assign writeBack_arbitration_haltItself = 1'b0;
  assign writeBack_arbitration_haltByOther = 1'b0;
  always @(*) begin
    writeBack_arbitration_removeIt = 1'b0;
    if(writeBack_arbitration_isFlushed) begin
      writeBack_arbitration_removeIt = 1'b1;
    end
  end

  assign writeBack_arbitration_flushIt = 1'b0;
  always @(*) begin
    writeBack_arbitration_flushNext = 1'b0;
    if(when_CsrPlugin_l1019) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
    if(when_CsrPlugin_l1064) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
  end

  assign lastStageInstruction = writeBack_INSTRUCTION;
  assign lastStagePc = writeBack_PC;
  assign lastStageIsValid = writeBack_arbitration_isValid;
  assign lastStageIsFiring = writeBack_arbitration_isFiring;
  always @(*) begin
    IBusCachedPlugin_fetcherHalt = 1'b0;
    if(when_CsrPlugin_l922) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_CsrPlugin_l1019) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_CsrPlugin_l1064) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_DebugPlugin_l284) begin
      if(when_DebugPlugin_l287) begin
        IBusCachedPlugin_fetcherHalt = 1'b1;
      end
    end
    if(DebugPlugin_haltIt) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_DebugPlugin_l300) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_incomingInstruction = 1'b0;
    if(when_Fetcher_l240) begin
      IBusCachedPlugin_incomingInstruction = 1'b1;
    end
  end

  assign CsrPlugin_csrMapping_allowCsrSignal = 1'b0;
  assign CsrPlugin_csrMapping_readDataSignal = CsrPlugin_csrMapping_readDataInit;
  assign CsrPlugin_inWfi = 1'b0;
  always @(*) begin
    CsrPlugin_thirdPartyWake = 1'b0;
    if(DebugPlugin_haltIt) begin
      CsrPlugin_thirdPartyWake = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_jumpInterface_valid = 1'b0;
    if(when_CsrPlugin_l1019) begin
      CsrPlugin_jumpInterface_valid = 1'b1;
    end
    if(when_CsrPlugin_l1064) begin
      CsrPlugin_jumpInterface_valid = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_jumpInterface_payload = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_CsrPlugin_l1019) begin
      CsrPlugin_jumpInterface_payload = {CsrPlugin_xtvec_base,2'b00};
    end
    if(when_CsrPlugin_l1064) begin
      case(switch_CsrPlugin_l1068)
        2'b11 : begin
          CsrPlugin_jumpInterface_payload = CsrPlugin_mepc;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    CsrPlugin_forceMachineWire = 1'b0;
    if(DebugPlugin_godmode) begin
      CsrPlugin_forceMachineWire = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_allowInterrupts = 1'b1;
    if(when_DebugPlugin_l316) begin
      CsrPlugin_allowInterrupts = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_allowException = 1'b1;
    if(DebugPlugin_godmode) begin
      CsrPlugin_allowException = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_allowEbreakException = 1'b1;
    if(DebugPlugin_allowEBreak) begin
      CsrPlugin_allowEbreakException = 1'b0;
    end
  end

  assign IBusCachedPlugin_externalFlush = ({writeBack_arbitration_flushNext,{memory_arbitration_flushNext,{execute_arbitration_flushNext,decode_arbitration_flushNext}}} != 4'b0000);
  assign IBusCachedPlugin_jump_pcLoad_valid = ({CsrPlugin_jumpInterface_valid,BranchPlugin_jumpInterface_valid} != 2'b00);
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload = {BranchPlugin_jumpInterface_valid,CsrPlugin_jumpInterface_valid};
  assign IBusCachedPlugin_jump_pcLoad_payload = (_zz_IBusCachedPlugin_jump_pcLoad_payload_1[0] ? CsrPlugin_jumpInterface_payload : BranchPlugin_jumpInterface_payload);
  always @(*) begin
    IBusCachedPlugin_fetchPc_correction = 1'b0;
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_correction = 1'b1;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_correction = 1'b1;
    end
  end

  assign IBusCachedPlugin_fetchPc_output_fire = (IBusCachedPlugin_fetchPc_output_valid && IBusCachedPlugin_fetchPc_output_ready);
  assign IBusCachedPlugin_fetchPc_corrected = (IBusCachedPlugin_fetchPc_correction || IBusCachedPlugin_fetchPc_correctionReg);
  always @(*) begin
    IBusCachedPlugin_fetchPc_pcRegPropagate = 1'b0;
    if(IBusCachedPlugin_iBusRsp_stages_1_input_ready) begin
      IBusCachedPlugin_fetchPc_pcRegPropagate = 1'b1;
    end
  end

  assign when_Fetcher_l131 = (IBusCachedPlugin_fetchPc_correction || IBusCachedPlugin_fetchPc_pcRegPropagate);
  assign IBusCachedPlugin_fetchPc_output_fire_1 = (IBusCachedPlugin_fetchPc_output_valid && IBusCachedPlugin_fetchPc_output_ready);
  assign when_Fetcher_l131_1 = ((! IBusCachedPlugin_fetchPc_output_valid) && IBusCachedPlugin_fetchPc_output_ready);
  always @(*) begin
    IBusCachedPlugin_fetchPc_pc = (IBusCachedPlugin_fetchPc_pcReg + _zz_IBusCachedPlugin_fetchPc_pc);
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_pc = IBusCachedPlugin_fetchPc_redo_payload;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_pc = IBusCachedPlugin_jump_pcLoad_payload;
    end
    IBusCachedPlugin_fetchPc_pc[0] = 1'b0;
    IBusCachedPlugin_fetchPc_pc[1] = 1'b0;
  end

  always @(*) begin
    IBusCachedPlugin_fetchPc_flushed = 1'b0;
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_flushed = 1'b1;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_flushed = 1'b1;
    end
  end

  assign when_Fetcher_l158 = (IBusCachedPlugin_fetchPc_booted && ((IBusCachedPlugin_fetchPc_output_ready || IBusCachedPlugin_fetchPc_correction) || IBusCachedPlugin_fetchPc_pcRegPropagate));
  assign IBusCachedPlugin_fetchPc_output_valid = ((! IBusCachedPlugin_fetcherHalt) && IBusCachedPlugin_fetchPc_booted);
  assign IBusCachedPlugin_fetchPc_output_payload = IBusCachedPlugin_fetchPc_pc;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_redoFetch = 1'b0;
    if(IBusCachedPlugin_rsp_redoFetch) begin
      IBusCachedPlugin_iBusRsp_redoFetch = 1'b1;
    end
  end

  assign IBusCachedPlugin_iBusRsp_stages_0_input_valid = IBusCachedPlugin_fetchPc_output_valid;
  assign IBusCachedPlugin_fetchPc_output_ready = IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  assign IBusCachedPlugin_iBusRsp_stages_0_input_payload = IBusCachedPlugin_fetchPc_output_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_0_halt = 1'b0;
    if(IBusCachedPlugin_cache_io_cpu_prefetch_haltIt) begin
      IBusCachedPlugin_iBusRsp_stages_0_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready = (! IBusCachedPlugin_iBusRsp_stages_0_halt);
  assign IBusCachedPlugin_iBusRsp_stages_0_input_ready = (IBusCachedPlugin_iBusRsp_stages_0_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_valid = (IBusCachedPlugin_iBusRsp_stages_0_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_payload = IBusCachedPlugin_iBusRsp_stages_0_input_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_1_halt = 1'b0;
    if(IBusCachedPlugin_mmuBus_busy) begin
      IBusCachedPlugin_iBusRsp_stages_1_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready = (! IBusCachedPlugin_iBusRsp_stages_1_halt);
  assign IBusCachedPlugin_iBusRsp_stages_1_input_ready = (IBusCachedPlugin_iBusRsp_stages_1_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_valid = (IBusCachedPlugin_iBusRsp_stages_1_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_payload = IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_2_halt = 1'b0;
    if(when_IBusCachedPlugin_l267) begin
      IBusCachedPlugin_iBusRsp_stages_2_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready = (! IBusCachedPlugin_iBusRsp_stages_2_halt);
  assign IBusCachedPlugin_iBusRsp_stages_2_input_ready = (IBusCachedPlugin_iBusRsp_stages_2_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_2_output_valid = (IBusCachedPlugin_iBusRsp_stages_2_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_2_output_payload = IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  assign IBusCachedPlugin_fetchPc_redo_valid = IBusCachedPlugin_iBusRsp_redoFetch;
  assign IBusCachedPlugin_fetchPc_redo_payload = IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  assign IBusCachedPlugin_iBusRsp_flush = ((decode_arbitration_removeIt || (decode_arbitration_flushNext && (! decode_arbitration_isStuck))) || IBusCachedPlugin_iBusRsp_redoFetch);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_ready = _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  assign _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready = ((1'b0 && (! _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1)) || IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1 = _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2;
  assign IBusCachedPlugin_iBusRsp_stages_1_input_valid = _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1;
  assign IBusCachedPlugin_iBusRsp_stages_1_input_payload = IBusCachedPlugin_fetchPc_pcReg;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_ready = ((1'b0 && (! IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid)) || IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid = _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload = _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  assign IBusCachedPlugin_iBusRsp_stages_2_input_valid = IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready = IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  assign IBusCachedPlugin_iBusRsp_stages_2_input_payload = IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_readyForError = 1'b1;
    if(when_Fetcher_l320) begin
      IBusCachedPlugin_iBusRsp_readyForError = 1'b0;
    end
  end

  assign when_Fetcher_l240 = (IBusCachedPlugin_iBusRsp_stages_1_input_valid || IBusCachedPlugin_iBusRsp_stages_2_input_valid);
  assign when_Fetcher_l320 = (! IBusCachedPlugin_pcValids_0);
  assign when_Fetcher_l329 = (! (! IBusCachedPlugin_iBusRsp_stages_1_input_ready));
  assign when_Fetcher_l329_1 = (! (! IBusCachedPlugin_iBusRsp_stages_2_input_ready));
  assign when_Fetcher_l329_2 = (! execute_arbitration_isStuck);
  assign when_Fetcher_l329_3 = (! memory_arbitration_isStuck);
  assign when_Fetcher_l329_4 = (! writeBack_arbitration_isStuck);
  assign IBusCachedPlugin_pcValids_0 = IBusCachedPlugin_injector_nextPcCalc_valids_1;
  assign IBusCachedPlugin_pcValids_1 = IBusCachedPlugin_injector_nextPcCalc_valids_2;
  assign IBusCachedPlugin_pcValids_2 = IBusCachedPlugin_injector_nextPcCalc_valids_3;
  assign IBusCachedPlugin_pcValids_3 = IBusCachedPlugin_injector_nextPcCalc_valids_4;
  assign IBusCachedPlugin_iBusRsp_output_ready = (! decode_arbitration_isStuck);
  always @(*) begin
    decode_arbitration_isValid = IBusCachedPlugin_iBusRsp_output_valid;
    case(switch_Fetcher_l362)
      3'b010 : begin
        decode_arbitration_isValid = 1'b1;
      end
      3'b011 : begin
        decode_arbitration_isValid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign iBus_cmd_valid = IBusCachedPlugin_cache_io_mem_cmd_valid;
  always @(*) begin
    iBus_cmd_payload_address = IBusCachedPlugin_cache_io_mem_cmd_payload_address;
    iBus_cmd_payload_address = IBusCachedPlugin_cache_io_mem_cmd_payload_address;
  end

  assign iBus_cmd_payload_size = IBusCachedPlugin_cache_io_mem_cmd_payload_size;
  assign IBusCachedPlugin_s0_tightlyCoupledHit = 1'b0;
  assign IBusCachedPlugin_cache_io_cpu_prefetch_isValid = (IBusCachedPlugin_iBusRsp_stages_0_input_valid && (! IBusCachedPlugin_s0_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_fetch_isValid = (IBusCachedPlugin_iBusRsp_stages_1_input_valid && (! IBusCachedPlugin_s1_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_fetch_isStuck = (! IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_mmuBus_cmd_0_isValid = IBusCachedPlugin_cache_io_cpu_fetch_isValid;
  assign IBusCachedPlugin_mmuBus_cmd_0_isStuck = (! IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_mmuBus_cmd_0_virtualAddress = IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  assign IBusCachedPlugin_mmuBus_cmd_0_bypassTranslation = 1'b0;
  assign IBusCachedPlugin_mmuBus_end = (IBusCachedPlugin_iBusRsp_stages_1_input_ready || IBusCachedPlugin_externalFlush);
  assign IBusCachedPlugin_cache_io_cpu_decode_isValid = (IBusCachedPlugin_iBusRsp_stages_2_input_valid && (! IBusCachedPlugin_s2_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_decode_isStuck = (! IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_cache_io_cpu_decode_isUser = (CsrPlugin_privilege == 2'b00);
  assign IBusCachedPlugin_rsp_iBusRspOutputHalt = 1'b0;
  assign IBusCachedPlugin_rsp_issueDetected = 1'b0;
  always @(*) begin
    IBusCachedPlugin_rsp_redoFetch = 1'b0;
    if(when_IBusCachedPlugin_l239) begin
      IBusCachedPlugin_rsp_redoFetch = 1'b1;
    end
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_rsp_redoFetch = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_cache_io_cpu_fill_valid = (IBusCachedPlugin_rsp_redoFetch && (! IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling));
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_cache_io_cpu_fill_valid = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_decodeExceptionPort_valid = 1'b0;
    if(when_IBusCachedPlugin_l244) begin
      IBusCachedPlugin_decodeExceptionPort_valid = IBusCachedPlugin_iBusRsp_readyForError;
    end
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_decodeExceptionPort_valid = IBusCachedPlugin_iBusRsp_readyForError;
    end
  end

  always @(*) begin
    IBusCachedPlugin_decodeExceptionPort_payload_code = 4'bxxxx;
    if(when_IBusCachedPlugin_l244) begin
      IBusCachedPlugin_decodeExceptionPort_payload_code = 4'b1100;
    end
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_decodeExceptionPort_payload_code = 4'b0001;
    end
  end

  assign IBusCachedPlugin_decodeExceptionPort_payload_badAddr = {IBusCachedPlugin_iBusRsp_stages_2_input_payload[31 : 2],2'b00};
  assign when_IBusCachedPlugin_l239 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling) && (! IBusCachedPlugin_rsp_issueDetected));
  assign when_IBusCachedPlugin_l244 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_mmuException) && (! IBusCachedPlugin_rsp_issueDetected_1));
  assign when_IBusCachedPlugin_l250 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_cacheMiss) && (! IBusCachedPlugin_rsp_issueDetected_2));
  assign when_IBusCachedPlugin_l256 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_error) && (! IBusCachedPlugin_rsp_issueDetected_3));
  assign when_IBusCachedPlugin_l267 = (IBusCachedPlugin_rsp_issueDetected_4 || IBusCachedPlugin_rsp_iBusRspOutputHalt);
  assign IBusCachedPlugin_iBusRsp_output_valid = IBusCachedPlugin_iBusRsp_stages_2_output_valid;
  assign IBusCachedPlugin_iBusRsp_stages_2_output_ready = IBusCachedPlugin_iBusRsp_output_ready;
  assign IBusCachedPlugin_iBusRsp_output_payload_rsp_inst = IBusCachedPlugin_cache_io_cpu_decode_data;
  assign IBusCachedPlugin_iBusRsp_output_payload_pc = IBusCachedPlugin_iBusRsp_stages_2_output_payload;
  assign IBusCachedPlugin_cache_io_flush = (decode_arbitration_isValid && decode_FLUSH_ALL);
  assign _zz_dBus_cmd_valid = 1'b0;
  always @(*) begin
    execute_DBusSimplePlugin_skipCmd = 1'b0;
    if(execute_ALIGNEMENT_FAULT) begin
      execute_DBusSimplePlugin_skipCmd = 1'b1;
    end
  end

  assign dBus_cmd_valid = (((((execute_arbitration_isValid && execute_MEMORY_ENABLE) && (! execute_arbitration_isStuckByOthers)) && (! execute_arbitration_isFlushed)) && (! execute_DBusSimplePlugin_skipCmd)) && (! _zz_dBus_cmd_valid));
  assign dBus_cmd_payload_wr = execute_MEMORY_STORE;
  assign dBus_cmd_payload_size = execute_INSTRUCTION[13 : 12];
  always @(*) begin
    case(dBus_cmd_payload_size)
      2'b00 : begin
        _zz_dBus_cmd_payload_data = {{{execute_RS2[7 : 0],execute_RS2[7 : 0]},execute_RS2[7 : 0]},execute_RS2[7 : 0]};
      end
      2'b01 : begin
        _zz_dBus_cmd_payload_data = {execute_RS2[15 : 0],execute_RS2[15 : 0]};
      end
      default : begin
        _zz_dBus_cmd_payload_data = execute_RS2[31 : 0];
      end
    endcase
  end

  assign dBus_cmd_payload_data = _zz_dBus_cmd_payload_data;
  assign when_DBusSimplePlugin_l426 = ((((execute_arbitration_isValid && execute_MEMORY_ENABLE) && (! dBus_cmd_ready)) && (! execute_DBusSimplePlugin_skipCmd)) && (! _zz_dBus_cmd_valid));
  always @(*) begin
    case(dBus_cmd_payload_size)
      2'b00 : begin
        _zz_execute_DBusSimplePlugin_formalMask = 4'b0001;
      end
      2'b01 : begin
        _zz_execute_DBusSimplePlugin_formalMask = 4'b0011;
      end
      default : begin
        _zz_execute_DBusSimplePlugin_formalMask = 4'b1111;
      end
    endcase
  end

  assign execute_DBusSimplePlugin_formalMask = (_zz_execute_DBusSimplePlugin_formalMask <<< dBus_cmd_payload_address[1 : 0]);
  assign dBus_cmd_payload_address = execute_SRC_ADD;
  assign when_DBusSimplePlugin_l479 = (((memory_arbitration_isValid && memory_MEMORY_ENABLE) && (! memory_MEMORY_STORE)) && ((! dBus_rsp_ready) || 1'b0));
  always @(*) begin
    DBusSimplePlugin_memoryExceptionPort_valid = 1'b0;
    if(when_DBusSimplePlugin_l486) begin
      DBusSimplePlugin_memoryExceptionPort_valid = 1'b1;
    end
    if(memory_ALIGNEMENT_FAULT) begin
      DBusSimplePlugin_memoryExceptionPort_valid = 1'b1;
    end
    if(when_DBusSimplePlugin_l512) begin
      DBusSimplePlugin_memoryExceptionPort_valid = 1'b0;
    end
  end

  always @(*) begin
    DBusSimplePlugin_memoryExceptionPort_payload_code = 4'bxxxx;
    if(when_DBusSimplePlugin_l486) begin
      DBusSimplePlugin_memoryExceptionPort_payload_code = 4'b0101;
    end
    if(memory_ALIGNEMENT_FAULT) begin
      DBusSimplePlugin_memoryExceptionPort_payload_code = {1'd0, _zz_DBusSimplePlugin_memoryExceptionPort_payload_code};
    end
  end

  assign DBusSimplePlugin_memoryExceptionPort_payload_badAddr = memory_REGFILE_WRITE_DATA;
  assign when_DBusSimplePlugin_l486 = ((dBus_rsp_ready && dBus_rsp_error) && (! memory_MEMORY_STORE));
  assign when_DBusSimplePlugin_l512 = (! ((memory_arbitration_isValid && memory_MEMORY_ENABLE) && (1'b1 || (! memory_arbitration_isStuckByOthers))));
  always @(*) begin
    writeBack_DBusSimplePlugin_rspShifted = writeBack_MEMORY_READ_DATA;
    case(writeBack_MEMORY_ADDRESS_LOW)
      2'b01 : begin
        writeBack_DBusSimplePlugin_rspShifted[7 : 0] = writeBack_MEMORY_READ_DATA[15 : 8];
      end
      2'b10 : begin
        writeBack_DBusSimplePlugin_rspShifted[15 : 0] = writeBack_MEMORY_READ_DATA[31 : 16];
      end
      2'b11 : begin
        writeBack_DBusSimplePlugin_rspShifted[7 : 0] = writeBack_MEMORY_READ_DATA[31 : 24];
      end
      default : begin
      end
    endcase
  end

  assign switch_Misc_l200 = writeBack_INSTRUCTION[13 : 12];
  assign _zz_writeBack_DBusSimplePlugin_rspFormated = (writeBack_DBusSimplePlugin_rspShifted[7] && (! writeBack_INSTRUCTION[14]));
  always @(*) begin
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[31] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[30] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[29] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[28] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[27] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[26] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[25] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[24] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[23] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[22] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[21] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[20] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[19] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[18] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[17] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[16] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[15] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[14] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[13] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[12] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[11] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[10] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[9] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[8] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[7 : 0] = writeBack_DBusSimplePlugin_rspShifted[7 : 0];
  end

  assign _zz_writeBack_DBusSimplePlugin_rspFormated_2 = (writeBack_DBusSimplePlugin_rspShifted[15] && (! writeBack_INSTRUCTION[14]));
  always @(*) begin
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[31] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[30] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[29] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[28] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[27] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[26] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[25] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[24] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[23] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[22] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[21] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[20] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[19] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[18] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[17] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[16] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[15 : 0] = writeBack_DBusSimplePlugin_rspShifted[15 : 0];
  end

  always @(*) begin
    case(switch_Misc_l200)
      2'b00 : begin
        writeBack_DBusSimplePlugin_rspFormated = _zz_writeBack_DBusSimplePlugin_rspFormated_1;
      end
      2'b01 : begin
        writeBack_DBusSimplePlugin_rspFormated = _zz_writeBack_DBusSimplePlugin_rspFormated_3;
      end
      default : begin
        writeBack_DBusSimplePlugin_rspFormated = writeBack_DBusSimplePlugin_rspShifted;
      end
    endcase
  end

  assign when_DBusSimplePlugin_l558 = (writeBack_arbitration_isValid && writeBack_MEMORY_ENABLE);
  assign IBusCachedPlugin_mmuBus_rsp_physicalAddress = IBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  assign IBusCachedPlugin_mmuBus_rsp_allowRead = 1'b1;
  assign IBusCachedPlugin_mmuBus_rsp_allowWrite = 1'b1;
  assign IBusCachedPlugin_mmuBus_rsp_allowExecute = 1'b1;
  assign IBusCachedPlugin_mmuBus_rsp_isIoAccess = IBusCachedPlugin_mmuBus_rsp_physicalAddress[31];
  assign IBusCachedPlugin_mmuBus_rsp_isPaging = 1'b0;
  assign IBusCachedPlugin_mmuBus_rsp_exception = 1'b0;
  assign IBusCachedPlugin_mmuBus_rsp_refilling = 1'b0;
  assign IBusCachedPlugin_mmuBus_busy = 1'b0;
  assign _zz_decode_ENV_CTRL_3 = ((decode_INSTRUCTION & 32'h00004050) == 32'h00004050);
  assign _zz_decode_ENV_CTRL_4 = ((decode_INSTRUCTION & 32'h00000004) == 32'h00000004);
  assign _zz_decode_ENV_CTRL_5 = ((decode_INSTRUCTION & 32'h00000050) == 32'h00000010);
  assign _zz_decode_ENV_CTRL_6 = ((decode_INSTRUCTION & 32'h00000048) == 32'h00000048);
  assign _zz_decode_ENV_CTRL_2 = {(((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2) == 32'h00100050) != 1'b0),{((_zz__zz_decode_ENV_CTRL_2_1 == _zz__zz_decode_ENV_CTRL_2_2) != 1'b0),{(_zz__zz_decode_ENV_CTRL_2_3 != 1'b0),{(_zz__zz_decode_ENV_CTRL_2_4 != _zz__zz_decode_ENV_CTRL_2_9),{_zz__zz_decode_ENV_CTRL_2_10,{_zz__zz_decode_ENV_CTRL_2_12,_zz__zz_decode_ENV_CTRL_2_14}}}}}};
  assign _zz_decode_SRC1_CTRL_2 = _zz_decode_ENV_CTRL_2[2 : 1];
  assign _zz_decode_SRC1_CTRL_1 = _zz_decode_SRC1_CTRL_2;
  assign _zz_decode_ALU_CTRL_2 = _zz_decode_ENV_CTRL_2[7 : 6];
  assign _zz_decode_ALU_CTRL_1 = _zz_decode_ALU_CTRL_2;
  assign _zz_decode_SRC2_CTRL_2 = _zz_decode_ENV_CTRL_2[9 : 8];
  assign _zz_decode_SRC2_CTRL_1 = _zz_decode_SRC2_CTRL_2;
  assign _zz_decode_ALU_BITWISE_CTRL_2 = _zz_decode_ENV_CTRL_2[18 : 17];
  assign _zz_decode_ALU_BITWISE_CTRL_1 = _zz_decode_ALU_BITWISE_CTRL_2;
  assign _zz_decode_SHIFT_CTRL_2 = _zz_decode_ENV_CTRL_2[21 : 20];
  assign _zz_decode_SHIFT_CTRL_1 = _zz_decode_SHIFT_CTRL_2;
  assign _zz_decode_BRANCH_CTRL_2 = _zz_decode_ENV_CTRL_2[23 : 22];
  assign _zz_decode_BRANCH_CTRL_1 = _zz_decode_BRANCH_CTRL_2;
  assign _zz_decode_ENV_CTRL_7 = _zz_decode_ENV_CTRL_2[26 : 25];
  assign _zz_decode_ENV_CTRL_1 = _zz_decode_ENV_CTRL_7;
  assign decodeExceptionPort_valid = (decode_arbitration_isValid && (! decode_LEGAL_INSTRUCTION));
  assign decodeExceptionPort_payload_code = 4'b0010;
  assign decodeExceptionPort_payload_badAddr = decode_INSTRUCTION;
  assign when_RegFilePlugin_l63 = (decode_INSTRUCTION[11 : 7] == 5'h0);
  assign decode_RegFilePlugin_regFileReadAddress1 = decode_INSTRUCTION_ANTICIPATED[19 : 15];
  assign decode_RegFilePlugin_regFileReadAddress2 = decode_INSTRUCTION_ANTICIPATED[24 : 20];
  assign decode_RegFilePlugin_rs1Data = _zz_RegFilePlugin_regFile_port0;
  assign decode_RegFilePlugin_rs2Data = _zz_RegFilePlugin_regFile_port1;
  always @(*) begin
    lastStageRegFileWrite_valid = (_zz_lastStageRegFileWrite_valid && writeBack_arbitration_isFiring);
    if(_zz_2) begin
      lastStageRegFileWrite_valid = 1'b1;
    end
  end

  always @(*) begin
    lastStageRegFileWrite_payload_address = _zz_lastStageRegFileWrite_payload_address[11 : 7];
    if(_zz_2) begin
      lastStageRegFileWrite_payload_address = 5'h0;
    end
  end

  always @(*) begin
    lastStageRegFileWrite_payload_data = _zz_lastStageRegFileWrite_payload_data;
    if(_zz_2) begin
      lastStageRegFileWrite_payload_data = 32'h0;
    end
  end

  always @(*) begin
    case(execute_ALU_BITWISE_CTRL)
      `AluBitwiseCtrlEnum_binary_sequential_AND_1 : begin
        execute_IntAluPlugin_bitwise = (execute_SRC1 & execute_SRC2);
      end
      `AluBitwiseCtrlEnum_binary_sequential_OR_1 : begin
        execute_IntAluPlugin_bitwise = (execute_SRC1 | execute_SRC2);
      end
      default : begin
        execute_IntAluPlugin_bitwise = (execute_SRC1 ^ execute_SRC2);
      end
    endcase
  end

  always @(*) begin
    case(execute_ALU_CTRL)
      `AluCtrlEnum_binary_sequential_BITWISE : begin
        _zz_execute_REGFILE_WRITE_DATA = execute_IntAluPlugin_bitwise;
      end
      `AluCtrlEnum_binary_sequential_SLT_SLTU : begin
        _zz_execute_REGFILE_WRITE_DATA = {31'd0, _zz__zz_execute_REGFILE_WRITE_DATA};
      end
      default : begin
        _zz_execute_REGFILE_WRITE_DATA = execute_SRC_ADD_SUB;
      end
    endcase
  end

  always @(*) begin
    case(execute_SRC1_CTRL)
      `Src1CtrlEnum_binary_sequential_RS : begin
        _zz_execute_SRC1 = execute_RS1;
      end
      `Src1CtrlEnum_binary_sequential_PC_INCREMENT : begin
        _zz_execute_SRC1 = {29'd0, _zz__zz_execute_SRC1};
      end
      `Src1CtrlEnum_binary_sequential_IMU : begin
        _zz_execute_SRC1 = {execute_INSTRUCTION[31 : 12],12'h0};
      end
      default : begin
        _zz_execute_SRC1 = {27'd0, _zz__zz_execute_SRC1_1};
      end
    endcase
  end

  assign _zz_execute_SRC2_1 = execute_INSTRUCTION[31];
  always @(*) begin
    _zz_execute_SRC2_2[19] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[18] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[17] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[16] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[15] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[14] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[13] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[12] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[11] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[10] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[9] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[8] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[7] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[6] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[5] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[4] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[3] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[2] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[1] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[0] = _zz_execute_SRC2_1;
  end

  assign _zz_execute_SRC2_3 = _zz__zz_execute_SRC2_3[11];
  always @(*) begin
    _zz_execute_SRC2_4[19] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[18] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[17] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[16] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[15] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[14] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[13] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[12] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[11] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[10] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[9] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[8] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[7] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[6] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[5] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[4] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[3] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[2] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[1] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[0] = _zz_execute_SRC2_3;
  end

  always @(*) begin
    case(execute_SRC2_CTRL)
      `Src2CtrlEnum_binary_sequential_RS : begin
        _zz_execute_SRC2_5 = execute_RS2;
      end
      `Src2CtrlEnum_binary_sequential_IMI : begin
        _zz_execute_SRC2_5 = {_zz_execute_SRC2_2,execute_INSTRUCTION[31 : 20]};
      end
      `Src2CtrlEnum_binary_sequential_IMS : begin
        _zz_execute_SRC2_5 = {_zz_execute_SRC2_4,{execute_INSTRUCTION[31 : 25],execute_INSTRUCTION[11 : 7]}};
      end
      default : begin
        _zz_execute_SRC2_5 = _zz_execute_SRC2;
      end
    endcase
  end

  always @(*) begin
    execute_SrcPlugin_addSub = _zz_execute_SrcPlugin_addSub;
    if(execute_SRC2_FORCE_ZERO) begin
      execute_SrcPlugin_addSub = execute_SRC1;
    end
  end

  assign execute_SrcPlugin_less = ((execute_SRC1[31] == execute_SRC2[31]) ? execute_SrcPlugin_addSub[31] : (execute_SRC_LESS_UNSIGNED ? execute_SRC2[31] : execute_SRC1[31]));
  assign execute_LightShifterPlugin_isShift = (execute_SHIFT_CTRL != `ShiftCtrlEnum_binary_sequential_DISABLE_1);
  assign execute_LightShifterPlugin_amplitude = (execute_LightShifterPlugin_isActive ? execute_LightShifterPlugin_amplitudeReg : execute_SRC2[4 : 0]);
  assign execute_LightShifterPlugin_shiftInput = (execute_LightShifterPlugin_isActive ? memory_REGFILE_WRITE_DATA : execute_SRC1);
  assign execute_LightShifterPlugin_done = (execute_LightShifterPlugin_amplitude[4 : 1] == 4'b0000);
  assign when_ShiftPlugins_l169 = ((execute_arbitration_isValid && execute_LightShifterPlugin_isShift) && (execute_SRC2[4 : 0] != 5'h0));
  always @(*) begin
    case(execute_SHIFT_CTRL)
      `ShiftCtrlEnum_binary_sequential_SLL_1 : begin
        _zz_execute_to_memory_REGFILE_WRITE_DATA_1 = (execute_LightShifterPlugin_shiftInput <<< 1);
      end
      default : begin
        _zz_execute_to_memory_REGFILE_WRITE_DATA_1 = _zz__zz_execute_to_memory_REGFILE_WRITE_DATA_1;
      end
    endcase
  end

  assign when_ShiftPlugins_l175 = (! execute_arbitration_isStuckByOthers);
  assign when_ShiftPlugins_l184 = (! execute_LightShifterPlugin_done);
  always @(*) begin
    HazardSimplePlugin_src0Hazard = 1'b0;
    if(HazardSimplePlugin_writeBackBuffer_valid) begin
      if(HazardSimplePlugin_addr0Match) begin
        HazardSimplePlugin_src0Hazard = 1'b1;
      end
    end
    if(when_HazardSimplePlugin_l57) begin
      if(when_HazardSimplePlugin_l58) begin
        if(when_HazardSimplePlugin_l59) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_1) begin
      if(when_HazardSimplePlugin_l58_1) begin
        if(when_HazardSimplePlugin_l59_1) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_2) begin
      if(when_HazardSimplePlugin_l58_2) begin
        if(when_HazardSimplePlugin_l59_2) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l105) begin
      HazardSimplePlugin_src0Hazard = 1'b0;
    end
  end

  always @(*) begin
    HazardSimplePlugin_src1Hazard = 1'b0;
    if(HazardSimplePlugin_writeBackBuffer_valid) begin
      if(HazardSimplePlugin_addr1Match) begin
        HazardSimplePlugin_src1Hazard = 1'b1;
      end
    end
    if(when_HazardSimplePlugin_l57) begin
      if(when_HazardSimplePlugin_l58) begin
        if(when_HazardSimplePlugin_l62) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_1) begin
      if(when_HazardSimplePlugin_l58_1) begin
        if(when_HazardSimplePlugin_l62_1) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_2) begin
      if(when_HazardSimplePlugin_l58_2) begin
        if(when_HazardSimplePlugin_l62_2) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l108) begin
      HazardSimplePlugin_src1Hazard = 1'b0;
    end
  end

  assign HazardSimplePlugin_writeBackWrites_valid = (_zz_lastStageRegFileWrite_valid && writeBack_arbitration_isFiring);
  assign HazardSimplePlugin_writeBackWrites_payload_address = _zz_lastStageRegFileWrite_payload_address[11 : 7];
  assign HazardSimplePlugin_writeBackWrites_payload_data = _zz_lastStageRegFileWrite_payload_data;
  assign HazardSimplePlugin_addr0Match = (HazardSimplePlugin_writeBackBuffer_payload_address == decode_INSTRUCTION[19 : 15]);
  assign HazardSimplePlugin_addr1Match = (HazardSimplePlugin_writeBackBuffer_payload_address == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l59 = (writeBack_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l62 = (writeBack_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l57 = (writeBack_arbitration_isValid && writeBack_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58 = (1'b1 || (! 1'b1));
  assign when_HazardSimplePlugin_l59_1 = (memory_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l62_1 = (memory_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l57_1 = (memory_arbitration_isValid && memory_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58_1 = (1'b1 || (! memory_BYPASSABLE_MEMORY_STAGE));
  assign when_HazardSimplePlugin_l59_2 = (execute_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l62_2 = (execute_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l57_2 = (execute_arbitration_isValid && execute_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58_2 = (1'b1 || (! execute_BYPASSABLE_EXECUTE_STAGE));
  assign when_HazardSimplePlugin_l105 = (! decode_RS1_USE);
  assign when_HazardSimplePlugin_l108 = (! decode_RS2_USE);
  assign when_HazardSimplePlugin_l113 = (decode_arbitration_isValid && (HazardSimplePlugin_src0Hazard || HazardSimplePlugin_src1Hazard));
  assign execute_BranchPlugin_eq = (execute_SRC1 == execute_SRC2);
  assign switch_Misc_l200_1 = execute_INSTRUCTION[14 : 12];
  always @(*) begin
    casez(switch_Misc_l200_1)
      3'b000 : begin
        _zz_execute_BRANCH_DO = execute_BranchPlugin_eq;
      end
      3'b001 : begin
        _zz_execute_BRANCH_DO = (! execute_BranchPlugin_eq);
      end
      3'b1?1 : begin
        _zz_execute_BRANCH_DO = (! execute_SRC_LESS);
      end
      default : begin
        _zz_execute_BRANCH_DO = execute_SRC_LESS;
      end
    endcase
  end

  always @(*) begin
    case(execute_BRANCH_CTRL)
      `BranchCtrlEnum_binary_sequential_INC : begin
        _zz_execute_BRANCH_DO_1 = 1'b0;
      end
      `BranchCtrlEnum_binary_sequential_JAL : begin
        _zz_execute_BRANCH_DO_1 = 1'b1;
      end
      `BranchCtrlEnum_binary_sequential_JALR : begin
        _zz_execute_BRANCH_DO_1 = 1'b1;
      end
      default : begin
        _zz_execute_BRANCH_DO_1 = _zz_execute_BRANCH_DO;
      end
    endcase
  end

  assign execute_BranchPlugin_branch_src1 = ((execute_BRANCH_CTRL == `BranchCtrlEnum_binary_sequential_JALR) ? execute_RS1 : execute_PC);
  assign _zz_execute_BranchPlugin_branch_src2 = _zz__zz_execute_BranchPlugin_branch_src2[19];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_1[10] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[9] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[8] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[7] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[6] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[5] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[4] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[3] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[2] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[1] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[0] = _zz_execute_BranchPlugin_branch_src2;
  end

  assign _zz_execute_BranchPlugin_branch_src2_2 = execute_INSTRUCTION[31];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_3[19] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[18] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[17] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[16] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[15] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[14] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[13] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[12] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[11] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[10] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[9] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[8] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[7] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[6] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[5] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[4] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[3] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[2] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[1] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[0] = _zz_execute_BranchPlugin_branch_src2_2;
  end

  assign _zz_execute_BranchPlugin_branch_src2_4 = _zz__zz_execute_BranchPlugin_branch_src2_4[11];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_5[18] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[17] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[16] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[15] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[14] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[13] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[12] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[11] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[10] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[9] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[8] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[7] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[6] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[5] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[4] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[3] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[2] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[1] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[0] = _zz_execute_BranchPlugin_branch_src2_4;
  end

  always @(*) begin
    case(execute_BRANCH_CTRL)
      `BranchCtrlEnum_binary_sequential_JAL : begin
        _zz_execute_BranchPlugin_branch_src2_6 = {{_zz_execute_BranchPlugin_branch_src2_1,{{{execute_INSTRUCTION[31],execute_INSTRUCTION[19 : 12]},execute_INSTRUCTION[20]},execute_INSTRUCTION[30 : 21]}},1'b0};
      end
      `BranchCtrlEnum_binary_sequential_JALR : begin
        _zz_execute_BranchPlugin_branch_src2_6 = {_zz_execute_BranchPlugin_branch_src2_3,execute_INSTRUCTION[31 : 20]};
      end
      default : begin
        _zz_execute_BranchPlugin_branch_src2_6 = {{_zz_execute_BranchPlugin_branch_src2_5,{{{execute_INSTRUCTION[31],execute_INSTRUCTION[7]},execute_INSTRUCTION[30 : 25]},execute_INSTRUCTION[11 : 8]}},1'b0};
      end
    endcase
  end

  assign execute_BranchPlugin_branch_src2 = _zz_execute_BranchPlugin_branch_src2_6;
  assign execute_BranchPlugin_branchAdder = (execute_BranchPlugin_branch_src1 + execute_BranchPlugin_branch_src2);
  assign BranchPlugin_jumpInterface_valid = ((memory_arbitration_isValid && memory_BRANCH_DO) && (! 1'b0));
  assign BranchPlugin_jumpInterface_payload = memory_BRANCH_CALC;
  assign BranchPlugin_branchExceptionPort_valid = ((memory_arbitration_isValid && memory_BRANCH_DO) && BranchPlugin_jumpInterface_payload[1]);
  assign BranchPlugin_branchExceptionPort_payload_code = 4'b0000;
  assign BranchPlugin_branchExceptionPort_payload_badAddr = BranchPlugin_jumpInterface_payload;
  always @(*) begin
    CsrPlugin_privilege = 2'b11;
    if(CsrPlugin_forceMachineWire) begin
      CsrPlugin_privilege = 2'b11;
    end
  end

  assign CsrPlugin_misa_base = 2'b01;
  assign CsrPlugin_misa_extensions = 26'h0000042;
  assign _zz_when_CsrPlugin_l952 = (CsrPlugin_mip_MTIP && CsrPlugin_mie_MTIE);
  assign _zz_when_CsrPlugin_l952_1 = (CsrPlugin_mip_MSIP && CsrPlugin_mie_MSIE);
  assign _zz_when_CsrPlugin_l952_2 = (CsrPlugin_mip_MEIP && CsrPlugin_mie_MEIE);
  assign CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped = 2'b11;
  assign CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege = ((CsrPlugin_privilege < CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped) ? CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped : CsrPlugin_privilege);
  assign _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code = {decodeExceptionPort_valid,IBusCachedPlugin_decodeExceptionPort_valid};
  assign _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 = _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1[0];
  assign _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_2 = {BranchPlugin_branchExceptionPort_valid,DBusSimplePlugin_memoryExceptionPort_valid};
  assign _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3 = _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3[0];
  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_decode = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
    if(_zz_when) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_decode = 1'b1;
    end
    if(decode_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_decode = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_execute = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
    if(CsrPlugin_selfException_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_execute = 1'b1;
    end
    if(execute_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_execute = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_memory = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
    if(_zz_when_1) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_memory = 1'b1;
    end
    if(memory_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_memory = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
    if(writeBack_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack = 1'b0;
    end
  end

  assign when_CsrPlugin_l909 = (! decode_arbitration_isStuck);
  assign when_CsrPlugin_l909_1 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l909_2 = (! memory_arbitration_isStuck);
  assign when_CsrPlugin_l909_3 = (! writeBack_arbitration_isStuck);
  assign when_CsrPlugin_l922 = ({CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack,{CsrPlugin_exceptionPortCtrl_exceptionValids_memory,{CsrPlugin_exceptionPortCtrl_exceptionValids_execute,CsrPlugin_exceptionPortCtrl_exceptionValids_decode}}} != 4'b0000);
  assign CsrPlugin_exceptionPendings_0 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
  assign CsrPlugin_exceptionPendings_1 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
  assign CsrPlugin_exceptionPendings_2 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
  assign CsrPlugin_exceptionPendings_3 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
  assign when_CsrPlugin_l946 = (CsrPlugin_mstatus_MIE || (CsrPlugin_privilege < 2'b11));
  assign when_CsrPlugin_l952 = ((_zz_when_CsrPlugin_l952 && 1'b1) && (! 1'b0));
  assign when_CsrPlugin_l952_1 = ((_zz_when_CsrPlugin_l952_1 && 1'b1) && (! 1'b0));
  assign when_CsrPlugin_l952_2 = ((_zz_when_CsrPlugin_l952_2 && 1'b1) && (! 1'b0));
  assign CsrPlugin_exception = (CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack && CsrPlugin_allowException);
  assign CsrPlugin_lastStageWasWfi = 1'b0;
  assign CsrPlugin_pipelineLiberator_active = ((CsrPlugin_interrupt_valid && CsrPlugin_allowInterrupts) && decode_arbitration_isValid);
  assign when_CsrPlugin_l980 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l980_1 = (! memory_arbitration_isStuck);
  assign when_CsrPlugin_l980_2 = (! writeBack_arbitration_isStuck);
  assign when_CsrPlugin_l985 = ((! CsrPlugin_pipelineLiberator_active) || decode_arbitration_removeIt);
  always @(*) begin
    CsrPlugin_pipelineLiberator_done = CsrPlugin_pipelineLiberator_pcValids_2;
    if(when_CsrPlugin_l991) begin
      CsrPlugin_pipelineLiberator_done = 1'b0;
    end
    if(CsrPlugin_hadException) begin
      CsrPlugin_pipelineLiberator_done = 1'b0;
    end
  end

  assign when_CsrPlugin_l991 = ({CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack,{CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory,CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute}} != 3'b000);
  assign CsrPlugin_interruptJump = ((CsrPlugin_interrupt_valid && CsrPlugin_pipelineLiberator_done) && CsrPlugin_allowInterrupts);
  always @(*) begin
    CsrPlugin_targetPrivilege = CsrPlugin_interrupt_targetPrivilege;
    if(CsrPlugin_hadException) begin
      CsrPlugin_targetPrivilege = CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege;
    end
  end

  always @(*) begin
    CsrPlugin_trapCause = CsrPlugin_interrupt_code;
    if(CsrPlugin_hadException) begin
      CsrPlugin_trapCause = CsrPlugin_exceptionPortCtrl_exceptionContext_code;
    end
  end

  always @(*) begin
    CsrPlugin_xtvec_mode = 2'bxx;
    case(CsrPlugin_targetPrivilege)
      2'b11 : begin
        CsrPlugin_xtvec_mode = CsrPlugin_mtvec_mode;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrPlugin_xtvec_base = 30'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(CsrPlugin_targetPrivilege)
      2'b11 : begin
        CsrPlugin_xtvec_base = CsrPlugin_mtvec_base;
      end
      default : begin
      end
    endcase
  end

  assign when_CsrPlugin_l1019 = (CsrPlugin_hadException || CsrPlugin_interruptJump);
  assign when_CsrPlugin_l1064 = (writeBack_arbitration_isValid && (writeBack_ENV_CTRL == `EnvCtrlEnum_binary_sequential_XRET));
  assign switch_CsrPlugin_l1068 = writeBack_INSTRUCTION[29 : 28];
  assign contextSwitching = CsrPlugin_jumpInterface_valid;
  assign when_CsrPlugin_l1116 = ({(writeBack_arbitration_isValid && (writeBack_ENV_CTRL == `EnvCtrlEnum_binary_sequential_XRET)),{(memory_arbitration_isValid && (memory_ENV_CTRL == `EnvCtrlEnum_binary_sequential_XRET)),(execute_arbitration_isValid && (execute_ENV_CTRL == `EnvCtrlEnum_binary_sequential_XRET))}} != 3'b000);
  assign execute_CsrPlugin_blockedBySideEffects = (({writeBack_arbitration_isValid,memory_arbitration_isValid} != 2'b00) || 1'b0);
  always @(*) begin
    execute_CsrPlugin_illegalAccess = 1'b1;
    if(execute_CsrPlugin_csr_768) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_836) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_772) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_773) begin
      if(execute_CSR_WRITE_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_833) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_834) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_835) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3008) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_4032) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(CsrPlugin_csrMapping_allowCsrSignal) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(when_CsrPlugin_l1297) begin
      execute_CsrPlugin_illegalAccess = 1'b1;
    end
    if(when_CsrPlugin_l1302) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
  end

  always @(*) begin
    execute_CsrPlugin_illegalInstruction = 1'b0;
    if(when_CsrPlugin_l1136) begin
      if(when_CsrPlugin_l1137) begin
        execute_CsrPlugin_illegalInstruction = 1'b1;
      end
    end
  end

  always @(*) begin
    CsrPlugin_selfException_valid = 1'b0;
    if(when_CsrPlugin_l1144) begin
      CsrPlugin_selfException_valid = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_selfException_payload_code = 4'bxxxx;
    if(when_CsrPlugin_l1144) begin
      case(CsrPlugin_privilege)
        2'b00 : begin
          CsrPlugin_selfException_payload_code = 4'b1000;
        end
        default : begin
          CsrPlugin_selfException_payload_code = 4'b1011;
        end
      endcase
    end
  end

  assign CsrPlugin_selfException_payload_badAddr = execute_INSTRUCTION;
  assign when_CsrPlugin_l1136 = (execute_arbitration_isValid && (execute_ENV_CTRL == `EnvCtrlEnum_binary_sequential_XRET));
  assign when_CsrPlugin_l1137 = (CsrPlugin_privilege < execute_INSTRUCTION[29 : 28]);
  assign when_CsrPlugin_l1144 = (execute_arbitration_isValid && (execute_ENV_CTRL == `EnvCtrlEnum_binary_sequential_ECALL));
  always @(*) begin
    execute_CsrPlugin_writeInstruction = ((execute_arbitration_isValid && execute_IS_CSR) && execute_CSR_WRITE_OPCODE);
    if(when_CsrPlugin_l1297) begin
      execute_CsrPlugin_writeInstruction = 1'b0;
    end
  end

  always @(*) begin
    execute_CsrPlugin_readInstruction = ((execute_arbitration_isValid && execute_IS_CSR) && execute_CSR_READ_OPCODE);
    if(when_CsrPlugin_l1297) begin
      execute_CsrPlugin_readInstruction = 1'b0;
    end
  end

  assign execute_CsrPlugin_writeEnable = (execute_CsrPlugin_writeInstruction && (! execute_arbitration_isStuck));
  assign execute_CsrPlugin_readEnable = (execute_CsrPlugin_readInstruction && (! execute_arbitration_isStuck));
  assign CsrPlugin_csrMapping_hazardFree = (! execute_CsrPlugin_blockedBySideEffects);
  assign execute_CsrPlugin_readToWriteData = CsrPlugin_csrMapping_readDataSignal;
  assign switch_Misc_l200_2 = execute_INSTRUCTION[13];
  always @(*) begin
    case(switch_Misc_l200_2)
      1'b0 : begin
        _zz_CsrPlugin_csrMapping_writeDataSignal = execute_SRC1;
      end
      default : begin
        _zz_CsrPlugin_csrMapping_writeDataSignal = (execute_INSTRUCTION[12] ? (execute_CsrPlugin_readToWriteData & (~ execute_SRC1)) : (execute_CsrPlugin_readToWriteData | execute_SRC1));
      end
    endcase
  end

  assign CsrPlugin_csrMapping_writeDataSignal = _zz_CsrPlugin_csrMapping_writeDataSignal;
  assign when_CsrPlugin_l1176 = (execute_arbitration_isValid && execute_IS_CSR);
  assign when_CsrPlugin_l1180 = (execute_arbitration_isValid && (execute_IS_CSR || 1'b0));
  assign execute_CsrPlugin_csrAddress = execute_INSTRUCTION[31 : 20];
  assign _zz_CsrPlugin_csrMapping_readDataInit_1 = (_zz_CsrPlugin_csrMapping_readDataInit & externalInterruptArray_regNext);
  assign externalInterrupt = (_zz_CsrPlugin_csrMapping_readDataInit_1 != 32'h0);
  assign when_DebugPlugin_l225 = (DebugPlugin_haltIt && (! DebugPlugin_isPipBusy));
  assign DebugPlugin_allowEBreak = (DebugPlugin_debugUsed && (! DebugPlugin_disableEbreak));
  always @(*) begin
    debug_bus_cmd_ready = 1'b1;
    if(debug_bus_cmd_valid) begin
      case(switch_DebugPlugin_l256)
        6'h01 : begin
          if(debug_bus_cmd_payload_wr) begin
            debug_bus_cmd_ready = IBusCachedPlugin_injectionPort_ready;
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    debug_bus_rsp_data = DebugPlugin_busReadDataReg;
    if(when_DebugPlugin_l244) begin
      debug_bus_rsp_data[0] = DebugPlugin_resetIt;
      debug_bus_rsp_data[1] = DebugPlugin_haltIt;
      debug_bus_rsp_data[2] = DebugPlugin_isPipBusy;
      debug_bus_rsp_data[3] = DebugPlugin_haltedByBreak;
      debug_bus_rsp_data[4] = DebugPlugin_stepIt;
    end
  end

  assign when_DebugPlugin_l244 = (! _zz_when_DebugPlugin_l244);
  always @(*) begin
    IBusCachedPlugin_injectionPort_valid = 1'b0;
    if(debug_bus_cmd_valid) begin
      case(switch_DebugPlugin_l256)
        6'h01 : begin
          if(debug_bus_cmd_payload_wr) begin
            IBusCachedPlugin_injectionPort_valid = 1'b1;
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign IBusCachedPlugin_injectionPort_payload = debug_bus_cmd_payload_data;
  assign switch_DebugPlugin_l256 = debug_bus_cmd_payload_address[7 : 2];
  assign when_DebugPlugin_l260 = debug_bus_cmd_payload_data[16];
  assign when_DebugPlugin_l260_1 = debug_bus_cmd_payload_data[24];
  assign when_DebugPlugin_l261 = debug_bus_cmd_payload_data[17];
  assign when_DebugPlugin_l261_1 = debug_bus_cmd_payload_data[25];
  assign when_DebugPlugin_l262 = debug_bus_cmd_payload_data[25];
  assign when_DebugPlugin_l263 = debug_bus_cmd_payload_data[25];
  assign when_DebugPlugin_l264 = debug_bus_cmd_payload_data[18];
  assign when_DebugPlugin_l264_1 = debug_bus_cmd_payload_data[26];
  assign when_DebugPlugin_l284 = (execute_arbitration_isValid && execute_DO_EBREAK);
  assign when_DebugPlugin_l287 = (({writeBack_arbitration_isValid,memory_arbitration_isValid} != 2'b00) == 1'b0);
  assign when_DebugPlugin_l300 = (DebugPlugin_stepIt && IBusCachedPlugin_incomingInstruction);
  assign debug_resetOut = DebugPlugin_resetIt_regNext;
  assign when_DebugPlugin_l316 = (DebugPlugin_haltIt || DebugPlugin_stepIt);
  assign when_Pipeline_l124 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_1 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_2 = ((! writeBack_arbitration_isStuck) && (! CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack));
  assign when_Pipeline_l124_3 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_4 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_5 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_6 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_7 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_8 = (! writeBack_arbitration_isStuck);
  assign _zz_decode_to_execute_SRC1_CTRL_1 = decode_SRC1_CTRL;
  assign _zz_decode_SRC1_CTRL = _zz_decode_SRC1_CTRL_1;
  assign when_Pipeline_l124_9 = (! execute_arbitration_isStuck);
  assign _zz_execute_SRC1_CTRL = decode_to_execute_SRC1_CTRL;
  assign when_Pipeline_l124_10 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_11 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_12 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_13 = (! writeBack_arbitration_isStuck);
  assign _zz_decode_to_execute_ALU_CTRL_1 = decode_ALU_CTRL;
  assign _zz_decode_ALU_CTRL = _zz_decode_ALU_CTRL_1;
  assign when_Pipeline_l124_14 = (! execute_arbitration_isStuck);
  assign _zz_execute_ALU_CTRL = decode_to_execute_ALU_CTRL;
  assign _zz_decode_to_execute_SRC2_CTRL_1 = decode_SRC2_CTRL;
  assign _zz_decode_SRC2_CTRL = _zz_decode_SRC2_CTRL_1;
  assign when_Pipeline_l124_15 = (! execute_arbitration_isStuck);
  assign _zz_execute_SRC2_CTRL = decode_to_execute_SRC2_CTRL;
  assign when_Pipeline_l124_16 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_17 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_18 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_19 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_20 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_21 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_22 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_23 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_24 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_25 = (! execute_arbitration_isStuck);
  assign _zz_decode_to_execute_ALU_BITWISE_CTRL_1 = decode_ALU_BITWISE_CTRL;
  assign _zz_decode_ALU_BITWISE_CTRL = _zz_decode_ALU_BITWISE_CTRL_1;
  assign when_Pipeline_l124_26 = (! execute_arbitration_isStuck);
  assign _zz_execute_ALU_BITWISE_CTRL = decode_to_execute_ALU_BITWISE_CTRL;
  assign _zz_decode_to_execute_SHIFT_CTRL_1 = decode_SHIFT_CTRL;
  assign _zz_decode_SHIFT_CTRL = _zz_decode_SHIFT_CTRL_1;
  assign when_Pipeline_l124_27 = (! execute_arbitration_isStuck);
  assign _zz_execute_SHIFT_CTRL = decode_to_execute_SHIFT_CTRL;
  assign _zz_decode_to_execute_BRANCH_CTRL_1 = decode_BRANCH_CTRL;
  assign _zz_decode_BRANCH_CTRL = _zz_decode_BRANCH_CTRL_1;
  assign when_Pipeline_l124_28 = (! execute_arbitration_isStuck);
  assign _zz_execute_BRANCH_CTRL = decode_to_execute_BRANCH_CTRL;
  assign when_Pipeline_l124_29 = (! execute_arbitration_isStuck);
  assign _zz_decode_to_execute_ENV_CTRL_1 = decode_ENV_CTRL;
  assign _zz_execute_to_memory_ENV_CTRL_1 = execute_ENV_CTRL;
  assign _zz_memory_to_writeBack_ENV_CTRL_1 = memory_ENV_CTRL;
  assign _zz_decode_ENV_CTRL = _zz_decode_ENV_CTRL_1;
  assign when_Pipeline_l124_30 = (! execute_arbitration_isStuck);
  assign _zz_execute_ENV_CTRL = decode_to_execute_ENV_CTRL;
  assign when_Pipeline_l124_31 = (! memory_arbitration_isStuck);
  assign _zz_memory_ENV_CTRL = execute_to_memory_ENV_CTRL;
  assign when_Pipeline_l124_32 = (! writeBack_arbitration_isStuck);
  assign _zz_writeBack_ENV_CTRL = memory_to_writeBack_ENV_CTRL;
  assign when_Pipeline_l124_33 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_34 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_35 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_36 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_37 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_38 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_39 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_40 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_41 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_42 = ((! memory_arbitration_isStuck) && (! execute_arbitration_isStuckByOthers));
  assign when_Pipeline_l124_43 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_44 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_45 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_46 = (! writeBack_arbitration_isStuck);
  assign decode_arbitration_isFlushed = (({writeBack_arbitration_flushNext,{memory_arbitration_flushNext,execute_arbitration_flushNext}} != 3'b000) || ({writeBack_arbitration_flushIt,{memory_arbitration_flushIt,{execute_arbitration_flushIt,decode_arbitration_flushIt}}} != 4'b0000));
  assign execute_arbitration_isFlushed = (({writeBack_arbitration_flushNext,memory_arbitration_flushNext} != 2'b00) || ({writeBack_arbitration_flushIt,{memory_arbitration_flushIt,execute_arbitration_flushIt}} != 3'b000));
  assign memory_arbitration_isFlushed = ((writeBack_arbitration_flushNext != 1'b0) || ({writeBack_arbitration_flushIt,memory_arbitration_flushIt} != 2'b00));
  assign writeBack_arbitration_isFlushed = (1'b0 || (writeBack_arbitration_flushIt != 1'b0));
  assign decode_arbitration_isStuckByOthers = (decode_arbitration_haltByOther || (((1'b0 || execute_arbitration_isStuck) || memory_arbitration_isStuck) || writeBack_arbitration_isStuck));
  assign decode_arbitration_isStuck = (decode_arbitration_haltItself || decode_arbitration_isStuckByOthers);
  assign decode_arbitration_isMoving = ((! decode_arbitration_isStuck) && (! decode_arbitration_removeIt));
  assign decode_arbitration_isFiring = ((decode_arbitration_isValid && (! decode_arbitration_isStuck)) && (! decode_arbitration_removeIt));
  assign execute_arbitration_isStuckByOthers = (execute_arbitration_haltByOther || ((1'b0 || memory_arbitration_isStuck) || writeBack_arbitration_isStuck));
  assign execute_arbitration_isStuck = (execute_arbitration_haltItself || execute_arbitration_isStuckByOthers);
  assign execute_arbitration_isMoving = ((! execute_arbitration_isStuck) && (! execute_arbitration_removeIt));
  assign execute_arbitration_isFiring = ((execute_arbitration_isValid && (! execute_arbitration_isStuck)) && (! execute_arbitration_removeIt));
  assign memory_arbitration_isStuckByOthers = (memory_arbitration_haltByOther || (1'b0 || writeBack_arbitration_isStuck));
  assign memory_arbitration_isStuck = (memory_arbitration_haltItself || memory_arbitration_isStuckByOthers);
  assign memory_arbitration_isMoving = ((! memory_arbitration_isStuck) && (! memory_arbitration_removeIt));
  assign memory_arbitration_isFiring = ((memory_arbitration_isValid && (! memory_arbitration_isStuck)) && (! memory_arbitration_removeIt));
  assign writeBack_arbitration_isStuckByOthers = (writeBack_arbitration_haltByOther || 1'b0);
  assign writeBack_arbitration_isStuck = (writeBack_arbitration_haltItself || writeBack_arbitration_isStuckByOthers);
  assign writeBack_arbitration_isMoving = ((! writeBack_arbitration_isStuck) && (! writeBack_arbitration_removeIt));
  assign writeBack_arbitration_isFiring = ((writeBack_arbitration_isValid && (! writeBack_arbitration_isStuck)) && (! writeBack_arbitration_removeIt));
  assign when_Pipeline_l151 = ((! execute_arbitration_isStuck) || execute_arbitration_removeIt);
  assign when_Pipeline_l154 = ((! decode_arbitration_isStuck) && (! decode_arbitration_removeIt));
  assign when_Pipeline_l151_1 = ((! memory_arbitration_isStuck) || memory_arbitration_removeIt);
  assign when_Pipeline_l154_1 = ((! execute_arbitration_isStuck) && (! execute_arbitration_removeIt));
  assign when_Pipeline_l151_2 = ((! writeBack_arbitration_isStuck) || writeBack_arbitration_removeIt);
  assign when_Pipeline_l154_2 = ((! memory_arbitration_isStuck) && (! memory_arbitration_removeIt));
  always @(*) begin
    IBusCachedPlugin_injectionPort_ready = 1'b0;
    case(switch_Fetcher_l362)
      3'b100 : begin
        IBusCachedPlugin_injectionPort_ready = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign when_Fetcher_l378 = (! decode_arbitration_isStuck);
  assign when_CsrPlugin_l1264 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_1 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_2 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_3 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_4 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_5 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_6 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_7 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_8 = (! execute_arbitration_isStuck);
  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_2 = 32'h0;
    if(execute_CsrPlugin_csr_768) begin
      _zz_CsrPlugin_csrMapping_readDataInit_2[12 : 11] = CsrPlugin_mstatus_MPP;
      _zz_CsrPlugin_csrMapping_readDataInit_2[7 : 7] = CsrPlugin_mstatus_MPIE;
      _zz_CsrPlugin_csrMapping_readDataInit_2[3 : 3] = CsrPlugin_mstatus_MIE;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_3 = 32'h0;
    if(execute_CsrPlugin_csr_836) begin
      _zz_CsrPlugin_csrMapping_readDataInit_3[11 : 11] = CsrPlugin_mip_MEIP;
      _zz_CsrPlugin_csrMapping_readDataInit_3[7 : 7] = CsrPlugin_mip_MTIP;
      _zz_CsrPlugin_csrMapping_readDataInit_3[3 : 3] = CsrPlugin_mip_MSIP;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_4 = 32'h0;
    if(execute_CsrPlugin_csr_772) begin
      _zz_CsrPlugin_csrMapping_readDataInit_4[11 : 11] = CsrPlugin_mie_MEIE;
      _zz_CsrPlugin_csrMapping_readDataInit_4[7 : 7] = CsrPlugin_mie_MTIE;
      _zz_CsrPlugin_csrMapping_readDataInit_4[3 : 3] = CsrPlugin_mie_MSIE;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_5 = 32'h0;
    if(execute_CsrPlugin_csr_833) begin
      _zz_CsrPlugin_csrMapping_readDataInit_5[31 : 0] = CsrPlugin_mepc;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_6 = 32'h0;
    if(execute_CsrPlugin_csr_834) begin
      _zz_CsrPlugin_csrMapping_readDataInit_6[31 : 31] = CsrPlugin_mcause_interrupt;
      _zz_CsrPlugin_csrMapping_readDataInit_6[3 : 0] = CsrPlugin_mcause_exceptionCode;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_7 = 32'h0;
    if(execute_CsrPlugin_csr_835) begin
      _zz_CsrPlugin_csrMapping_readDataInit_7[31 : 0] = CsrPlugin_mtval;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_8 = 32'h0;
    if(execute_CsrPlugin_csr_3008) begin
      _zz_CsrPlugin_csrMapping_readDataInit_8[31 : 0] = _zz_CsrPlugin_csrMapping_readDataInit;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_9 = 32'h0;
    if(execute_CsrPlugin_csr_4032) begin
      _zz_CsrPlugin_csrMapping_readDataInit_9[31 : 0] = _zz_CsrPlugin_csrMapping_readDataInit_1;
    end
  end

  assign CsrPlugin_csrMapping_readDataInit = (((_zz_CsrPlugin_csrMapping_readDataInit_2 | _zz_CsrPlugin_csrMapping_readDataInit_3) | (_zz_CsrPlugin_csrMapping_readDataInit_4 | _zz_CsrPlugin_csrMapping_readDataInit_5)) | ((_zz_CsrPlugin_csrMapping_readDataInit_6 | _zz_CsrPlugin_csrMapping_readDataInit_7) | (_zz_CsrPlugin_csrMapping_readDataInit_8 | _zz_CsrPlugin_csrMapping_readDataInit_9)));
  assign when_CsrPlugin_l1297 = (CsrPlugin_privilege < execute_CsrPlugin_csrAddress[9 : 8]);
  assign when_CsrPlugin_l1302 = ((! execute_arbitration_isValid) || (! execute_IS_CSR));
  assign iBusWishbone_ADR = {_zz_iBusWishbone_ADR_1,_zz_iBusWishbone_ADR};
  assign iBusWishbone_CTI = ((_zz_iBusWishbone_ADR == 3'b111) ? 3'b111 : 3'b010);
  assign iBusWishbone_BTE = 2'b00;
  assign iBusWishbone_SEL = 4'b1111;
  assign iBusWishbone_WE = 1'b0;
  assign iBusWishbone_DAT_MOSI = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  always @(*) begin
    iBusWishbone_CYC = 1'b0;
    if(when_InstructionCache_l239) begin
      iBusWishbone_CYC = 1'b1;
    end
  end

  always @(*) begin
    iBusWishbone_STB = 1'b0;
    if(when_InstructionCache_l239) begin
      iBusWishbone_STB = 1'b1;
    end
  end

  assign when_InstructionCache_l239 = (iBus_cmd_valid || (_zz_iBusWishbone_ADR != 3'b000));
  assign iBus_cmd_ready = (iBus_cmd_valid && iBusWishbone_ACK);
  assign iBus_rsp_valid = _zz_iBus_rsp_valid;
  assign iBus_rsp_payload_data = iBusWishbone_DAT_MISO_regNext;
  assign iBus_rsp_payload_error = 1'b0;
  assign dBus_cmd_halfPipe_fire = (dBus_cmd_halfPipe_valid && dBus_cmd_halfPipe_ready);
  assign dBus_cmd_ready = (! dBus_cmd_rValid);
  assign dBus_cmd_halfPipe_valid = dBus_cmd_rValid;
  assign dBus_cmd_halfPipe_payload_wr = dBus_cmd_rData_wr;
  assign dBus_cmd_halfPipe_payload_address = dBus_cmd_rData_address;
  assign dBus_cmd_halfPipe_payload_data = dBus_cmd_rData_data;
  assign dBus_cmd_halfPipe_payload_size = dBus_cmd_rData_size;
  assign dBusWishbone_ADR = (dBus_cmd_halfPipe_payload_address >>> 2);
  assign dBusWishbone_CTI = 3'b000;
  assign dBusWishbone_BTE = 2'b00;
  always @(*) begin
    case(dBus_cmd_halfPipe_payload_size)
      2'b00 : begin
        _zz_dBusWishbone_SEL = 4'b0001;
      end
      2'b01 : begin
        _zz_dBusWishbone_SEL = 4'b0011;
      end
      default : begin
        _zz_dBusWishbone_SEL = 4'b1111;
      end
    endcase
  end

  always @(*) begin
    dBusWishbone_SEL = (_zz_dBusWishbone_SEL <<< dBus_cmd_halfPipe_payload_address[1 : 0]);
    if(when_DBusSimplePlugin_l189) begin
      dBusWishbone_SEL = 4'b1111;
    end
  end

  assign when_DBusSimplePlugin_l189 = (! dBus_cmd_halfPipe_payload_wr);
  assign dBusWishbone_WE = dBus_cmd_halfPipe_payload_wr;
  assign dBusWishbone_DAT_MOSI = dBus_cmd_halfPipe_payload_data;
  assign dBus_cmd_halfPipe_ready = (dBus_cmd_halfPipe_valid && dBusWishbone_ACK);
  assign dBusWishbone_CYC = dBus_cmd_halfPipe_valid;
  assign dBusWishbone_STB = dBus_cmd_halfPipe_valid;
  assign dBus_rsp_ready = ((dBus_cmd_halfPipe_valid && (! dBusWishbone_WE)) && dBusWishbone_ACK);
  assign dBus_rsp_data = dBusWishbone_DAT_MISO;
  assign dBus_rsp_error = 1'b0;
  always @(posedge clk) begin
    if(reset) begin
      IBusCachedPlugin_fetchPc_pcReg <= externalResetVector;
      IBusCachedPlugin_fetchPc_correctionReg <= 1'b0;
      IBusCachedPlugin_fetchPc_booted <= 1'b0;
      IBusCachedPlugin_fetchPc_inc <= 1'b0;
      _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2 <= 1'b0;
      _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_1 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_2 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_3 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_4 <= 1'b0;
      IBusCachedPlugin_rspCounter <= _zz_IBusCachedPlugin_rspCounter;
      IBusCachedPlugin_rspCounter <= 32'h0;
      _zz_2 <= 1'b1;
      execute_LightShifterPlugin_isActive <= 1'b0;
      HazardSimplePlugin_writeBackBuffer_valid <= 1'b0;
      CsrPlugin_mstatus_MIE <= 1'b0;
      CsrPlugin_mstatus_MPIE <= 1'b0;
      CsrPlugin_mstatus_MPP <= 2'b11;
      CsrPlugin_mie_MEIE <= 1'b0;
      CsrPlugin_mie_MTIE <= 1'b0;
      CsrPlugin_mie_MSIE <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= 1'b0;
      CsrPlugin_interrupt_valid <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_1 <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_2 <= 1'b0;
      CsrPlugin_hadException <= 1'b0;
      execute_CsrPlugin_wfiWake <= 1'b0;
      _zz_CsrPlugin_csrMapping_readDataInit <= 32'h0;
      execute_arbitration_isValid <= 1'b0;
      memory_arbitration_isValid <= 1'b0;
      writeBack_arbitration_isValid <= 1'b0;
      switch_Fetcher_l362 <= 3'b000;
      _zz_iBusWishbone_ADR <= 3'b000;
      _zz_iBus_rsp_valid <= 1'b0;
      dBus_cmd_rValid <= 1'b0;
    end else begin
      if(IBusCachedPlugin_fetchPc_correction) begin
        IBusCachedPlugin_fetchPc_correctionReg <= 1'b1;
      end
      if(IBusCachedPlugin_fetchPc_output_fire) begin
        IBusCachedPlugin_fetchPc_correctionReg <= 1'b0;
      end
      IBusCachedPlugin_fetchPc_booted <= 1'b1;
      if(when_Fetcher_l131) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b0;
      end
      if(IBusCachedPlugin_fetchPc_output_fire_1) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b1;
      end
      if(when_Fetcher_l131_1) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b0;
      end
      if(when_Fetcher_l158) begin
        IBusCachedPlugin_fetchPc_pcReg <= IBusCachedPlugin_fetchPc_pc;
      end
      if(IBusCachedPlugin_iBusRsp_flush) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2 <= 1'b0;
      end
      if(_zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2 <= (IBusCachedPlugin_iBusRsp_stages_0_output_valid && (! 1'b0));
      end
      if(IBusCachedPlugin_iBusRsp_flush) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= 1'b0;
      end
      if(IBusCachedPlugin_iBusRsp_stages_1_output_ready) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= (IBusCachedPlugin_iBusRsp_stages_1_output_valid && (! IBusCachedPlugin_iBusRsp_flush));
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b0;
      end
      if(when_Fetcher_l329) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b1;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= 1'b0;
      end
      if(when_Fetcher_l329_1) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= IBusCachedPlugin_injector_nextPcCalc_valids_0;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= 1'b0;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= 1'b0;
      end
      if(when_Fetcher_l329_2) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= IBusCachedPlugin_injector_nextPcCalc_valids_1;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= 1'b0;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= 1'b0;
      end
      if(when_Fetcher_l329_3) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= IBusCachedPlugin_injector_nextPcCalc_valids_2;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= 1'b0;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_4 <= 1'b0;
      end
      if(when_Fetcher_l329_4) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_4 <= IBusCachedPlugin_injector_nextPcCalc_valids_3;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_4 <= 1'b0;
      end
      if(iBus_rsp_valid) begin
        IBusCachedPlugin_rspCounter <= (IBusCachedPlugin_rspCounter + 32'h00000001);
      end

      _zz_2 <= 1'b0;
      if(when_ShiftPlugins_l169) begin
        if(when_ShiftPlugins_l175) begin
          execute_LightShifterPlugin_isActive <= 1'b1;
          if(execute_LightShifterPlugin_done) begin
            execute_LightShifterPlugin_isActive <= 1'b0;
          end
        end
      end
      if(execute_arbitration_removeIt) begin
        execute_LightShifterPlugin_isActive <= 1'b0;
      end
      HazardSimplePlugin_writeBackBuffer_valid <= HazardSimplePlugin_writeBackWrites_valid;
      if(when_CsrPlugin_l909) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= 1'b0;
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= CsrPlugin_exceptionPortCtrl_exceptionValids_decode;
      end
      if(when_CsrPlugin_l909_1) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= (CsrPlugin_exceptionPortCtrl_exceptionValids_decode && (! decode_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= CsrPlugin_exceptionPortCtrl_exceptionValids_execute;
      end
      if(when_CsrPlugin_l909_2) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= (CsrPlugin_exceptionPortCtrl_exceptionValids_execute && (! execute_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= CsrPlugin_exceptionPortCtrl_exceptionValids_memory;
      end
      if(when_CsrPlugin_l909_3) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= (CsrPlugin_exceptionPortCtrl_exceptionValids_memory && (! memory_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= 1'b0;
      end
      CsrPlugin_interrupt_valid <= 1'b0;
      if(when_CsrPlugin_l946) begin
        if(when_CsrPlugin_l952) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
        if(when_CsrPlugin_l952_1) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
        if(when_CsrPlugin_l952_2) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
      end
      if(CsrPlugin_pipelineLiberator_active) begin
        if(when_CsrPlugin_l980) begin
          CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b1;
        end
        if(when_CsrPlugin_l980_1) begin
          CsrPlugin_pipelineLiberator_pcValids_1 <= CsrPlugin_pipelineLiberator_pcValids_0;
        end
        if(when_CsrPlugin_l980_2) begin
          CsrPlugin_pipelineLiberator_pcValids_2 <= CsrPlugin_pipelineLiberator_pcValids_1;
        end
      end
      if(when_CsrPlugin_l985) begin
        CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b0;
        CsrPlugin_pipelineLiberator_pcValids_1 <= 1'b0;
        CsrPlugin_pipelineLiberator_pcValids_2 <= 1'b0;
      end
      if(CsrPlugin_interruptJump) begin
        CsrPlugin_interrupt_valid <= 1'b0;
      end
      CsrPlugin_hadException <= CsrPlugin_exception;
      if(when_CsrPlugin_l1019) begin
        case(CsrPlugin_targetPrivilege)
          2'b11 : begin
            CsrPlugin_mstatus_MIE <= 1'b0;
            CsrPlugin_mstatus_MPIE <= CsrPlugin_mstatus_MIE;
            CsrPlugin_mstatus_MPP <= CsrPlugin_privilege;
          end
          default : begin
          end
        endcase
      end
      if(when_CsrPlugin_l1064) begin
        case(switch_CsrPlugin_l1068)
          2'b11 : begin
            CsrPlugin_mstatus_MPP <= 2'b00;
            CsrPlugin_mstatus_MIE <= CsrPlugin_mstatus_MPIE;
            CsrPlugin_mstatus_MPIE <= 1'b1;
          end
          default : begin
          end
        endcase
      end
      execute_CsrPlugin_wfiWake <= (({_zz_when_CsrPlugin_l952_2,{_zz_when_CsrPlugin_l952_1,_zz_when_CsrPlugin_l952}} != 3'b000) || CsrPlugin_thirdPartyWake);
      if(when_Pipeline_l151) begin
        execute_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154) begin
        execute_arbitration_isValid <= decode_arbitration_isValid;
      end
      if(when_Pipeline_l151_1) begin
        memory_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154_1) begin
        memory_arbitration_isValid <= execute_arbitration_isValid;
      end
      if(when_Pipeline_l151_2) begin
        writeBack_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154_2) begin
        writeBack_arbitration_isValid <= memory_arbitration_isValid;
      end
      case(switch_Fetcher_l362)
        3'b000 : begin
          if(IBusCachedPlugin_injectionPort_valid) begin
            switch_Fetcher_l362 <= 3'b001;
          end
        end
        3'b001 : begin
          switch_Fetcher_l362 <= 3'b010;
        end
        3'b010 : begin
          switch_Fetcher_l362 <= 3'b011;
        end
        3'b011 : begin
          if(when_Fetcher_l378) begin
            switch_Fetcher_l362 <= 3'b100;
          end
        end
        3'b100 : begin
          switch_Fetcher_l362 <= 3'b000;
        end
        default : begin
        end
      endcase
      if(execute_CsrPlugin_csr_768) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_mstatus_MPP <= CsrPlugin_csrMapping_writeDataSignal[12 : 11];
          CsrPlugin_mstatus_MPIE <= CsrPlugin_csrMapping_writeDataSignal[7];
          CsrPlugin_mstatus_MIE <= CsrPlugin_csrMapping_writeDataSignal[3];
        end
      end
      if(execute_CsrPlugin_csr_772) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_mie_MEIE <= CsrPlugin_csrMapping_writeDataSignal[11];
          CsrPlugin_mie_MTIE <= CsrPlugin_csrMapping_writeDataSignal[7];
          CsrPlugin_mie_MSIE <= CsrPlugin_csrMapping_writeDataSignal[3];
        end
      end
      if(execute_CsrPlugin_csr_3008) begin
        if(execute_CsrPlugin_writeEnable) begin
          _zz_CsrPlugin_csrMapping_readDataInit <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
        end
      end
      if(when_InstructionCache_l239) begin
        if(iBusWishbone_ACK) begin
          _zz_iBusWishbone_ADR <= (_zz_iBusWishbone_ADR + 3'b001);
        end
      end
      _zz_iBus_rsp_valid <= (iBusWishbone_CYC && iBusWishbone_ACK);
      if(dBus_cmd_valid) begin
        dBus_cmd_rValid <= 1'b1;
      end
      if(dBus_cmd_halfPipe_fire) begin
        dBus_cmd_rValid <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(IBusCachedPlugin_iBusRsp_stages_1_output_ready) begin
      _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload <= IBusCachedPlugin_iBusRsp_stages_1_output_payload;
    end
    if(IBusCachedPlugin_iBusRsp_stages_1_input_ready) begin
      IBusCachedPlugin_s1_tightlyCoupledHit <= IBusCachedPlugin_s0_tightlyCoupledHit;
    end
    if(IBusCachedPlugin_iBusRsp_stages_2_input_ready) begin
      IBusCachedPlugin_s2_tightlyCoupledHit <= IBusCachedPlugin_s1_tightlyCoupledHit;
    end
    if(when_ShiftPlugins_l169) begin
      if(when_ShiftPlugins_l175) begin
        execute_LightShifterPlugin_amplitudeReg <= (execute_LightShifterPlugin_amplitude - 5'h01);
      end
    end
    HazardSimplePlugin_writeBackBuffer_payload_address <= HazardSimplePlugin_writeBackWrites_payload_address;
    HazardSimplePlugin_writeBackBuffer_payload_data <= HazardSimplePlugin_writeBackWrites_payload_data;
    CsrPlugin_mip_MEIP <= externalInterrupt;
    CsrPlugin_mip_MTIP <= timerInterrupt;
    CsrPlugin_mip_MSIP <= softwareInterrupt;
    CsrPlugin_mcycle <= (CsrPlugin_mcycle + 64'h0000000000000001);
    if(writeBack_arbitration_isFiring) begin
      CsrPlugin_minstret <= (CsrPlugin_minstret + 64'h0000000000000001);
    end
    if(_zz_when) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 ? IBusCachedPlugin_decodeExceptionPort_payload_code : decodeExceptionPort_payload_code);
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 ? IBusCachedPlugin_decodeExceptionPort_payload_badAddr : decodeExceptionPort_payload_badAddr);
    end
    if(CsrPlugin_selfException_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= CsrPlugin_selfException_payload_code;
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= CsrPlugin_selfException_payload_badAddr;
    end
    if(_zz_when_1) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3 ? DBusSimplePlugin_memoryExceptionPort_payload_code : BranchPlugin_branchExceptionPort_payload_code);
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3 ? DBusSimplePlugin_memoryExceptionPort_payload_badAddr : BranchPlugin_branchExceptionPort_payload_badAddr);
    end
    if(when_CsrPlugin_l946) begin
      if(when_CsrPlugin_l952) begin
        CsrPlugin_interrupt_code <= 4'b0111;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
      if(when_CsrPlugin_l952_1) begin
        CsrPlugin_interrupt_code <= 4'b0011;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
      if(when_CsrPlugin_l952_2) begin
        CsrPlugin_interrupt_code <= 4'b1011;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
    end
    if(when_CsrPlugin_l1019) begin
      case(CsrPlugin_targetPrivilege)
        2'b11 : begin
          CsrPlugin_mcause_interrupt <= (! CsrPlugin_hadException);
          CsrPlugin_mcause_exceptionCode <= CsrPlugin_trapCause;
          CsrPlugin_mepc <= writeBack_PC;
          if(CsrPlugin_hadException) begin
            CsrPlugin_mtval <= CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr;
          end
        end
        default : begin
        end
      endcase
    end
    externalInterruptArray_regNext <= externalInterruptArray;
    if(when_Pipeline_l124) begin
      decode_to_execute_PC <= decode_PC;
    end
    if(when_Pipeline_l124_1) begin
      execute_to_memory_PC <= _zz_execute_SRC2;
    end
    if(when_Pipeline_l124_2) begin
      memory_to_writeBack_PC <= memory_PC;
    end
    if(when_Pipeline_l124_3) begin
      decode_to_execute_INSTRUCTION <= decode_INSTRUCTION;
    end
    if(when_Pipeline_l124_4) begin
      execute_to_memory_INSTRUCTION <= execute_INSTRUCTION;
    end
    if(when_Pipeline_l124_5) begin
      memory_to_writeBack_INSTRUCTION <= memory_INSTRUCTION;
    end
    if(when_Pipeline_l124_6) begin
      decode_to_execute_FORMAL_PC_NEXT <= decode_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_7) begin
      execute_to_memory_FORMAL_PC_NEXT <= execute_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_8) begin
      memory_to_writeBack_FORMAL_PC_NEXT <= _zz_memory_to_writeBack_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_9) begin
      decode_to_execute_SRC1_CTRL <= _zz_decode_to_execute_SRC1_CTRL;
    end
    if(when_Pipeline_l124_10) begin
      decode_to_execute_SRC_USE_SUB_LESS <= decode_SRC_USE_SUB_LESS;
    end
    if(when_Pipeline_l124_11) begin
      decode_to_execute_MEMORY_ENABLE <= decode_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_12) begin
      execute_to_memory_MEMORY_ENABLE <= execute_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_13) begin
      memory_to_writeBack_MEMORY_ENABLE <= memory_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_14) begin
      decode_to_execute_ALU_CTRL <= _zz_decode_to_execute_ALU_CTRL;
    end
    if(when_Pipeline_l124_15) begin
      decode_to_execute_SRC2_CTRL <= _zz_decode_to_execute_SRC2_CTRL;
    end
    if(when_Pipeline_l124_16) begin
      decode_to_execute_REGFILE_WRITE_VALID <= decode_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_17) begin
      execute_to_memory_REGFILE_WRITE_VALID <= execute_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_18) begin
      memory_to_writeBack_REGFILE_WRITE_VALID <= memory_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_19) begin
      decode_to_execute_BYPASSABLE_EXECUTE_STAGE <= decode_BYPASSABLE_EXECUTE_STAGE;
    end
    if(when_Pipeline_l124_20) begin
      decode_to_execute_BYPASSABLE_MEMORY_STAGE <= decode_BYPASSABLE_MEMORY_STAGE;
    end
    if(when_Pipeline_l124_21) begin
      execute_to_memory_BYPASSABLE_MEMORY_STAGE <= execute_BYPASSABLE_MEMORY_STAGE;
    end
    if(when_Pipeline_l124_22) begin
      decode_to_execute_MEMORY_STORE <= decode_MEMORY_STORE;
    end
    if(when_Pipeline_l124_23) begin
      execute_to_memory_MEMORY_STORE <= execute_MEMORY_STORE;
    end
    if(when_Pipeline_l124_24) begin
      memory_to_writeBack_MEMORY_STORE <= memory_MEMORY_STORE;
    end
    if(when_Pipeline_l124_25) begin
      decode_to_execute_SRC_LESS_UNSIGNED <= decode_SRC_LESS_UNSIGNED;
    end
    if(when_Pipeline_l124_26) begin
      decode_to_execute_ALU_BITWISE_CTRL <= _zz_decode_to_execute_ALU_BITWISE_CTRL;
    end
    if(when_Pipeline_l124_27) begin
      decode_to_execute_SHIFT_CTRL <= _zz_decode_to_execute_SHIFT_CTRL;
    end
    if(when_Pipeline_l124_28) begin
      decode_to_execute_BRANCH_CTRL <= _zz_decode_to_execute_BRANCH_CTRL;
    end
    if(when_Pipeline_l124_29) begin
      decode_to_execute_IS_CSR <= decode_IS_CSR;
    end
    if(when_Pipeline_l124_30) begin
      decode_to_execute_ENV_CTRL <= _zz_decode_to_execute_ENV_CTRL;
    end
    if(when_Pipeline_l124_31) begin
      execute_to_memory_ENV_CTRL <= _zz_execute_to_memory_ENV_CTRL;
    end
    if(when_Pipeline_l124_32) begin
      memory_to_writeBack_ENV_CTRL <= _zz_memory_to_writeBack_ENV_CTRL;
    end
    if(when_Pipeline_l124_33) begin
      decode_to_execute_RS1 <= decode_RS1;
    end
    if(when_Pipeline_l124_34) begin
      decode_to_execute_RS2 <= decode_RS2;
    end
    if(when_Pipeline_l124_35) begin
      decode_to_execute_SRC2_FORCE_ZERO <= decode_SRC2_FORCE_ZERO;
    end
    if(when_Pipeline_l124_36) begin
      decode_to_execute_CSR_WRITE_OPCODE <= decode_CSR_WRITE_OPCODE;
    end
    if(when_Pipeline_l124_37) begin
      decode_to_execute_CSR_READ_OPCODE <= decode_CSR_READ_OPCODE;
    end
    if(when_Pipeline_l124_38) begin
      decode_to_execute_DO_EBREAK <= decode_DO_EBREAK;
    end
    if(when_Pipeline_l124_39) begin
      execute_to_memory_ALIGNEMENT_FAULT <= execute_ALIGNEMENT_FAULT;
    end
    if(when_Pipeline_l124_40) begin
      execute_to_memory_MEMORY_ADDRESS_LOW <= execute_MEMORY_ADDRESS_LOW;
    end
    if(when_Pipeline_l124_41) begin
      memory_to_writeBack_MEMORY_ADDRESS_LOW <= memory_MEMORY_ADDRESS_LOW;
    end
    if(when_Pipeline_l124_42) begin
      execute_to_memory_REGFILE_WRITE_DATA <= _zz_execute_to_memory_REGFILE_WRITE_DATA;
    end
    if(when_Pipeline_l124_43) begin
      memory_to_writeBack_REGFILE_WRITE_DATA <= memory_REGFILE_WRITE_DATA;
    end
    if(when_Pipeline_l124_44) begin
      execute_to_memory_BRANCH_DO <= execute_BRANCH_DO;
    end
    if(when_Pipeline_l124_45) begin
      execute_to_memory_BRANCH_CALC <= execute_BRANCH_CALC;
    end
    if(when_Pipeline_l124_46) begin
      memory_to_writeBack_MEMORY_READ_DATA <= memory_MEMORY_READ_DATA;
    end
    if(when_CsrPlugin_l1264) begin
      execute_CsrPlugin_csr_768 <= (decode_INSTRUCTION[31 : 20] == 12'h300);
    end
    if(when_CsrPlugin_l1264_1) begin
      execute_CsrPlugin_csr_836 <= (decode_INSTRUCTION[31 : 20] == 12'h344);
    end
    if(when_CsrPlugin_l1264_2) begin
      execute_CsrPlugin_csr_772 <= (decode_INSTRUCTION[31 : 20] == 12'h304);
    end
    if(when_CsrPlugin_l1264_3) begin
      execute_CsrPlugin_csr_773 <= (decode_INSTRUCTION[31 : 20] == 12'h305);
    end
    if(when_CsrPlugin_l1264_4) begin
      execute_CsrPlugin_csr_833 <= (decode_INSTRUCTION[31 : 20] == 12'h341);
    end
    if(when_CsrPlugin_l1264_5) begin
      execute_CsrPlugin_csr_834 <= (decode_INSTRUCTION[31 : 20] == 12'h342);
    end
    if(when_CsrPlugin_l1264_6) begin
      execute_CsrPlugin_csr_835 <= (decode_INSTRUCTION[31 : 20] == 12'h343);
    end
    if(when_CsrPlugin_l1264_7) begin
      execute_CsrPlugin_csr_3008 <= (decode_INSTRUCTION[31 : 20] == 12'hbc0);
    end
    if(when_CsrPlugin_l1264_8) begin
      execute_CsrPlugin_csr_4032 <= (decode_INSTRUCTION[31 : 20] == 12'hfc0);
    end
    if(execute_CsrPlugin_csr_836) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mip_MSIP <= CsrPlugin_csrMapping_writeDataSignal[3];
      end
    end
    if(execute_CsrPlugin_csr_773) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mtvec_base <= CsrPlugin_csrMapping_writeDataSignal[31 : 2];
        CsrPlugin_mtvec_mode <= CsrPlugin_csrMapping_writeDataSignal[1 : 0];
      end
    end
    if(execute_CsrPlugin_csr_833) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mepc <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
      end
    end
    iBusWishbone_DAT_MISO_regNext <= iBusWishbone_DAT_MISO;
    if(dBus_cmd_ready) begin
      dBus_cmd_rData_wr <= dBus_cmd_payload_wr;
      dBus_cmd_rData_address <= dBus_cmd_payload_address;
      dBus_cmd_rData_data <= dBus_cmd_payload_data;
      dBus_cmd_rData_size <= dBus_cmd_payload_size;
    end
  end

  always @(posedge clk) begin
    DebugPlugin_firstCycle <= 1'b0;
    if(debug_bus_cmd_ready) begin
      DebugPlugin_firstCycle <= 1'b1;
    end
    DebugPlugin_secondCycle <= DebugPlugin_firstCycle;
    DebugPlugin_isPipBusy <= (({writeBack_arbitration_isValid,{memory_arbitration_isValid,{execute_arbitration_isValid,decode_arbitration_isValid}}} != 4'b0000) || IBusCachedPlugin_incomingInstruction);
    if(writeBack_arbitration_isValid) begin
      DebugPlugin_busReadDataReg <= _zz_lastStageRegFileWrite_payload_data;
    end
    _zz_when_DebugPlugin_l244 <= debug_bus_cmd_payload_address[2];
    if(when_DebugPlugin_l284) begin
      DebugPlugin_busReadDataReg <= execute_PC;
    end
    DebugPlugin_resetIt_regNext <= DebugPlugin_resetIt;
  end

  always @(posedge clk) begin
    if(debugReset) begin
      DebugPlugin_resetIt <= 1'b0;
      DebugPlugin_haltIt <= 1'b0;
      DebugPlugin_stepIt <= 1'b0;
      DebugPlugin_godmode <= 1'b0;
      DebugPlugin_haltedByBreak <= 1'b0;
      DebugPlugin_debugUsed <= 1'b0;
      DebugPlugin_disableEbreak <= 1'b0;
    end else begin
      if(when_DebugPlugin_l225) begin
        DebugPlugin_godmode <= 1'b1;
      end
      if(debug_bus_cmd_valid) begin
        DebugPlugin_debugUsed <= 1'b1;
      end
      if(debug_bus_cmd_valid) begin
        case(switch_DebugPlugin_l256)
          6'h0 : begin
            if(debug_bus_cmd_payload_wr) begin
              DebugPlugin_stepIt <= debug_bus_cmd_payload_data[4];
              if(when_DebugPlugin_l260) begin
                DebugPlugin_resetIt <= 1'b1;
              end
              if(when_DebugPlugin_l260_1) begin
                DebugPlugin_resetIt <= 1'b0;
              end
              if(when_DebugPlugin_l261) begin
                DebugPlugin_haltIt <= 1'b1;
              end
              if(when_DebugPlugin_l261_1) begin
                DebugPlugin_haltIt <= 1'b0;
              end
              if(when_DebugPlugin_l262) begin
                DebugPlugin_haltedByBreak <= 1'b0;
              end
              if(when_DebugPlugin_l263) begin
                DebugPlugin_godmode <= 1'b0;
              end
              if(when_DebugPlugin_l264) begin
                DebugPlugin_disableEbreak <= 1'b1;
              end
              if(when_DebugPlugin_l264_1) begin
                DebugPlugin_disableEbreak <= 1'b0;
              end
            end
          end
          default : begin
          end
        endcase
      end
      if(when_DebugPlugin_l284) begin
        if(when_DebugPlugin_l287) begin
          DebugPlugin_haltIt <= 1'b1;
          DebugPlugin_haltedByBreak <= 1'b1;
        end
      end
      if(when_DebugPlugin_l300) begin
        if(decode_arbitration_isValid) begin
          DebugPlugin_haltIt <= 1'b1;
        end
      end
    end
  end


endmodule

module InstructionCache (
  input               io_flush,
  input               io_cpu_prefetch_isValid,
  output reg          io_cpu_prefetch_haltIt,
  input      [31:0]   io_cpu_prefetch_pc,
  input               io_cpu_fetch_isValid,
  input               io_cpu_fetch_isStuck,
  input               io_cpu_fetch_isRemoved,
  input      [31:0]   io_cpu_fetch_pc,
  output     [31:0]   io_cpu_fetch_data,
  input      [31:0]   io_cpu_fetch_mmuRsp_physicalAddress,
  input               io_cpu_fetch_mmuRsp_isIoAccess,
  input               io_cpu_fetch_mmuRsp_isPaging,
  input               io_cpu_fetch_mmuRsp_allowRead,
  input               io_cpu_fetch_mmuRsp_allowWrite,
  input               io_cpu_fetch_mmuRsp_allowExecute,
  input               io_cpu_fetch_mmuRsp_exception,
  input               io_cpu_fetch_mmuRsp_refilling,
  input               io_cpu_fetch_mmuRsp_bypassTranslation,
  output     [31:0]   io_cpu_fetch_physicalAddress,
  input               io_cpu_decode_isValid,
  input               io_cpu_decode_isStuck,
  input      [31:0]   io_cpu_decode_pc,
  output     [31:0]   io_cpu_decode_physicalAddress,
  output     [31:0]   io_cpu_decode_data,
  output              io_cpu_decode_cacheMiss,
  output              io_cpu_decode_error,
  output              io_cpu_decode_mmuRefilling,
  output              io_cpu_decode_mmuException,
  input               io_cpu_decode_isUser,
  input               io_cpu_fill_valid,
  input      [31:0]   io_cpu_fill_payload,
  output              io_mem_cmd_valid,
  input               io_mem_cmd_ready,
  output     [31:0]   io_mem_cmd_payload_address,
  output     [2:0]    io_mem_cmd_payload_size,
  input               io_mem_rsp_valid,
  input      [31:0]   io_mem_rsp_payload_data,
  input               io_mem_rsp_payload_error,
  input      [2:0]    _zz_when_Fetcher_l398,
  input      [31:0]   _zz_io_cpu_fetch_data_regNextWhen,
  input               clk,
  input               reset
);
  reg        [31:0]   _zz_banks_0_port1;
  reg        [27:0]   _zz_ways_0_tags_port1;
  wire       [27:0]   _zz_ways_0_tags_port;
  reg                 _zz_1;
  reg                 _zz_2;
  reg                 lineLoader_fire;
  reg                 lineLoader_valid;
  (* keep , syn_keep *) reg        [31:0]   lineLoader_address /* synthesis syn_keep = 1 */ ;
  reg                 lineLoader_hadError;
  reg                 lineLoader_flushPending;
  reg        [1:0]    lineLoader_flushCounter;
  wire                when_InstructionCache_l338;
  reg                 _zz_when_InstructionCache_l342;
  wire                when_InstructionCache_l342;
  wire                when_InstructionCache_l351;
  reg                 lineLoader_cmdSent;
  wire                io_mem_cmd_fire;
  wire                when_Utils_l357;
  reg                 lineLoader_wayToAllocate_willIncrement;
  wire                lineLoader_wayToAllocate_willClear;
  wire                lineLoader_wayToAllocate_willOverflowIfInc;
  wire                lineLoader_wayToAllocate_willOverflow;
  (* keep , syn_keep *) reg        [2:0]    lineLoader_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                lineLoader_write_tag_0_valid;
  wire       [0:0]    lineLoader_write_tag_0_payload_address;
  wire                lineLoader_write_tag_0_payload_data_valid;
  wire                lineLoader_write_tag_0_payload_data_error;
  wire       [25:0]   lineLoader_write_tag_0_payload_data_address;
  wire                lineLoader_write_data_0_valid;
  wire       [3:0]    lineLoader_write_data_0_payload_address;
  wire       [31:0]   lineLoader_write_data_0_payload_data;
  wire                when_InstructionCache_l401;
  wire       [3:0]    _zz_fetchStage_read_banksValue_0_dataMem;
  wire                _zz_fetchStage_read_banksValue_0_dataMem_1;
  wire       [31:0]   fetchStage_read_banksValue_0_dataMem;
  wire       [31:0]   fetchStage_read_banksValue_0_data;
  wire       [0:0]    _zz_fetchStage_read_waysValues_0_tag_valid;
  wire                _zz_fetchStage_read_waysValues_0_tag_valid_1;
  wire                fetchStage_read_waysValues_0_tag_valid;
  wire                fetchStage_read_waysValues_0_tag_error;
  wire       [25:0]   fetchStage_read_waysValues_0_tag_address;
  wire       [27:0]   _zz_fetchStage_read_waysValues_0_tag_valid_2;
  wire                fetchStage_hit_hits_0;
  wire                fetchStage_hit_valid;
  wire                fetchStage_hit_error;
  wire       [31:0]   fetchStage_hit_data;
  wire       [31:0]   fetchStage_hit_word;
  wire                when_InstructionCache_l435;
  reg        [31:0]   io_cpu_fetch_data_regNextWhen;
  wire                when_InstructionCache_l459;
  reg        [31:0]   decodeStage_mmuRsp_physicalAddress;
  reg                 decodeStage_mmuRsp_isIoAccess;
  reg                 decodeStage_mmuRsp_isPaging;
  reg                 decodeStage_mmuRsp_allowRead;
  reg                 decodeStage_mmuRsp_allowWrite;
  reg                 decodeStage_mmuRsp_allowExecute;
  reg                 decodeStage_mmuRsp_exception;
  reg                 decodeStage_mmuRsp_refilling;
  reg                 decodeStage_mmuRsp_bypassTranslation;
  wire                when_InstructionCache_l459_1;
  reg                 decodeStage_hit_valid;
  wire                when_InstructionCache_l459_2;
  reg                 decodeStage_hit_error;
  wire                when_Fetcher_l398;
  (* ram_style = "block" *) reg [31:0] banks_0 [0:15];
  (* ram_style = "block" *) reg [27:0] ways_0_tags [0:1];

  assign _zz_ways_0_tags_port = {lineLoader_write_tag_0_payload_data_address,{lineLoader_write_tag_0_payload_data_error,lineLoader_write_tag_0_payload_data_valid}};
  always @(posedge clk) begin
    if(_zz_1) begin
      banks_0[lineLoader_write_data_0_payload_address] <= lineLoader_write_data_0_payload_data;
    end
  end

  always @(posedge clk) begin
    if(_zz_fetchStage_read_banksValue_0_dataMem_1) begin
      _zz_banks_0_port1 <= banks_0[_zz_fetchStage_read_banksValue_0_dataMem];
    end
  end

  always @(posedge clk) begin
    if(_zz_2) begin
      ways_0_tags[lineLoader_write_tag_0_payload_address] <= _zz_ways_0_tags_port;
    end
  end

  always @(posedge clk) begin
    if(_zz_fetchStage_read_waysValues_0_tag_valid_1) begin
      _zz_ways_0_tags_port1 <= ways_0_tags[_zz_fetchStage_read_waysValues_0_tag_valid];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(lineLoader_write_data_0_valid) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(lineLoader_write_tag_0_valid) begin
      _zz_2 = 1'b1;
    end
  end

  always @(*) begin
    lineLoader_fire = 1'b0;
    if(io_mem_rsp_valid) begin
      if(when_InstructionCache_l401) begin
        lineLoader_fire = 1'b1;
      end
    end
  end

  always @(*) begin
    io_cpu_prefetch_haltIt = (lineLoader_valid || lineLoader_flushPending);
    if(when_InstructionCache_l338) begin
      io_cpu_prefetch_haltIt = 1'b1;
    end
    if(when_InstructionCache_l342) begin
      io_cpu_prefetch_haltIt = 1'b1;
    end
    if(io_flush) begin
      io_cpu_prefetch_haltIt = 1'b1;
    end
  end

  assign when_InstructionCache_l338 = (! lineLoader_flushCounter[1]);
  assign when_InstructionCache_l342 = (! _zz_when_InstructionCache_l342);
  assign when_InstructionCache_l351 = (lineLoader_flushPending && (! (lineLoader_valid || io_cpu_fetch_isValid)));
  assign io_mem_cmd_fire = (io_mem_cmd_valid && io_mem_cmd_ready);
  assign io_mem_cmd_valid = (lineLoader_valid && (! lineLoader_cmdSent));
  assign io_mem_cmd_payload_address = {lineLoader_address[31 : 5],5'h0};
  assign io_mem_cmd_payload_size = 3'b101;
  assign when_Utils_l357 = (! lineLoader_valid);
  always @(*) begin
    lineLoader_wayToAllocate_willIncrement = 1'b0;
    if(when_Utils_l357) begin
      lineLoader_wayToAllocate_willIncrement = 1'b1;
    end
  end

  assign lineLoader_wayToAllocate_willClear = 1'b0;
  assign lineLoader_wayToAllocate_willOverflowIfInc = 1'b1;
  assign lineLoader_wayToAllocate_willOverflow = (lineLoader_wayToAllocate_willOverflowIfInc && lineLoader_wayToAllocate_willIncrement);
  assign lineLoader_write_tag_0_valid = ((1'b1 && lineLoader_fire) || (! lineLoader_flushCounter[1]));
  assign lineLoader_write_tag_0_payload_address = (lineLoader_flushCounter[1] ? lineLoader_address[5 : 5] : lineLoader_flushCounter[0 : 0]);
  assign lineLoader_write_tag_0_payload_data_valid = lineLoader_flushCounter[1];
  assign lineLoader_write_tag_0_payload_data_error = (lineLoader_hadError || io_mem_rsp_payload_error);
  assign lineLoader_write_tag_0_payload_data_address = lineLoader_address[31 : 6];
  assign lineLoader_write_data_0_valid = (io_mem_rsp_valid && 1'b1);
  assign lineLoader_write_data_0_payload_address = {lineLoader_address[5 : 5],lineLoader_wordIndex};
  assign lineLoader_write_data_0_payload_data = io_mem_rsp_payload_data;
  assign when_InstructionCache_l401 = (lineLoader_wordIndex == 3'b111);
  assign _zz_fetchStage_read_banksValue_0_dataMem = io_cpu_prefetch_pc[5 : 2];
  assign _zz_fetchStage_read_banksValue_0_dataMem_1 = (! io_cpu_fetch_isStuck);
  assign fetchStage_read_banksValue_0_dataMem = _zz_banks_0_port1;
  assign fetchStage_read_banksValue_0_data = fetchStage_read_banksValue_0_dataMem[31 : 0];
  assign _zz_fetchStage_read_waysValues_0_tag_valid = io_cpu_prefetch_pc[5 : 5];
  assign _zz_fetchStage_read_waysValues_0_tag_valid_1 = (! io_cpu_fetch_isStuck);
  assign _zz_fetchStage_read_waysValues_0_tag_valid_2 = _zz_ways_0_tags_port1;
  assign fetchStage_read_waysValues_0_tag_valid = _zz_fetchStage_read_waysValues_0_tag_valid_2[0];
  assign fetchStage_read_waysValues_0_tag_error = _zz_fetchStage_read_waysValues_0_tag_valid_2[1];
  assign fetchStage_read_waysValues_0_tag_address = _zz_fetchStage_read_waysValues_0_tag_valid_2[27 : 2];
  assign fetchStage_hit_hits_0 = (fetchStage_read_waysValues_0_tag_valid && (fetchStage_read_waysValues_0_tag_address == io_cpu_fetch_mmuRsp_physicalAddress[31 : 6]));
  assign fetchStage_hit_valid = (fetchStage_hit_hits_0 != 1'b0);
  assign fetchStage_hit_error = fetchStage_read_waysValues_0_tag_error;
  assign fetchStage_hit_data = fetchStage_read_banksValue_0_data;
  assign fetchStage_hit_word = fetchStage_hit_data;
  assign io_cpu_fetch_data = fetchStage_hit_word;
  assign when_InstructionCache_l435 = (! io_cpu_decode_isStuck);
  assign io_cpu_decode_data = io_cpu_fetch_data_regNextWhen;
  assign io_cpu_fetch_physicalAddress = io_cpu_fetch_mmuRsp_physicalAddress;
  assign when_InstructionCache_l459 = (! io_cpu_decode_isStuck);
  assign when_InstructionCache_l459_1 = (! io_cpu_decode_isStuck);
  assign when_InstructionCache_l459_2 = (! io_cpu_decode_isStuck);
  assign io_cpu_decode_cacheMiss = (! decodeStage_hit_valid);
  assign io_cpu_decode_error = (decodeStage_hit_error || ((! decodeStage_mmuRsp_isPaging) && (decodeStage_mmuRsp_exception || (! decodeStage_mmuRsp_allowExecute))));
  assign io_cpu_decode_mmuRefilling = decodeStage_mmuRsp_refilling;
  assign io_cpu_decode_mmuException = (((! decodeStage_mmuRsp_refilling) && decodeStage_mmuRsp_isPaging) && (decodeStage_mmuRsp_exception || (! decodeStage_mmuRsp_allowExecute)));
  assign io_cpu_decode_physicalAddress = decodeStage_mmuRsp_physicalAddress;
  assign when_Fetcher_l398 = (_zz_when_Fetcher_l398 != 3'b000);
  always @(posedge clk) begin
    if(reset) begin
      lineLoader_valid <= 1'b0;
      lineLoader_hadError <= 1'b0;
      lineLoader_flushPending <= 1'b1;
      lineLoader_cmdSent <= 1'b0;
      lineLoader_wordIndex <= 3'b000;
    end else begin
      if(lineLoader_fire) begin
        lineLoader_valid <= 1'b0;
      end
      if(lineLoader_fire) begin
        lineLoader_hadError <= 1'b0;
      end
      if(io_cpu_fill_valid) begin
        lineLoader_valid <= 1'b1;
      end
      if(io_flush) begin
        lineLoader_flushPending <= 1'b1;
      end
      if(when_InstructionCache_l351) begin
        lineLoader_flushPending <= 1'b0;
      end
      if(io_mem_cmd_fire) begin
        lineLoader_cmdSent <= 1'b1;
      end
      if(lineLoader_fire) begin
        lineLoader_cmdSent <= 1'b0;
      end
      if(io_mem_rsp_valid) begin
        lineLoader_wordIndex <= (lineLoader_wordIndex + 3'b001);
        if(io_mem_rsp_payload_error) begin
          lineLoader_hadError <= 1'b1;
        end
      end
    end
  end

  always @(posedge clk) begin
    if(io_cpu_fill_valid) begin
      lineLoader_address <= io_cpu_fill_payload;
    end
    if(when_InstructionCache_l338) begin
      lineLoader_flushCounter <= (lineLoader_flushCounter + 2'b01);
    end
    _zz_when_InstructionCache_l342 <= lineLoader_flushCounter[1];
    if(when_InstructionCache_l351) begin
      lineLoader_flushCounter <= 2'b00;
    end
    if(when_InstructionCache_l435) begin
      io_cpu_fetch_data_regNextWhen <= io_cpu_fetch_data;
    end
    if(when_InstructionCache_l459) begin
      decodeStage_mmuRsp_physicalAddress <= io_cpu_fetch_mmuRsp_physicalAddress;
      decodeStage_mmuRsp_isIoAccess <= io_cpu_fetch_mmuRsp_isIoAccess;
      decodeStage_mmuRsp_isPaging <= io_cpu_fetch_mmuRsp_isPaging;
      decodeStage_mmuRsp_allowRead <= io_cpu_fetch_mmuRsp_allowRead;
      decodeStage_mmuRsp_allowWrite <= io_cpu_fetch_mmuRsp_allowWrite;
      decodeStage_mmuRsp_allowExecute <= io_cpu_fetch_mmuRsp_allowExecute;
      decodeStage_mmuRsp_exception <= io_cpu_fetch_mmuRsp_exception;
      decodeStage_mmuRsp_refilling <= io_cpu_fetch_mmuRsp_refilling;
      decodeStage_mmuRsp_bypassTranslation <= io_cpu_fetch_mmuRsp_bypassTranslation;
    end
    if(when_InstructionCache_l459_1) begin
      decodeStage_hit_valid <= fetchStage_hit_valid;
    end
    if(when_InstructionCache_l459_2) begin
      decodeStage_hit_error <= fetchStage_hit_error;
    end
    if(when_Fetcher_l398) begin
      io_cpu_fetch_data_regNextWhen <= _zz_io_cpu_fetch_data_regNextWhen;
    end
  end


endmodule
//////////////////////////////////////////////////////////////////////////////////
// Author : Tony Ho
//
// Create Date: 11/17/2023
// Design Name:
// Module Name: FSIC
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module FSIC #( 
    parameter BITS=32,
    parameter pUSER_PROJECT_SIDEBAND_WIDTH   = 5,
      parameter pSERIALIO_WIDTH   = 13,
  
    parameter pADDR_WIDTH   = 15,
    parameter pDATA_WIDTH   = 32,
    parameter pRxFIFO_DEPTH = 5,
    parameter pCLK_RATIO =4
  ) (
  input  wire          vccd,
  input  wire          vssd,
  input  wire          wb_rst,
  input  wire          wb_clk,
  input  wire  [31: 0] wbs_adr,
  input  wire  [31: 0] wbs_wdata,
  input  wire   [3: 0] wbs_sel,
  input  wire          wbs_cyc,
  input  wire          wbs_stb,
  input  wire          wbs_we,
  input  wire  [37: 0] io_in,
  output wire          wbs_ack,
  output wire  [31: 0] wbs_rdata,
  output wire   [2: 0] user_irq,
  output wire  [37: 0] io_out,
  output wire  [37: 0] io_oeb,
  input  wire          user_clock2
);


wire           m_awvalid_aa_cfg_awvalid;
wire   [31: 0] m_awaddr_aa_cfg_awaddr;
wire           m_wvalid_aa_cfg_wvalid;
wire   [31: 0] m_wdata_aa_cfg_wdata;
wire    [3: 0] m_wstrb_aa_cfg_wstrb;
wire           m_arvalid_aa_cfg_arvalid;
wire   [31: 0] m_araddr_aa_cfg_araddr;
wire           m_rready_aa_cfg_rready;
wire           s_wready_axi_wready1;
wire           s_awready_axi_awready1;
wire           s_arready_axi_arready1;
wire   [31: 0] s_rdata_axi_rdata1;
wire           s_rvalid_axi_rvalid1;
wire           axi_awready_axi_awready4;
wire           axi_wready_axi_wready4;
wire           axi_arready_axi_arready4;
wire   [31: 0] axi_rdata_axi_rdata4;
wire           axi_rvalid_axi_rvalid4;
wire           axi_awready_axi_awready3;
wire           axi_wready_axi_wready3;
wire           axi_arready_axi_arready3;
wire   [31: 0] axi_rdata_axi_rdata3;
wire           axi_rvalid_axi_rvalid3;
wire           axi_awready_axi_awready0;
wire           axi_wready_axi_wready0;
wire           axi_arready_axi_arready0;
wire   [31: 0] axi_rdata_axi_rdata0;
wire           axi_rvalid_axi_rvalid0;
wire           axi_awready_axi_awready2;
wire           axi_wready_axi_wready2;
wire           axi_arready_axi_arready2;
wire   [31: 0] axi_rdata_axi_rdata2;
wire           axi_rvalid_axi_rvalid2;
wire           axi_awvalid_s_awvalid;
wire   [14: 0] axi_awaddr_s_awaddr;
wire           axi_wvalid_s_wvalid;
wire   [31: 0] axi_wdata_s_wdata;
wire    [3: 0] axi_wstrb_s_wstrb;
wire           axi_arvalid_s_arvalid;
wire   [14: 0] axi_araddr_s_araddr;
wire           axi_rready_s_rready;
wire   [31: 0] aa_cfg_rdata_m_rdata;
wire           aa_cfg_rvalid_m_rvalid;
wire           aa_cfg_awready_m_awready;
wire           aa_cfg_wready_m_wready;
wire           aa_cfg_arready_m_arready;
wire           cc_aa_enable;
wire   [31: 0] as_aa_tdata;
wire    [3: 0] as_aa_tstrb;
wire    [3: 0] as_aa_tkeep;
wire           as_aa_tlast;
wire           as_aa_tvalid;
wire    [1: 0] as_aa_tuser;
wire           as_aa_tready;
//wire           axi_awvalid;
//wire   [14: 0] axi_awaddr;
//wire           axi_wvalid;
//wire   [31: 0] axi_wdata;
//wire    [3: 0] axi_wstrb;
//wire           axi_arvalid;
//wire   [14: 0] axi_araddr;
//wire           axi_rready;
wire           cc_as_enable;
wire   [31: 0] aa_as_tdata;
wire    [3: 0] aa_as_tstrb;
wire    [3: 0] aa_as_tkeep;
wire           aa_as_tlast;
wire           aa_as_tvalid;
wire    [1: 0] aa_as_tuser;
wire           aa_as_tready;
wire   [31: 0] is_as_tdata;
wire    [3: 0] is_as_tstrb;
wire    [3: 0] is_as_tkeep;
wire           is_as_tlast;
wire    [1: 0] is_as_tid;
wire           is_as_tvalid;
wire    [1: 0] is_as_tuser;
wire           is_as_tready;

  wire   [pUSER_PROJECT_SIDEBAND_WIDTH-1:0] is_as_tupsb;

wire   [31: 0] m_tdata_la_as_tdata;
wire    [3: 0] m_tstrb_la_as_tstrb;
wire    [3: 0] m_tkeep_la_as_tkeep;
wire           m_tlast_la_as_tlast;
wire           m_tvalid_la_as_tvalid;
wire    [1: 0] m_tuser_la_as_tuser;
wire           la_hpri_req;
wire   [31: 0] m_tdata_up_as_tdata;

  wire   [pUSER_PROJECT_SIDEBAND_WIDTH-1:0] m_tupsb_up_as_tupsb;

wire    [3: 0] m_tstrb_up_as_tstrb;
wire    [3: 0] m_tkeep_up_as_tkeep;
wire           m_tlast_up_as_tlast;
wire           m_tvalid_up_as_tvalid;
wire    [1: 0] m_tuser_up_as_tuser;
wire           s_tready_up_as_tready;
wire           high_pri_irq_up_hpri_req;
wire           cc_is_enable;
wire   [31: 0] as_is_tdata;
wire    [3: 0] as_is_tstrb;
wire    [3: 0] as_is_tkeep;
wire           as_is_tlast;
wire    [1: 0] as_is_tid;
wire           as_is_tvalid;
wire    [1: 0] as_is_tuser;
wire           as_is_tready;

  wire   [pUSER_PROJECT_SIDEBAND_WIDTH-1:0] as_is_tupsb;

wire           ioclk;
wire   [pSERIALIO_WIDTH-1: 0] serial_rxd;
wire           serial_rclk;
wire           cc_la_enable;
wire           as_la_tready_m_tready;
wire   [23: 0] up_la_data;
wire           cc_up_enable;
wire    [4: 0] user_prj_sel;
wire   [31: 0] as_up_tdata_s_tdata;

  wire   [pUSER_PROJECT_SIDEBAND_WIDTH-1:0] as_up_tupsb_s_tupsb;

wire    [3: 0] as_up_tstrb_s_tstrb;
wire    [3: 0] as_up_tkeep_s_tkeep;
wire           as_up_tlast_s_tlast;
wire           as_up_tvalid_s_tvalid;
wire    [1: 0] as_up_tuser_s_tuser;
wire           as_up_tready_m_tready;
wire           mb_irq;
wire           low__pri_irq;
wire           high_pri_irq;
wire           io_clk;
wire   [pSERIALIO_WIDTH-1: 0] serial_txd;
wire           serial_tclk;
wire           axi_clk;
wire           axi_reset_n;
wire           axis_clk;
wire           uck2_rst_n;
wire           axis_rst_n;


// This code snippet was auto generated by xls2vlog.py from source file: /home/josh/Downloads/Interface-Definition.xlsx
// User: josh
// Date: Sep-22-23



CFG_CTRL #(.pADDR_WIDTH( pADDR_WIDTH ),
           .pDATA_WIDTH( 32 )) U_CFG_CTRL0 (
                                            .aa_cfg_awvalid (m_awvalid_aa_cfg_awvalid),// I  
                                            .aa_cfg_awaddr  (m_awaddr_aa_cfg_awaddr),  // I  32
                                            .aa_cfg_wvalid  (m_wvalid_aa_cfg_wvalid),  // I  
                                            .aa_cfg_wdata   (m_wdata_aa_cfg_wdata),    // I  32
                                            .aa_cfg_wstrb   (m_wstrb_aa_cfg_wstrb),    // I  4
                                            .aa_cfg_arvalid (m_arvalid_aa_cfg_arvalid),// I  
                                            .aa_cfg_araddr  (m_araddr_aa_cfg_araddr),  // I  32
                                            .aa_cfg_rready  (m_rready_aa_cfg_rready),  // I  
                                            .axi_wready1    (s_wready_axi_wready1),    // I  
                                            .axi_awready1   (s_awready_axi_awready1),  // I  
                                            .axi_arready1   (s_arready_axi_arready1),  // I  
                                            .axi_rdata1     (s_rdata_axi_rdata1),      // I  32
                                            .axi_rvalid1    (s_rvalid_axi_rvalid1),    // I  
                                            .axi_awready4   (axi_awready_axi_awready4),// I  
                                            .axi_wready4    (axi_wready_axi_wready4),  // I  
                                            .axi_arready4   (axi_arready_axi_arready4),// I  
                                            .axi_rdata4     (axi_rdata_axi_rdata4),    // I  32
                                            .axi_rvalid4    (axi_rvalid_axi_rvalid4),  // I  
                                            .axi_awready3   (axi_awready_axi_awready3),// I  
                                            .axi_wready3    (axi_wready_axi_wready3),  // I  
                                            .axi_arready3   (axi_arready_axi_arready3),// I  
                                            .axi_rdata3     (axi_rdata_axi_rdata3),    // I  32
                                            .axi_rvalid3    (axi_rvalid_axi_rvalid3),  // I  
                                            .axi_awready0   (axi_awready_axi_awready0),// I  
                                            .axi_wready0    (axi_wready_axi_wready0),  // I  
                                            .axi_arready0   (axi_arready_axi_arready0),// I  
                                            .axi_rdata0     (axi_rdata_axi_rdata0),    // I  32
                                            .axi_rvalid0    (axi_rvalid_axi_rvalid0),  // I  
                                            .axi_awready2   (axi_awready_axi_awready2),// I  
                                            .axi_wready2    (axi_wready_axi_wready2),  // I  
                                            .axi_arready2   (axi_arready_axi_arready2),// I  
                                            .axi_rdata2     (axi_rdata_axi_rdata2),    // I  32
                                            .axi_rvalid2    (axi_rvalid_axi_rvalid2),  // I  
                                            .axi_awvalid    (axi_awvalid_s_awvalid),   // O  
                                            .axi_awaddr     (axi_awaddr_s_awaddr),     // O  15
                                            .axi_wvalid     (axi_wvalid_s_wvalid),     // O  
                                            .axi_wdata      (axi_wdata_s_wdata),       // O  32
                                            .axi_wstrb      (axi_wstrb_s_wstrb),       // O  4
                                            .axi_arvalid    (axi_arvalid_s_arvalid),   // O  
                                            .axi_araddr     (axi_araddr_s_araddr),     // O  15
                                            .axi_rready     (axi_rready_s_rready),     // O  
                                            .aa_cfg_rdata   (aa_cfg_rdata_m_rdata),    // O  32
                                            .aa_cfg_rvalid  (aa_cfg_rvalid_m_rvalid),  // O  
                                            .aa_cfg_awready (aa_cfg_awready_m_awready),// O  
                                            .aa_cfg_wready  (aa_cfg_wready_m_wready),  // O  
                                            .aa_cfg_arready (aa_cfg_arready_m_arready),// O  
                                            .cc_aa_enable   (cc_aa_enable),            // O  
                                            .cc_as_enable   (cc_as_enable),            // O  
                                            .cc_is_enable   (cc_is_enable),            // O  
                                            .cc_la_enable   (cc_la_enable),            // O  
                                            .cc_up_enable   (cc_up_enable),            // O  
                                            .user_prj_sel   (user_prj_sel),            // O  5
                                            .wb_rst         (wb_rst),                  // I  
                                            .wb_clk         (wb_clk),                  // I  
                                            .wbs_adr        (wbs_adr),                 // I  32
                                            .wbs_wdata      (wbs_wdata),               // I  32
                                            .wbs_sel        (wbs_sel),                 // I  4
                                            .wbs_cyc        (wbs_cyc),                 // I  
                                            .wbs_stb        (wbs_stb),                 // I  
                                            .wbs_we         (wbs_we),                  // I  
                                            .wbs_ack        (wbs_ack),                 // O  
                                            .wbs_rdata      (wbs_rdata),               // O  32
                                            .user_clock2    (user_clock2),             // I  
                                            .axi_clk        (axi_clk),                 // I  
                                            .axi_reset_n    (axi_reset_n),             // I  
                                            .uck2_rst_n     (uck2_rst_n)               // I  
                                           );


// This code snippet was auto generated by xls2vlog.py from source file: /home/josh/Downloads/Interface-Definition.xlsx
// User: josh
// Date: Sep-22-23



AXIL_AXIS #(.pADDR_WIDTH( pADDR_WIDTH ),
            .pDATA_WIDTH( 32 )) U_AXIL_AXIS0 (
                                              .m_awvalid    (m_awvalid_aa_cfg_awvalid),// O  
                                              .m_awaddr     (m_awaddr_aa_cfg_awaddr),  // O  32
                                              .m_wvalid     (m_wvalid_aa_cfg_wvalid),  // O  
                                              .m_wdata      (m_wdata_aa_cfg_wdata),    // O  32
                                              .m_wstrb      (m_wstrb_aa_cfg_wstrb),    // O  4
                                              .m_arvalid    (m_arvalid_aa_cfg_arvalid),// O  
                                              .m_araddr     (m_araddr_aa_cfg_araddr),  // O  32
                                              .m_rready     (m_rready_aa_cfg_rready),  // O  
                                              .s_wready     (s_wready_axi_wready1),    // O  
                                              .s_awready    (s_awready_axi_awready1),  // O  
                                              .s_arready    (s_arready_axi_arready1),  // O  
                                              .s_rdata      (s_rdata_axi_rdata1),      // O  32
                                              .s_rvalid     (s_rvalid_axi_rvalid1),    // O  
                                              .s_awvalid    (axi_awvalid_s_awvalid),   // I  
                                              .s_awaddr     (axi_awaddr_s_awaddr),     // I  15
                                              .s_wvalid     (axi_wvalid_s_wvalid),     // I  
                                              .s_wdata      (axi_wdata_s_wdata),       // I  32
                                              .s_wstrb      (axi_wstrb_s_wstrb),       // I  4
                                              .s_arvalid    (axi_arvalid_s_arvalid),   // I  
                                              .s_araddr     (axi_araddr_s_araddr),     // I  15
                                              .s_rready     (axi_rready_s_rready),     // I  
                                              .m_rdata      (aa_cfg_rdata_m_rdata),    // I  32
                                              .m_rvalid     (aa_cfg_rvalid_m_rvalid),  // I  
                                              .m_awready    (aa_cfg_awready_m_awready),// I  
                                              .m_wready     (aa_cfg_wready_m_wready),  // I  
                                              .m_arready    (aa_cfg_arready_m_arready),// I  
                                              .cc_aa_enable (cc_aa_enable),            // I  
                                              .as_aa_tdata  (as_aa_tdata),             // I  32
                                              .as_aa_tstrb  (as_aa_tstrb),             // I  4
                                              .as_aa_tkeep  (as_aa_tkeep),             // I  4
                                              .as_aa_tlast  (as_aa_tlast),             // I  
                                              .as_aa_tvalid (as_aa_tvalid),            // I  
                                              .as_aa_tuser  (as_aa_tuser),             // I  2
                                              .as_aa_tready (as_aa_tready),            // I  
                                              .aa_as_tdata  (aa_as_tdata),             // O  32
                                              .aa_as_tstrb  (aa_as_tstrb),             // O  4
                                              .aa_as_tkeep  (aa_as_tkeep),             // O  4
                                              .aa_as_tlast  (aa_as_tlast),             // O  
                                              .aa_as_tvalid (aa_as_tvalid),            // O  
                                              .aa_as_tuser  (aa_as_tuser),             // O  2
                                              .aa_as_tready (aa_as_tready),            // O  
                                              .mb_irq       (mb_irq),                  // O  
                                              .axi_clk      (axi_clk),                 // I  
                                              .axi_reset_n  (axi_reset_n),             // I  
                                              .axis_clk     (axis_clk),                // I  
                                              .axis_rst_n   (axis_rst_n)               // I  
                                             );


// This code snippet was auto generated by xls2vlog.py from source file: /home/josh/Downloads/Interface-Definition.xlsx
// User: josh
// Date: Sep-22-23



AXIS_SW #(  .pUSER_PROJECT_SIDEBAND_WIDTH( pUSER_PROJECT_SIDEBAND_WIDTH ),
      .pADDR_WIDTH( pADDR_WIDTH ),
      .pDATA_WIDTH( 32 )) AXIS_SW0 (
                                        .axi_awready  (axi_awready_axi_awready4),// O  
                                        .axi_wready   (axi_wready_axi_wready4),  // O  
                                        .axi_arready  (axi_arready_axi_arready4),// O  
                                        .axi_rdata    (axi_rdata_axi_rdata4),    // O  32
                                        .axi_rvalid   (axi_rvalid_axi_rvalid4),  // O  
                                        .as_aa_tdata  (as_aa_tdata),             // O  32
                                        .as_aa_tstrb  (as_aa_tstrb),             // O  4
                                        .as_aa_tkeep  (as_aa_tkeep),             // O  4
                                        .as_aa_tlast  (as_aa_tlast),             // O  
                                        .as_aa_tvalid (as_aa_tvalid),            // O  
                                        .as_aa_tuser  (as_aa_tuser),             // O  2
                                        .as_aa_tready (as_aa_tready),            // O  
                                        .axi_awvalid  (axi_awvalid_s_awvalid),   // I  
                                        .axi_awaddr   (axi_awaddr_s_awaddr),     // I  15
                                        .axi_wvalid   (axi_wvalid_s_wvalid),     // I  
                                        .axi_wdata    (axi_wdata_s_wdata),       // I  32
                                        .axi_wstrb    (axi_wstrb_s_wstrb),       // I  4
                                        .axi_arvalid  (axi_arvalid_s_arvalid),   // I  
                                        .axi_araddr   (axi_araddr_s_araddr),     // I  15
                                        .axi_rready   (axi_rready_s_rready),     // I  
                                        .cc_as_enable (cc_as_enable),            // I  
                                        .aa_as_tdata  (aa_as_tdata),             // I  32
                                        .aa_as_tstrb  (aa_as_tstrb),             // I  4
                                        .aa_as_tkeep  (aa_as_tkeep),             // I  4
                                        .aa_as_tlast  (aa_as_tlast),             // I  
                                        .aa_as_tvalid (aa_as_tvalid),            // I  
                                        .aa_as_tuser  (aa_as_tuser),             // I  2
                                        .aa_as_tready (aa_as_tready),            // I  
                                        .is_as_tdata  (is_as_tdata),             // I  32

                      .is_as_tupsb  (is_as_tupsb),     // I  5

                                        .is_as_tstrb  (is_as_tstrb),             // I  4
                                        .is_as_tkeep  (is_as_tkeep),             // I  4
                                        .is_as_tlast  (is_as_tlast),             // I  
                                        .is_as_tid    (is_as_tid),               // I  2
                                        .is_as_tvalid (is_as_tvalid),            // I  
                                        .is_as_tuser  (is_as_tuser),             // I  2
                                        .is_as_tready (is_as_tready),            // I  
                                        .la_as_tdata  (m_tdata_la_as_tdata),     // I  32
                                        .la_as_tstrb  (m_tstrb_la_as_tstrb),     // I  4
                                        .la_as_tkeep  (m_tkeep_la_as_tkeep),     // I  4
                                        .la_as_tlast  (m_tlast_la_as_tlast),     // I  
                                        .la_as_tvalid (m_tvalid_la_as_tvalid),   // I  
                                        .la_as_tuser  (m_tuser_la_as_tuser),     // I  2
                                        .la_hpri_req  (la_hpri_req),             // I  
                                        .up_as_tdata  (m_tdata_up_as_tdata),     // I  32

                      .up_as_tupsb  (m_tupsb_up_as_tupsb),     // I  5

                                        .up_as_tstrb  (m_tstrb_up_as_tstrb),     // I  4
                                        .up_as_tkeep  (m_tkeep_up_as_tkeep),     // I  4
                                        .up_as_tlast  (m_tlast_up_as_tlast),     // I  
                                        .up_as_tvalid (m_tvalid_up_as_tvalid),   // I  
                                        .up_as_tuser  (m_tuser_up_as_tuser),     // I  2
                                        .up_as_tready (s_tready_up_as_tready),   // I  
                                        .up_hpri_req  (high_pri_irq_up_hpri_req),// I  
                                        .as_is_tdata  (as_is_tdata),             // O  32

                      .as_is_tupsb  (as_is_tupsb),     // O  5

                                        .as_is_tstrb  (as_is_tstrb),             // O  4
                                        .as_is_tkeep  (as_is_tkeep),             // O  4
                                        .as_is_tlast  (as_is_tlast),             // O  
                                        .as_is_tid    (as_is_tid),               // O  2
                                        .as_is_tvalid (as_is_tvalid),            // O  
                                        .as_is_tuser  (as_is_tuser),             // O  2
                                        .as_is_tready (as_is_tready),            // O  
                                        .as_la_tready (as_la_tready_m_tready),   // O  
                                        .as_up_tdata  (as_up_tdata_s_tdata),     // O  32

                      .as_up_tupsb  (as_up_tupsb_s_tupsb),     // O  5

                                        .as_up_tstrb  (as_up_tstrb_s_tstrb),     // O  4
                                        .as_up_tkeep  (as_up_tkeep_s_tkeep),     // O  4
                                        .as_up_tlast  (as_up_tlast_s_tlast),     // O  
                                        .as_up_tvalid (as_up_tvalid_s_tvalid),   // O  
                                        .as_up_tuser  (as_up_tuser_s_tuser),     // O  2
                                        .as_up_tready (as_up_tready_m_tready),   // O  
                                        .axi_reset_n  (axi_reset_n),             // I  
                                        .axis_clk     (axis_clk),                // I  
                                        .axis_rst_n   (axis_rst_n)               // I  
                                       );


// This code snippet was auto generated by xls2vlog.py from source file: /home/josh/Downloads/Interface-Definition.xlsx
// User: josh
// Date: Sep-22-23



IO_SERDES #(.pUSER_PROJECT_SIDEBAND_WIDTH( pUSER_PROJECT_SIDEBAND_WIDTH ),
      .pSERIALIO_WIDTH( pSERIALIO_WIDTH ),
            .pADDR_WIDTH( pADDR_WIDTH ),
            .pDATA_WIDTH( pDATA_WIDTH ),
            .pRxFIFO_DEPTH( pRxFIFO_DEPTH ),
            .pCLK_RATIO      ( pCLK_RATIO)) U_IO_SERDES0 (
                                                  .axi_awready  (axi_awready_axi_awready3),// O  
                                                  .axi_wready   (axi_wready_axi_wready3),  // O  
                                                  .axi_arready  (axi_arready_axi_arready3),// O  
                                                  .axi_rdata    (axi_rdata_axi_rdata3),    // O  32
                                                  .axi_rvalid   (axi_rvalid_axi_rvalid3),  // O  
                                                  .is_as_tdata  (is_as_tdata),             // O  32

                           .is_as_tupsb  (is_as_tupsb),     // O  5

                          .is_as_tstrb  (is_as_tstrb),             // O  4
                                                  .is_as_tkeep  (is_as_tkeep),             // O  4
                                                  .is_as_tlast  (is_as_tlast),             // O  
                                                  .is_as_tid    (is_as_tid),               // O  2
                                                  .is_as_tvalid (is_as_tvalid),            // O  
                                                  .is_as_tuser  (is_as_tuser),             // O  2
                                                  .is_as_tready (is_as_tready),            // O  
                                                  .axi_awvalid  (axi_awvalid_s_awvalid),   // I  
                                                  .axi_awaddr   (axi_awaddr_s_awaddr),     // I  15
                                                  .axi_wvalid   (axi_wvalid_s_wvalid),     // I  
                                                  .axi_wdata    (axi_wdata_s_wdata),       // I  32
                                                  .axi_wstrb    (axi_wstrb_s_wstrb),       // I  4
                                                  .axi_arvalid  (axi_arvalid_s_arvalid),   // I  
                                                  .axi_araddr   (axi_araddr_s_araddr),     // I  15
                                                  .axi_rready   (axi_rready_s_rready),     // I  
                                                  .cc_is_enable (cc_is_enable),            // I  
                                                  .as_is_tdata  (as_is_tdata),             // I  32

                           .as_is_tupsb  (as_is_tupsb),     // I  5

                                                  .as_is_tstrb  (as_is_tstrb),             // I  4
                                                  .as_is_tkeep  (as_is_tkeep),             // I  4
                                                  .as_is_tlast  (as_is_tlast),             // I  
                                                  .as_is_tid    (as_is_tid),               // I  2
                                                  .as_is_tvalid (as_is_tvalid),            // I  
                                                  .as_is_tuser  (as_is_tuser),             // I  2
                                                  .as_is_tready (as_is_tready),            // I  
                                                  .ioclk        (ioclk),                   // I  
                                                  .serial_rxd   (serial_rxd),              // I  12
                                                  .serial_rclk  (serial_rclk),             // I  
                                                  .serial_txd   (serial_txd),              // O  12
                                                  .serial_tclk  (serial_tclk),             // O  
                                                  .axi_clk      (axi_clk),                 // I  
                                                  .axi_reset_n  (axi_reset_n),             // I  
                                                  .axis_clk     (axis_clk),                // I  
                                                  .axis_rst_n   (axis_rst_n)               // I  
                                                 );


// This code snippet was auto generated by xls2vlog.py from source file: /home/josh/Downloads/Interface-Definition.xlsx
// User: josh
// Date: Sep-22-23



LOGIC_ANLZ #(.pADDR_WIDTH( pADDR_WIDTH ),
             .pDATA_WIDTH( 32 )) U_LOGIC_ANLZ0 (
                                                .axi_awready  (axi_awready_axi_awready0),// O  
                                                .axi_wready   (axi_wready_axi_wready0),  // O  
                                                .axi_arready  (axi_arready_axi_arready0),// O  
                                                .axi_rdata    (axi_rdata_axi_rdata0),    // O  32
                                                .axi_rvalid   (axi_rvalid_axi_rvalid0),  // O  
                                                .m_tdata      (m_tdata_la_as_tdata),     // O  32
                                                .m_tstrb      (m_tstrb_la_as_tstrb),     // O  4
                                                .m_tkeep      (m_tkeep_la_as_tkeep),     // O  4
                                                .m_tlast      (m_tlast_la_as_tlast),     // O  
                                                .m_tvalid     (m_tvalid_la_as_tvalid),   // O  
                                                .m_tuser      (m_tuser_la_as_tuser),     // O  2
                                                .la_hpri_req  (la_hpri_req),             // O  
                                                .axi_awvalid  (axi_awvalid_s_awvalid),   // I  
                                                .axi_awaddr   (axi_awaddr_s_awaddr),     // I  15
                                                .axi_wvalid   (axi_wvalid_s_wvalid),     // I  
                                                .axi_wdata    (axi_wdata_s_wdata),       // I  32
                                                .axi_wstrb    (axi_wstrb_s_wstrb),       // I  4
                                                .axi_arvalid  (axi_arvalid_s_arvalid),   // I  
                                                .axi_araddr   (axi_araddr_s_araddr),     // I  15
                                                .axi_rready   (axi_rready_s_rready),     // I  
                                                .cc_la_enable (cc_la_enable),            // I  
                                                .m_tready     (as_la_tready_m_tready),   // I  
                                                .up_la_data   (up_la_data),              // I  24
                                                .user_clock2  (user_clock2),             // I  
                                                .axi_clk      (axi_clk),                 // I  
                                                .axi_reset_n  (axi_reset_n),             // I  
                                                .axis_clk     (axis_clk),                // I  
                                                .uck2_rst_n   (uck2_rst_n),              // I  
                                                .axis_rst_n   (axis_rst_n)               // I  
                                               );


// This code snippet was auto generated by xls2vlog.py from source file: /home/josh/Downloads/Interface-Definition.xlsx
// User: josh
// Date: Sep-22-23



USER_SUBSYS #(  .pUSER_PROJECT_SIDEBAND_WIDTH( pUSER_PROJECT_SIDEBAND_WIDTH ),
        .pADDR_WIDTH( pADDR_WIDTH ),
        .pDATA_WIDTH( 32 )) U_USER_SUBSYS0 (
                                                  .axi_awready  (axi_awready_axi_awready2),// O  
                                                  .axi_wready   (axi_wready_axi_wready2),  // O  
                                                  .axi_arready  (axi_arready_axi_arready2),// O  
                                                  .axi_rdata    (axi_rdata_axi_rdata2),    // O  32
                                                  .axi_rvalid   (axi_rvalid_axi_rvalid2),  // O  
                                                  .m_tdata      (m_tdata_up_as_tdata),     // O  32

                            .m_tupsb    (m_tupsb_up_as_tupsb),     // O  5

                                                  .m_tstrb      (m_tstrb_up_as_tstrb),     // O  4
                                                  .m_tkeep      (m_tkeep_up_as_tkeep),     // O  4
                                                  .m_tlast      (m_tlast_up_as_tlast),     // O  
                                                  .m_tvalid     (m_tvalid_up_as_tvalid),   // O  
                                                  .m_tuser      (m_tuser_up_as_tuser),     // O  2
                                                  .s_tready     (s_tready_up_as_tready),   // O  
                                                  .high_pri_irq (high_pri_irq_up_hpri_req),// O  
                                                  .up_la_data   (up_la_data),              // O  24
                                                  .axi_awvalid  (axi_awvalid_s_awvalid),   // I  
                                                  .axi_awaddr   (axi_awaddr_s_awaddr),     // I  15
                                                  .axi_wvalid   (axi_wvalid_s_wvalid),     // I  
                                                  .axi_wdata    (axi_wdata_s_wdata),       // I  32
                                                  .axi_wstrb    (axi_wstrb_s_wstrb),       // I  4
                                                  .axi_arvalid  (axi_arvalid_s_arvalid),   // I  
                                                  .axi_araddr   (axi_araddr_s_araddr),     // I  15
                                                  .axi_rready   (axi_rready_s_rready),     // I  
                                                  .cc_up_enable (cc_up_enable),            // I  
                                                  .user_prj_sel (user_prj_sel),            // I  5
                                                  .s_tdata      (as_up_tdata_s_tdata),     // I  32

                            .s_tupsb   (as_up_tupsb_s_tupsb),     // I  5

                                                  .s_tstrb      (as_up_tstrb_s_tstrb),     // I  4
                                                  .s_tkeep      (as_up_tkeep_s_tkeep),     // I  4
                                                  .s_tlast      (as_up_tlast_s_tlast),     // I  
                                                  .s_tvalid     (as_up_tvalid_s_tvalid),   // I  
                                                  .s_tuser      (as_up_tuser_s_tuser),     // I  2
                                                  .m_tready     (as_up_tready_m_tready),   // I  
                                                  .low__pri_irq (low__pri_irq),            // O  
                                                  .user_clock2  (user_clock2),             // I  
                                                  .axi_clk      (axi_clk),                 // I  
                                                  .axi_reset_n  (axi_reset_n),             // I  
                                                  .axis_clk     (axis_clk),                // I  
                                                  .uck2_rst_n   (uck2_rst_n),              // I  
                                                  .axis_rst_n   (axis_rst_n)               // I  
                                                 );


// This code snippet was auto generated by xls2vlog.py from source file: /home/josh/Downloads/Interface-Definition.xlsx
// User: josh
// Date: Sep-22-23



FSIC_CLKRST  U_FSIC_CLKRST0 (
                             .ioclk        (ioclk),                   // O  
                             .user_prj_sel (user_prj_sel),            // I  5
                             .mb_irq       (mb_irq),                  // I  
                             .low__pri_irq (low__pri_irq),            // I  
                             .high_pri_irq (high_pri_irq_up_hpri_req),// I  
                             .io_clk       (io_clk),                  // I  
                             .wb_rst       (wb_rst),                  // I  
                             .wb_clk       (wb_clk),                  // I  
                             .user_irq     (user_irq),                // O  3
                             .user_clock2  (user_clock2),             // I  
                             .axi_clk      (axi_clk),                 // O  
                             .axi_reset_n  (axi_reset_n),             // O  
                             .axis_clk     (axis_clk),                // O  
                             .uck2_rst_n   (uck2_rst_n),              // O  
                             .axis_rst_n   (axis_rst_n)               // O  
                            );


// This code snippet was auto generated by xls2vlog.py from source file: /home/josh/Downloads/Interface-Definition.xlsx
// User: josh
// Date: Sep-22-23


MPRJ_IO #(
      .pUSER_PROJECT_SIDEBAND_WIDTH( pUSER_PROJECT_SIDEBAND_WIDTH ),
      .pSERIALIO_WIDTH ( pSERIALIO_WIDTH ),
      .pADDR_WIDTH( pADDR_WIDTH ),
      .pDATA_WIDTH( 32 )) U_MPRJ_IO0 (
                                          .serial_rxd   (serial_rxd),              // O  12
                                          .serial_rclk  (serial_rclk),             // O  
                                          .io_clk       (io_clk),                  // O  
                                          .user_prj_sel (user_prj_sel),            // I  5
                                          .serial_txd   (serial_txd),              // I  12
                                          .serial_tclk  (serial_tclk),             // I  
                                          .io_in        (io_in),                   // I  38
                                          .vccd         (vccd),                    // I  
                                          .vssd         (vssd),                    // I  
                                          .io_out       (io_out),                  // O  38
                                          .io_oeb       (io_oeb),                  // O  38
                                          .user_clock2  (user_clock2),             // I  
                                          .axi_clk      (axi_clk),                 // I  
                                          .axi_reset_n  (axi_reset_n),             // I  
                                          .axis_clk     (axis_clk),                // I  
                                          .uck2_rst_n   (uck2_rst_n),              // I  
                                          .axis_rst_n   (axis_rst_n)               // I  
                                         );




endmodule // FSIC
// This code snippet was auto generated by xls2vlog.py from source file: /home/patrick/Downloads/Interface-Definition.xlsx
// User: patrick
// Date: Jun-06-23


module FSIC_CLKRST (
  input  wire  [4: 0] user_prj_sel,
  input  wire         mb_irq,
  input  wire         wb_rst,
  input  wire         wb_clk,
  output wire  [2: 0] user_irq,

  input  wire         low__pri_irq,
  input  wire         high_pri_irq,

  input  wire         user_clock2,
  output wire         uck2_rst_n,

  output  wire         axi_clk,
  output wire         axi_reset_n,

  output  wire         axis_clk,
  output wire         axis_rst_n,

  input  wire         io_clk,
  output wire         ioclk
);


  assign axi_clk = wb_clk;
  assign axis_clk = wb_clk;  

// ----------------------------------------------------------
// AXI-Lite
reg [2:0] axi_reset_nr; 
always @(posedge axi_clk or posedge wb_rst)
  if( wb_rst )
    axi_reset_nr <= 3'b000;
  else
    axi_reset_nr <= {axi_reset_nr[1:0], 1'b1};

assign axi_reset_n = axi_reset_nr[2];


// ----------------------------------------------------------
// AXIS
reg [2:0] axis_rst_nr; 
always @(posedge axis_clk or posedge wb_rst)
  if( wb_rst )
    axis_rst_nr <= 3'b000;
  else
    axis_rst_nr <= {axis_rst_nr[1:0], 1'b1};

assign axis_rst_n = axis_rst_nr[2];


// ----------------------------------------------------------
// user_clock2
reg [2:0] uck2_rst_nr; 
always @(posedge user_clock2 or posedge wb_rst)
  if( wb_rst )
    uck2_rst_nr <= 3'b000;
  else
    uck2_rst_nr <= {uck2_rst_nr[1:0], 1'b1};

assign uck2_rst_n = uck2_rst_nr[2];


// ----------------------------------------------------------
// IRQ
assign user_irq[2] = high_pri_irq;
assign user_irq[1] = low__pri_irq;
assign user_irq[0] = mb_irq;


// ----------------------------------------------------------
// IOCLK for IO_SERDES

/*
// TBD
reg div2_clk;
always @(posedge user_clock2 or negedge uck2_rst_n)
  if( ~uck2_rst_n )
    div2_clk <= 1'b0;
  else
    div2_clk <= ~div2_clk; 
*/

// TBD
assign ioclk = io_clk;

endmodule // FSIC_CLKRST

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Author : Tony Ho
//
//
// Create Date: 07/10/2023 11:39:49 AM
// Design Name:
// Module Name: fsic_coreclk_phase_cnt
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module fsic_coreclk_phase_cnt#(
		parameter pCLK_RATIO =4
	) (
		input wire 	axis_rst_n,
		input wire 	ioclk,
		input wire 	coreclk,
		output wire	[$clog2(pCLK_RATIO)-1:0] phase_cnt_out
	);

    reg [pCLK_RATIO-1:0] clk_seq;
    reg [$clog2(pCLK_RATIO)-1:0] phase_cnt;
    assign phase_cnt_out = phase_cnt;

	reg core_clk_toggle;
    always @(posedge coreclk or negedge axis_rst_n) begin
        if ( !axis_rst_n ) begin
            core_clk_toggle <= 0;
        end
        else begin
            core_clk_toggle <= ~core_clk_toggle;
        end
    end

	reg pre_core_clk_toggle;
	reg sync_core_clk_toggle;
	
    always @(posedge ioclk or negedge axis_rst_n) begin
        if ( !axis_rst_n ) begin
            pre_core_clk_toggle <= 0;
            sync_core_clk_toggle <= 0;
        end
        else begin
			pre_core_clk_toggle <= core_clk_toggle;
			sync_core_clk_toggle <= pre_core_clk_toggle;		//avoid metastable issue.
        end
    end


    always @(posedge ioclk or negedge axis_rst_n) begin
        if ( !axis_rst_n ) begin
            clk_seq <= 0;
        end
        else begin
            clk_seq[pCLK_RATIO-1:1] <=  clk_seq[pCLK_RATIO-2:0];
            clk_seq[0] <=  sync_core_clk_toggle;
        end
    end


    always @(posedge ioclk or negedge axis_rst_n) begin
        if ( !axis_rst_n) begin
            phase_cnt <= 0;
        end
        else begin
            if ( (clk_seq == 4'h3) || (clk_seq == 4'hc) )
                phase_cnt <= 0;
            else
                phase_cnt <= phase_cnt + 1;
        end
    end

endmodule
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Author : Tony Ho
//
//
// Create Date: 07/10/2023 11:45:06 AM
// Design Name:
// Module Name: fsic_io_serdes_rx
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
//20230724
//1. rx_sync_fifo output to rxdata_out for reduce 1T.

module fsic_io_serdes_rx#(
		parameter pRxFIFO_DEPTH = 5,
		parameter pCLK_RATIO =4
	) (
		input wire 	axis_rst_n,
		input wire 	rxclk,
		input wire   rxen,
		input wire 	ioclk,
		input wire 	coreclk,
		input wire 	Serial_Data_in,
		output wire 	[pCLK_RATIO-1:0] rxdata_out,
		output wire 	rxdata_out_valid
	);


	reg [$clog2(pRxFIFO_DEPTH)-1:0] w_ptr;
	reg w_ptr_pre;
	reg w_ptr_sync;
	wire rx_shift_reg_valid;

	wire w_ptr_graycode_bit0;

	assign w_ptr_graycode_bit0 = w_ptr[1] ^  w_ptr[0];

	wire rxen_rst_n = axis_rst_n & rxen;

	always @(negedge rxclk or negedge rxen_rst_n)  begin
		if ( !rxen_rst_n ) begin
			w_ptr <= 0;
		end
		else begin
			if (w_ptr == 4)
				w_ptr <= 0;
			else
				w_ptr <= w_ptr+1;
		end
	end


	reg [pRxFIFO_DEPTH-1:0] RxFifo;


	always @(negedge rxclk or negedge rxen_rst_n) begin
		if ( !rxen_rst_n ) begin
			RxFifo <= 0;
		end
		else begin
			RxFifo[w_ptr] <= Serial_Data_in;
		end
	end



	always @(posedge ioclk or negedge axis_rst_n)  begin
		if ( !axis_rst_n ) begin
			w_ptr_pre <= 0;
			w_ptr_sync <= 0;
		end
		else begin
			w_ptr_pre <= w_ptr_graycode_bit0;		//use gray code
			w_ptr_sync <= w_ptr_pre;				//avoid metastable issue
		end
	end

	reg rx_start;
	always @(posedge ioclk or negedge axis_rst_n)  begin
		if ( !axis_rst_n ) begin
			rx_start <= 0;
		end
		else begin
			if (w_ptr_sync != 0 )
				rx_start <= 1;
			else
				rx_start <= rx_start;
		end
	end


	reg [$clog2(pRxFIFO_DEPTH)-1:0] r_ptr;

	always @(posedge ioclk or negedge axis_rst_n)  begin
		if ( !axis_rst_n ) begin
			r_ptr <= 0;
		end
		else begin
			if (rx_start) begin
				if ( r_ptr == 4 )
					r_ptr <= 0;
				else
					r_ptr <= r_ptr + 1;
			end
			else
				r_ptr <= r_ptr;
		end
	end

	reg [pCLK_RATIO-1:0] rx_shift_reg;

	always @(posedge ioclk or negedge axis_rst_n)  begin
		if ( !axis_rst_n ) begin
			rx_shift_reg <= 0;
		end
		else begin
			if (rx_start) begin
				rx_shift_reg[3] <= RxFifo[r_ptr];		//r_ptr get from LSB to MSB
				rx_shift_reg[2:0] <= rx_shift_reg[3:1];
			end
		end
	end

	reg [$clog2(pCLK_RATIO)-1:0] rx_shift_phase_cnt;

	always @(posedge ioclk or negedge axis_rst_n)  begin
		if ( !axis_rst_n ) begin
			rx_shift_phase_cnt <= pCLK_RATIO-1;
		end
		else begin
			if (rx_start)
				rx_shift_phase_cnt <= rx_shift_phase_cnt+1;
			else
				rx_shift_phase_cnt <= rx_shift_phase_cnt;
		end
	end

	reg [2:0] rx_start_delay;

	always @(posedge ioclk or negedge axis_rst_n)  begin
		if ( !axis_rst_n ) begin
			rx_start_delay <= 0;
		end
		else begin
			rx_start_delay[0] <= rx_start;
			rx_start_delay[2:1] <= rx_start_delay[1:0];
		end
	end

	assign rx_shift_reg_valid = (rx_shift_phase_cnt == pCLK_RATIO-1) && rx_start_delay[2] ; //rx_shift_reg is ready to move.

	//write by ioclk in negedge and read by coreclk in posedge then simulation result is ok.

	reg [pCLK_RATIO-1:0] rx_sync_fifo;
	reg rx_sync_fifo_valid;

	always @(negedge ioclk or negedge axis_rst_n)  begin		// Note : the FPGA provide both coreclk and ioclk to FSIC_SOC, the skew of coreclk and ioclk maybe impact by FPGA output timining -> PCB -> FSIC_SOC input timing.
																// when ioclok early then coreclk in fsic_io_serdes_rx, it may cause hold time issue in rx_shift_reg to rx_sync_fifo.
																// use negdege ioclk to improve the hold time, but it sacrifice the setup time. 
		if ( !axis_rst_n ) begin
			rx_sync_fifo <= 0;
			rx_sync_fifo_valid <= 0;
		end
		else begin
			if (rx_start && rx_shift_reg_valid)  begin
				rx_sync_fifo <= rx_shift_reg;
				rx_sync_fifo_valid <= 1;
			end
			else begin
				rx_sync_fifo <= rx_sync_fifo;
				rx_sync_fifo_valid <= rx_sync_fifo_valid;
			end
		end
	end

	assign rxdata_out = rx_sync_fifo;
	assign rxdata_out_valid = rx_sync_fifo_valid;

/*
	reg [pCLK_RATIO-1:0] rxdata;
	reg rxdata_valid;

	assign rxdata_out = rxdata;
	assign rxdata_out_valid = rxdata_valid;

	always @(posedge coreclk or negedge axis_rst_n)  begin
		if ( !axis_rst_n ) begin
			rxdata <= 0;
			rxdata_valid <= 0;
		end
		else begin
				rxdata <= rx_sync_fifo;
				rxdata_valid <= rx_sync_fifo_valid;
		end
	end
*/


endmodule

// This code snippet was auto generated by xls2vlog.py from source file: /home/patrick/Downloads/Interface-Definition.xlsx
// User: patrick
// Date: Jul-19-23



module MPRJ_IO #(   parameter pUSER_PROJECT_SIDEBAND_WIDTH   = 5,
          parameter pSERIALIO_WIDTH   = 13,
          parameter pADDR_WIDTH   = 12,
          parameter pDATA_WIDTH   = 32
                )
(
  input  wire          vccd,
  input  wire          vssd,
  output wire  [pSERIALIO_WIDTH-1: 0] serial_rxd,
  output wire          serial_rclk,
  input  wire   [4: 0] user_prj_sel,
  input  wire  [pSERIALIO_WIDTH-1: 0] serial_txd,
  input  wire          serial_tclk,
  input  wire  [37: 0] io_in,
  output wire  [37: 0] io_out,
  output wire  [37: 0] io_oeb,
  output wire          io_clk,
  input  wire          user_clock2,
  input  wire          axi_clk,
  input  wire          axi_reset_n,
  input  wire          axis_clk,
  input  wire          uck2_rst_n,
  input  wire          axis_rst_n
);

  localparam BASE_OFFSET = 8;
  localparam RXD_OFFSET = BASE_OFFSET;
  localparam RXCLK_OFFSET = RXD_OFFSET + pSERIALIO_WIDTH;
  localparam TXD_OFFSET = RXCLK_OFFSET + 1;
  localparam TXCLK_OFFSET = TXD_OFFSET + pSERIALIO_WIDTH;
  localparam IOCLK_OFFSET = TXCLK_OFFSET + 1;
  localparam TXRX_WIDTH = IOCLK_OFFSET - BASE_OFFSET + 1;

// MPRJ_IO PIN PLANNING when pSERIALIO_WIDTH=13
// --------------------------------
// [20: 8]  I   RXD
// [   21]  I   RXCLK

// --------------------------------
// [34:22]  O   TXD
// [   35]  O   TXCLK

// --------------------------------
// [   36]  I   IO_CLK

// MPRJ_IO PIN PLANNING when pSERIALIO_WIDTH=12
// --------------------------------
// [19: 8]  I   RXD
// [   20]  I   RXCLK

// --------------------------------
// [32:21]  O   TXD
// [   33]  O   TXCLK

// --------------------------------
// [   34]  I   IO_CLK

/*
assign serial_rxd    = 12'b0;
assign serial_rclk   = 1'b0;
assign io_out        = 38'b0;
assign io_oeb        = 38'b0;
*/

assign io_clk = io_in[IOCLK_OFFSET];

assign io_oeb[ 7: 0]   =  8'h00;

assign io_oeb[RXD_OFFSET +: pSERIALIO_WIDTH]   = ~32'b0;  // RXD
assign io_oeb[RXCLK_OFFSET]   =  1'b1;    // RX_CLK

assign io_oeb[TXD_OFFSET +: pSERIALIO_WIDTH]   = 32'b0;  // TXD
assign io_oeb[TXCLK_OFFSET]   =  1'b0;    // TX_CLK

assign io_oeb[IOCLK_OFFSET]   =  1'b1;    // IO_CLK (from FPGA)

//assign value to avoid dc_shell report warning
//below setting only for pSERIALIO_WIDTH=13, for pSERIALIO_WIDTH=12 need change the hard code setting.
assign io_oeb[ 37]   =  1'b0; 		//for pSERIALIO_WIDTH=13
//assign io_oeb[ 37:35]   =  3'b0; 		//for pSERIALIO_WIDTH=12

assign serial_rxd  = io_in[RXD_OFFSET +: pSERIALIO_WIDTH];
assign serial_rclk = io_in[RXCLK_OFFSET];

assign io_out[TXD_OFFSET +: pSERIALIO_WIDTH] = serial_txd;
assign io_out[TXCLK_OFFSET] = serial_tclk;

//assign value to avoid dc_shell report warning
assign io_out[21:0] = 32'b0; 			//for pSERIALIO_WIDTH=13
assign io_out[37:36] = 2'b0; 			//for pSERIALIO_WIDTH=13
//assign io_out[20:0] = 32'b0; 		//for pSERIALIO_WIDTH=12
//assign io_out[37:34] = 4'b0; 		//for pSERIALIO_WIDTH=12

endmodule // MPRJ_IO


`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Author : Tony Ho
//
// Create Date: 06/18/2023 10:44:18 PM
// Design Name:
// Module Name: IO_SERDES
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
// 20230720
// 1. change pADDR_WIDTH=15 and use [pADDR_WIDTH-1:0] for *_axi_awaddr and *_axi_araddr
// 20230714
// 1. change [pADDR_WIDTH-1:0] axi_awaddr to [pADDR_WIDTH+1:2] axi_awaddr for DW base address
// 2. add pSERIALIO_WIDTH and pSERIALIO_TDATA_WIDTH
// 3. add is_as_dummy for remove WARNING message
// 4. update typo in pSERIALIO_TDATA_WIDTH
// 5. update tpyo, change cc_ls_enable to cc_is_enable
// 20230712
// 1. axi_awaddr is DW address, pADDR_WIDTH change from 12 to 10
// 2. define USE_FOR_LOOP_Serial_Data_Out_tdata and update coding error in for loop

`define USE_FOR_LOOP_Serial_Data_Out_tdata 1

module IO_SERDES #(
    parameter pUSER_PROJECT_SIDEBAND_WIDTH   = 5,
    parameter pSERIALIO_WIDTH   = 13,
    parameter pADDR_WIDTH   = 15,
    parameter pDATA_WIDTH   = 32,
    parameter pRxFIFO_DEPTH = 5,
    parameter pCLK_RATIO =4      //[TODO]: use pCLK_RATIO for register define
  ) (


    input wire   ioclk,

    input wire   axi_reset_n,
    input wire   axi_clk,

    input wire   axis_rst_n,
    input wire   axis_clk,

    //write addr channel
    input wire   axi_awvalid,
    input wire   [pADDR_WIDTH-1:0] axi_awaddr,    //axi_awaddr is DW address
    output wire  axi_awready,

    //write data channel
    input wire   axi_wvalid,
    input wire   [pDATA_WIDTH-1:0] axi_wdata,
    input wire   [(pDATA_WIDTH/8)-1:0] axi_wstrb,
    output wire  axi_wready,

    //read addr channel
    input wire   axi_arvalid,
    input wire   [pADDR_WIDTH-1:0] axi_araddr,
    output wire   axi_arready,

    //read data channel
    output wire   axi_rvalid,
    output wire   [pDATA_WIDTH-1:0] axi_rdata,
    input wire   axi_rready,

    input wire   cc_is_enable,    //axi_lite enable



    //TX path
    input wire   [pDATA_WIDTH-1:0] as_is_tdata,
    input wire   [pUSER_PROJECT_SIDEBAND_WIDTH-1:0] as_is_tupsb,
    input wire   [(pDATA_WIDTH/8)-1:0] as_is_tstrb,
    input wire   [(pDATA_WIDTH/8)-1:0] as_is_tkeep,
    input wire   as_is_tlast,
    input wire   [1:0] as_is_tid,
    input wire   as_is_tvalid,
    input wire   [1:0] as_is_tuser,
    input wire   as_is_tready,    //when local side axis switch Rxfifo size <= threshold then as_is_tready=0, this flow control mechanism is for notify remote side do not provide data with is_as_tvalid=1
    output wire rxen_out,   //output rxen for post synthsis simultation

    output wire      serial_tclk,
    output wire  [pSERIALIO_WIDTH-1: 0] serial_txd,

    //Rx path
    input  wire      serial_rclk,
    input  wire  [pSERIALIO_WIDTH-1: 0] serial_rxd,

    output wire   [pDATA_WIDTH-1:0] is_as_tdata,
    output wire   [pUSER_PROJECT_SIDEBAND_WIDTH-1:0] is_as_tupsb,
    output wire   [(pDATA_WIDTH/8)-1:0] is_as_tstrb,
    output wire   [(pDATA_WIDTH/8)-1:0] is_as_tkeep,
    output wire   is_as_tlast,
    output wire   [1:0] is_as_tid,
    output wire   is_as_tvalid,
    output wire   [1:0] is_as_tuser,
    output wire   is_as_tready    //when remote side axis switch Rxfifo size <= threshold then is_as_tready=0, this flow control mechanism is for notify local side do not provide data with as_is_tvalid=1

  );

  localparam pSERIALIO_TDATA_WIDTH  = pDATA_WIDTH/pCLK_RATIO;
  
  wire coreclk;
  wire txclk;
  wire rxclk;
  wire axi_awvalid_in;
  wire axi_wvalid_in;
  wire txen_out;
  wire is_as_tready_remote;
  
  assign coreclk = axis_clk;
  assign serial_tclk = txclk;
  assign rxclk = serial_rclk;


  wire Serial_Data_Out_tupsb_4_1;
  wire Serial_Data_Out_tupsb_tlast_tvalid_tready;
  wire Serial_Data_Out_tid_tuser;
  wire Serial_Data_Out_tkeep;
  wire Serial_Data_Out_tstrb;
  wire [pSERIALIO_TDATA_WIDTH-1:0] Serial_Data_Out_tdata;

    assign   serial_txd[pSERIALIO_WIDTH-1:0] = {Serial_Data_Out_tupsb_4_1, Serial_Data_Out_tupsb_tlast_tvalid_tready, Serial_Data_Out_tid_tuser, Serial_Data_Out_tkeep, Serial_Data_Out_tstrb, Serial_Data_Out_tdata[pSERIALIO_TDATA_WIDTH-1:0]};



    wire Serial_Data_In_tupsb_4_1;
    wire Serial_Data_In_tupsb_tlast_tvalid_tready;

  wire Serial_Data_In_tid_tuser;
  wire Serial_Data_In_tkeep;
  wire Serial_Data_In_tstrb;
  wire [pSERIALIO_TDATA_WIDTH-1:0] Serial_Data_In_tdata;

    assign {Serial_Data_In_tupsb_4_1, Serial_Data_In_tupsb_tlast_tvalid_tready, Serial_Data_In_tid_tuser, Serial_Data_In_tkeep, Serial_Data_In_tstrb, Serial_Data_In_tdata[pSERIALIO_TDATA_WIDTH-1:0] } = serial_rxd[pSERIALIO_WIDTH-1:0];



  reg  txen;

  //register offset 0
  reg rxen_ctl;  //bit 0
  reg txen_ctl;  //bit 1

  //write addr channel
  assign   axi_awvalid_in  = axi_awvalid && cc_is_enable;
  wire axi_awready_out;
  assign axi_awready = axi_awready_out;

  //write data channel
  assign   axi_wvalid_in  = axi_wvalid && cc_is_enable;
  wire axi_wready_out;
  assign axi_wready = axi_wready_out;

  // if both axi_awvalid_in=1 and axi_wvalid_in=1 then output axi_awready_out = 1 and axi_wready_out = 1
  assign axi_awready_out = (axi_awvalid_in && axi_wvalid_in) ? 1'b1 : 1'b0;
  assign axi_wready_out = (axi_awvalid_in && axi_wvalid_in) ? 1'b1 : 1'b0;


  //write register
  always @(posedge axi_clk or negedge axi_reset_n)  begin
    if ( !axi_reset_n ) begin
      rxen_ctl <= 0;
      txen_ctl <= 0;
    end
    else begin
      if ( axi_awvalid_in && axi_wvalid_in ) begin    //when axi_awvalid_in=1 and axi_wvalid_in=1 means axi_awready_out=1 and axi_wready_out=1
        if (axi_awaddr[11:2] == 10'h000 && (axi_wstrb[0] == 1) ) begin //offset 0
          rxen_ctl <= axi_wdata[0];
          txen_ctl <= axi_wdata[1];
        end
        else begin
          rxen_ctl <= rxen_ctl;
          txen_ctl <= txen_ctl;
        end
      end
    end
  end


  // io serdes always output axi_arready = 1 and don't care the axi_arvalid & axi_araddr
  // io serdes only support 2 register bits in offset 0. config read other address offset is reserved.
  assign axi_arready = 1;
  // io serdes always output axi_rvalid = 1 and axi_rdata =  { 30'b0, txen_ctl, rxen_ctl }
  assign axi_rvalid = 1;
  assign axi_rdata =  { 30'b0, txen_ctl, rxen_ctl };



  assign txen_out = txen;

  wire [$clog2(pCLK_RATIO)-1:0] phase_cnt;

  fsic_coreclk_phase_cnt  #(
    .pCLK_RATIO(pCLK_RATIO)
  )
  fsic_coreclk_phase_cnt_0(
    .axis_rst_n(axis_rst_n),
    .ioclk(ioclk),
    .coreclk(coreclk),
    .phase_cnt_out(phase_cnt)
  );


// For Tx Path

  wire  rx_received_data;


  always @(negedge ioclk or negedge axis_rst_n)  begin
    if ( !axis_rst_n ) begin
      txen <= 0;
    end
    else begin
      if ( (txen_ctl || rx_received_data) && phase_cnt == 3   )  // set txen=1 when timeout or rx_received_data==1
                                      // if rx_received_data==1 before timeout, it means remote side txen is ealry then local side.
                                      // then we should set local site txen=1 to allow local site provide ready signal to remote side in tx path.
                                      // It is to avoid local site rx fifo full in axis switch.
        txen <= 1;
      else
        txen <= txen;
    end
  end

  reg [$clog2(pCLK_RATIO)-1:0] tx_shift_phase_cnt;


  always @(posedge ioclk or negedge axis_rst_n)  begin
    if ( !axis_rst_n ) begin
      tx_shift_phase_cnt <= 3;
    end
    else begin
      if (txen)
        tx_shift_phase_cnt <= tx_shift_phase_cnt + 1;
      else
        tx_shift_phase_cnt <= tx_shift_phase_cnt;
    end
  end

  reg [pDATA_WIDTH-1:0] pre_as_is_tdata_buf;
  reg [(pDATA_WIDTH/8)-1:0] pre_as_is_tstrb_buf;
  reg [(pDATA_WIDTH/8)-1:0] pre_as_is_tkeep_buf;
  reg [(pDATA_WIDTH/8)-1:0] pre_as_is_tid_tuser_buf;


    reg [3:0] pre_as_is_tupsb_4_1_buf;
    reg [(pDATA_WIDTH/8)-1:0] pre_as_is_tupsb_tlast_tvalid_tready_buf;


  wire txen_rst_n = axis_rst_n & txen;

  always @(negedge coreclk or negedge txen_rst_n)  begin

    if ( !txen_rst_n ) begin
      pre_as_is_tdata_buf <= 0;
      pre_as_is_tstrb_buf <= 0;
      pre_as_is_tkeep_buf <= 0;
      pre_as_is_tid_tuser_buf <= 0;

        pre_as_is_tupsb_4_1_buf <= 0;
        pre_as_is_tupsb_tlast_tvalid_tready_buf <= 0;

    end 
    else begin
      pre_as_is_tdata_buf <= as_is_tdata;
      pre_as_is_tstrb_buf <= as_is_tstrb;
      pre_as_is_tkeep_buf <= as_is_tkeep;
      pre_as_is_tid_tuser_buf[3:2] <= as_is_tid;
      pre_as_is_tid_tuser_buf[1:0] <= as_is_tuser;

        pre_as_is_tupsb_4_1_buf <= as_is_tupsb[pUSER_PROJECT_SIDEBAND_WIDTH-1:1];
        pre_as_is_tupsb_tlast_tvalid_tready_buf[3] <= as_is_tupsb[0];
        pre_as_is_tupsb_tlast_tvalid_tready_buf[2] <= as_is_tlast;
        pre_as_is_tupsb_tlast_tvalid_tready_buf[1] <= as_is_tvalid;
        pre_as_is_tupsb_tlast_tvalid_tready_buf[0] <= as_is_tready;

      
      if (is_as_tready && as_is_tvalid) begin      //data transfer from Axis siwtch to io serdes when is_as_tready=1 and as_is_tvalid=1
        

          pre_as_is_tupsb_tlast_tvalid_tready_buf[1] <= as_is_tvalid;

      end
      else begin

          pre_as_is_tupsb_tlast_tvalid_tready_buf[1] <= 0;      // set as_is_tvalid =0 to remote side

      end
    end
  end

  reg [pDATA_WIDTH-1:0] as_is_tdata_buf;
  reg [(pDATA_WIDTH/8)-1:0] as_is_tstrb_buf;
  reg [(pDATA_WIDTH/8)-1:0] as_is_tkeep_buf;
  reg [(pDATA_WIDTH/8)-1:0] as_is_tid_tuser_buf;

    reg [pCLK_RATIO-1:0] as_is_tupsb_4_1_buf;
    reg [pCLK_RATIO-1:0] as_is_tupsb_tlast_tvalid_tready_buf;    


  always @(posedge ioclk or negedge axis_rst_n)  begin
    if ( !axis_rst_n ) begin
      as_is_tdata_buf <= 0;
      as_is_tstrb_buf <= 0;
      as_is_tkeep_buf <= 0;
      as_is_tid_tuser_buf <= 0;

        as_is_tupsb_4_1_buf <= 0;
        as_is_tupsb_tlast_tvalid_tready_buf <= 0;

    end
    else begin
      if (phase_cnt == 3) begin      //update as_is_*_buf when phase_cnt == 3
        as_is_tdata_buf <= pre_as_is_tdata_buf;
        as_is_tstrb_buf <= pre_as_is_tstrb_buf;
        as_is_tkeep_buf <= pre_as_is_tkeep_buf;
        as_is_tid_tuser_buf <= pre_as_is_tid_tuser_buf;
          as_is_tupsb_4_1_buf <= pre_as_is_tupsb_4_1_buf;
          as_is_tupsb_tlast_tvalid_tready_buf <= pre_as_is_tupsb_tlast_tvalid_tready_buf;

      end
    end
  end

  assign txclk = ioclk&txen;    //use negedge to avoid glitch in txclk.



  genvar j;
  generate
    for (j=0; j<pSERIALIO_TDATA_WIDTH; j=j+1 ) begin
      assign Serial_Data_Out_tdata[j] = as_is_tdata_buf[j*4+tx_shift_phase_cnt] & txen ;
    end
  endgenerate



  assign Serial_Data_Out_tstrb = as_is_tstrb_buf[tx_shift_phase_cnt] & txen ;
  assign Serial_Data_Out_tkeep = as_is_tkeep_buf[tx_shift_phase_cnt] & txen ;
  assign Serial_Data_Out_tid_tuser = as_is_tid_tuser_buf[tx_shift_phase_cnt] & txen ;

    assign Serial_Data_Out_tupsb_4_1 = as_is_tupsb_4_1_buf[tx_shift_phase_cnt] & txen ;
    assign Serial_Data_Out_tupsb_tlast_tvalid_tready = as_is_tupsb_tlast_tvalid_tready_buf[tx_shift_phase_cnt] & txen ;




// For Rx Path

    wire rxdata_out_valid[pSERIALIO_TDATA_WIDTH+3:0];    //add dummy connection to avoid WARNING message by xelab


  reg  rxen;
  assign rxen_out = rxen;

  always @(negedge ioclk or negedge axis_rst_n)  begin
    if ( !axis_rst_n ) begin
      rxen <= 0;
    end
    else begin
      if (rxen_ctl)
        rxen <= 1;
      else
        rxen <= rxen;
    end
  end


  genvar i;
  generate
    for (i=0; i<pSERIALIO_TDATA_WIDTH; i=i+1 ) begin

      fsic_io_serdes_rx  #(
        .pRxFIFO_DEPTH(pRxFIFO_DEPTH),
        .pCLK_RATIO(pCLK_RATIO)
      )
      fsic_io_serdes_rx_tdata(
        .axis_rst_n(axis_rst_n),
        .rxclk(rxclk),
        .rxen(rxen),
        .ioclk(ioclk),
        .coreclk(coreclk),
        .Serial_Data_in(Serial_Data_In_tdata[i]),
        .rxdata_out(is_as_tdata[i*4+3:i*4]),
        .rxdata_out_valid(rxdata_out_valid[i])
      );

    end
  endgenerate


  fsic_io_serdes_rx  #(
    .pRxFIFO_DEPTH(pRxFIFO_DEPTH),
    .pCLK_RATIO(pCLK_RATIO)
  )
  fsic_io_serdes_rx_tstrb(
    .axis_rst_n(axis_rst_n),
    .rxclk(rxclk),
    .rxen(rxen),
    .ioclk(ioclk),
    .coreclk(coreclk),
    .Serial_Data_in(Serial_Data_In_tstrb),
    .rxdata_out(is_as_tstrb),
    .rxdata_out_valid(rxdata_out_valid[pSERIALIO_TDATA_WIDTH])
  );


  fsic_io_serdes_rx  #(
    .pRxFIFO_DEPTH(pRxFIFO_DEPTH),
    .pCLK_RATIO(pCLK_RATIO)
  )
  fsic_io_serdes_rx_tkeep(
    .axis_rst_n(axis_rst_n),
    .rxclk(rxclk),
    .rxen(rxen),
    .ioclk(ioclk),
    .coreclk(coreclk),
    .Serial_Data_in(Serial_Data_In_tkeep),
    .rxdata_out(is_as_tkeep),
    .rxdata_out_valid(rxdata_out_valid[pSERIALIO_TDATA_WIDTH+1])
  );

  fsic_io_serdes_rx  #(
    .pRxFIFO_DEPTH(pRxFIFO_DEPTH),
    .pCLK_RATIO(pCLK_RATIO)
  )
  fsic_io_serdes_rx_tid_tuser(
    .axis_rst_n(axis_rst_n),
    .rxclk(rxclk),
    .rxen(rxen),
    .ioclk(ioclk),
    .coreclk(coreclk),
    .Serial_Data_in(Serial_Data_In_tid_tuser),
    .rxdata_out( {is_as_tid[1:0], is_as_tuser[1:0]}),
    .rxdata_out_valid(rxdata_out_valid[pSERIALIO_TDATA_WIDTH+2])
  );


    fsic_io_serdes_rx  #(
      .pRxFIFO_DEPTH(pRxFIFO_DEPTH),
      .pCLK_RATIO(pCLK_RATIO)
    )
    fsic_io_serdes_rx_upsb(
      .axis_rst_n(axis_rst_n),
      .rxclk(rxclk),
      .rxen(rxen),
      .ioclk(ioclk),
      .coreclk(coreclk),
      .Serial_Data_in(Serial_Data_In_tupsb_4_1),
      .rxdata_out( is_as_tupsb[4:1]),    
      .rxdata_out_valid(rxdata_out_valid[pSERIALIO_TDATA_WIDTH+3])
    );
  
    fsic_io_serdes_rx  #(
      .pRxFIFO_DEPTH(pRxFIFO_DEPTH),
      .pCLK_RATIO(pCLK_RATIO)
    )
    fsic_io_serdes_rx_fc(
      .axis_rst_n(axis_rst_n),
      .rxclk(rxclk),
      .rxen(rxen),
      .ioclk(ioclk),
      .coreclk(coreclk),
      .Serial_Data_in(Serial_Data_In_tupsb_tlast_tvalid_tready),
      .rxdata_out( {is_as_tupsb[0], is_as_tlast, is_as_tvalid, is_as_tready_remote}),    
      .rxdata_out_valid(rx_received_data)
    );


  reg is_as_tready_out;
  assign is_as_tready = is_as_tready_out;

  always @(posedge coreclk or negedge txen_rst_n )  begin
    if ( !txen_rst_n ) begin
      is_as_tready_out <= 0;        //set is_as_tready_out=0 when txen == 0
    end
    else begin
      if (rx_received_data == 0) is_as_tready_out <= 1;    // when txen==1 and still not recevies data from remote side then set is_as_tready_out=1 to avoid dead lock issue.
      else  is_as_tready_out <= is_as_tready_remote;        // when txen == 1 and rx_received_data==1 (received data from remote side) then is_as_tready_out come from is_as_tready_remote (remote side)
    end
  end


endmodule




//////////////////////////////////////////////////////////////////////////////////
// Author : Tony Ho
//
// Create Date: 11/20/2023
// Design Name:
// Module Name: IRQ_MUX
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module IRQ_MUX #( parameter pADDR_WIDTH=10
                )
(
  input  wire         low__pri_irq_0,
  input  wire         High_pri_req_0,
  input  wire         low__pri_irq_1,
  input  wire         High_pri_req_1,
  input  wire         low__pri_irq_2,
  input  wire         High_pri_req_2,
  input  wire         low__pri_irq_3,
  input  wire         High_pri_req_3,
  output wire         low__pri_irq,
  output wire         high_pri_irq,
  input  wire         axi_clk,
  input  wire         axi_reset_n,
  input  wire         axis_rst_n,
  input  wire  [4: 0] user_prj_sel
);


assign low__pri_irq = (user_prj_sel == 5'b00000) ? low__pri_irq_0 :
                      (user_prj_sel == 5'b00001) ? low__pri_irq_1 :
                      (user_prj_sel == 5'b00010) ? low__pri_irq_2 :
                      (user_prj_sel == 5'b00011) ? low__pri_irq_3 :
                      1'b0;
                      
assign high_pri_irq = (user_prj_sel == 5'b00000) ? High_pri_req_0 :
                      (user_prj_sel == 5'b00001) ? High_pri_req_1 :
                      (user_prj_sel == 5'b00010) ? High_pri_req_2 :
                      (user_prj_sel == 5'b00011) ? High_pri_req_3 :
                      1'b0;


endmodule // IRQ_MUX

//////////////////////////////////////////////////////////////////////////////////
// Author : Tony Ho
//
// Create Date: 11/20/2023
// Design Name:
// Module Name: LA_MUX
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module LA_MUX #( parameter pADDR_WIDTH   = 12,
                 parameter pDATA_WIDTH   = 32
               )
(
  input  wire  [23: 0] la_data_0,
  input  wire  [23: 0] la_data_1,
  input  wire  [23: 0] la_data_2,
  input  wire  [23: 0] la_data_3,
  output wire  [23: 0] up_la_data,
  input  wire          axi_clk,
  input  wire          axis_clk,
  input  wire          axi_reset_n,
  input  wire          axis_rst_n,
  input  wire   [4: 0] user_prj_sel
);


assign up_la_data = (user_prj_sel == 5'b00000) ? la_data_0 :
                    (user_prj_sel == 5'b00001) ? la_data_1 :
                    (user_prj_sel == 5'b00010) ? la_data_2 :
                    (user_prj_sel == 5'b00011) ? la_data_3 :
                    24'b0;

endmodule // LA_MUX

`timescale 1ns / 1ps
module AXIS_SW #(
				parameter pUSER_PROJECT_SIDEBAND_WIDTH   = 5,
				parameter pADDR_WIDTH   = 10,
                parameter pDATA_WIDTH   = 32
                )
(
    input  wire                             axi_reset_n,    
    input  wire                             axis_clk,
    input  wire                             axis_rst_n,
 
    //axi_lite slave interface
    //write addr channel
    input wire 	axi_awvalid,
    input wire 	[14:0] axi_awaddr,		
	output wire	axi_awready,
	//write data channel
	input wire 	axi_wvalid,
	input wire 	[pDATA_WIDTH-1:0] axi_wdata,
	input wire 	[(pDATA_WIDTH/8)-1:0] axi_wstrb,
	output wire	axi_wready,
	//read addr channel
	input wire 	axi_arvalid,
	input wire 	[14:0] axi_araddr,
	output wire axi_arready,
	//read data channel
	output wire axi_rvalid,
	output wire [pDATA_WIDTH-1:0] axi_rdata,
	input wire 	axi_rready,
	input wire 	cc_as_enable,		//axi_lite enable        
    //AXI Stream inputs for User Project grant 0
    input  wire [pDATA_WIDTH-1:0]           up_as_tdata,
		input wire 	[pUSER_PROJECT_SIDEBAND_WIDTH-1:0] up_as_tupsb,
    input  wire [pDATA_WIDTH/8-1:0]         up_as_tstrb,
    input  wire [pDATA_WIDTH/8-1:0]         up_as_tkeep,  
    input  wire                             up_as_tlast,      
    input  wire                             up_as_tvalid,
    input  wire [1:0]                       up_as_tuser, 
	input  wire                             up_hpri_req,
    output wire                             as_up_tready,
    //AXI Stream inputs for Axis Axilite grant 1
    input  wire [pDATA_WIDTH-1:0]           aa_as_tdata,
    input  wire [pDATA_WIDTH/8-1:0]         aa_as_tstrb,
    input  wire [pDATA_WIDTH/8-1:0]         aa_as_tkeep,   
    input  wire                             aa_as_tlast,       
    input  wire                             aa_as_tvalid,
    input  wire [1:0]                       aa_as_tuser,       
    output wire                             as_aa_tready,
    //AXI Stream inputs for Logic Analyzer grant 2
    input  wire [pDATA_WIDTH-1:0]           la_as_tdata,
    input  wire [pDATA_WIDTH/8-1:0]         la_as_tstrb,
    input  wire [pDATA_WIDTH/8-1:0]         la_as_tkeep, 
    input  wire                             la_as_tlast,          
    input  wire                             la_as_tvalid,
    input  wire [1:0]                       la_as_tuser,      
	input  wire                             la_hpri_req,
    output wire                             as_la_tready,
    //AXI Stream outputs for IO Serdes
    output  wire [pDATA_WIDTH-1:0]          as_is_tdata,

		output wire 	[pUSER_PROJECT_SIDEBAND_WIDTH-1:0] as_is_tupsb,
    output  wire [pDATA_WIDTH/8-1:0]        as_is_tstrb,
    output  wire [pDATA_WIDTH/8-1:0]        as_is_tkeep, 
    output  wire                            as_is_tlast,        
    output  wire [1:0]                      as_is_tid, 
    output  wire                            as_is_tvalid,
    output  wire [1:0]                      as_is_tuser,     
    input	wire                            is_as_tready,
    //Demux
    //AXI Input Stream for IO_Serdes
    input  wire [pDATA_WIDTH-1:0]           is_as_tdata,

		input wire 	[pUSER_PROJECT_SIDEBAND_WIDTH-1:0] is_as_tupsb,

    input  wire [pDATA_WIDTH/8-1:0]         is_as_tstrb,    
    input  wire [pDATA_WIDTH/8-1:0]         is_as_tkeep,
    input  wire                             is_as_tlast,
    input  wire [1:0]                       is_as_tid,
    input  wire                             is_as_tvalid,
    input  wire [1:0]                       is_as_tuser,
    output wire                             as_is_tready,
    //AXI Output Stream for User Project
    output wire [pDATA_WIDTH-1:0]           as_up_tdata,

		output wire 	[pUSER_PROJECT_SIDEBAND_WIDTH-1:0] as_up_tupsb,

    output wire [pDATA_WIDTH/8-1:0]         as_up_tstrb,    
    output wire [pDATA_WIDTH/8-1:0]         as_up_tkeep,
    output wire                             as_up_tlast,
    output wire                             as_up_tvalid,
    output wire [1:0]                       as_up_tuser,    
    input  wire                             up_as_tready,   
    //AXI Output Stream for Axis_Axilite
    output wire [pDATA_WIDTH-1:0]           as_aa_tdata,
    output wire [pDATA_WIDTH/8-1:0]         as_aa_tstrb,    
    output wire [pDATA_WIDTH/8-1:0]         as_aa_tkeep,
    output wire                             as_aa_tlast,    
    output wire                             as_aa_tvalid,
    output wire [1:0]                       as_aa_tuser, 
    input  wire                             aa_as_tready
);
localparam  USER_WIDTH = 2;
localparam  TID_WIDTH = 2;   
//for arbiter
localparam N = 3; //Upstream master Num for Input port
//source 0 support req/hi_req for user project
//source 1 support req for axilite_axis
//source 2 support req/hi_req for Logic Analyzer
localparam req_mask = 3'b111; //normal request mask for Upstream
localparam hi_req_mask = 3'b101; //high request mask for Upstream 
localparam last_support = 3'b000; //last signal support for hi request
//for Demux
// FIFO depth
localparam  FIFO_DEPTH = 16;   
//FIFO address width
localparam ADDR_WIDTH   = $clog2(FIFO_DEPTH);
//field offset for mem unit 

	localparam UPSB_OFFSET  = pDATA_WIDTH;
	localparam STRB_OFFSET  = UPSB_OFFSET + pUSER_PROJECT_SIDEBAND_WIDTH;

localparam KEEP_OFFSET  = STRB_OFFSET + pDATA_WIDTH/8;
localparam LAST_OFFSET  = KEEP_OFFSET + pDATA_WIDTH/8;
localparam TID_OFFSET   = LAST_OFFSET + 1;
localparam USER_OFFSET  = TID_OFFSET  + TID_WIDTH;
localparam WIDTH        = USER_OFFSET + USER_WIDTH;


/////////////////////////////////////////////////////for axi_lite/////////////////////////////////////////
//write addr channel

//axi_lite reg
//FIFO threshold setting
reg [ADDR_WIDTH-1:0] TH_reg; //offset0, bit3:0
wire axi_awvalid_in;
wire axi_wvalid_in;
wire axi_awready_out;
wire axi_wready_out;

assign axi_awvalid_in = axi_awvalid && cc_as_enable;
assign axi_awready = axi_awready_out;
//write data channel
assign axi_wvalid_in = axi_wvalid && cc_as_enable;
assign axi_wready = axi_wready_out;
// if both axi_awvalid_in=1 and axi_wvalid_in=1 then output axi_awready_out = 1 and axi_wready_out = 1
assign axi_awready_out = (axi_awvalid_in && axi_wvalid_in) ? 1'b1 : 1'b0;
assign axi_wready_out = (axi_awvalid_in && axi_wvalid_in) ? 1'b1 : 1'b0;
//write register
always @(posedge axis_clk or negedge axi_reset_n)  begin
	if ( !axi_reset_n ) begin
		TH_reg <= 4'h6;
	end
	else begin
		if ( axi_awvalid_in && axi_wvalid_in ) begin		//when axi_awvalid_in=1 and axi_wvalid_in=1 means axi_awready_out=1 and axi_wready_out=1
			if (axi_awaddr[11:2] == 10'h000 && (axi_wstrb[0] == 1) ) begin //offset 0 //axi_awaddr is DW address
				TH_reg <= axi_wdata[3:0];
			end
			else begin
				TH_reg <= TH_reg;
			end
		end
	end
end
//axis_switch always output axi_arready = 1 and don't care the axi_arvalid & axi_araddr
//axis_switch only support 1 register bits in offset 0. config read other address offset is reserved.
assign axi_arready = 1;
// axis_switch  always output axi_rvalid = 1 and axi_rdata =  { 28'b0, TH_reg}
assign axi_rvalid = 1;
assign axi_rdata =  { 28'b0, TH_reg };

/////////////////////////////////////////////////////////////////////////////////////////////////////////




//////////////////////////////////////////////////Upstream///////////////////////////////////////////
//For Arbiter
wire [N-1:0]                req, hi_req;
wire  [N-1:0]                grant;


reg [pDATA_WIDTH-1:0]       m_axis_tdata_reg;

	reg [pUSER_PROJECT_SIDEBAND_WIDTH-1:0]     m_axis_tupsb_reg;

reg [pDATA_WIDTH/8-1:0]     m_axis_tstrb_reg;
reg [pDATA_WIDTH/8-1:0]     m_axis_tkeep_reg; 
reg                         m_axis_tlast_reg;        
reg                         m_axis_tvalid_reg;
reg [USER_WIDTH-1:0]        m_axis_tuser_reg;     
reg [TID_WIDTH-1:0]         m_axis_tid_reg;






//for Abiter
assign  req[0] = up_as_tvalid & req_mask[0];
assign  req[1] = aa_as_tvalid & req_mask[1];
assign  req[2] = la_as_tvalid & req_mask[2];
assign  hi_req[0] = up_hpri_req & hi_req_mask[0];
assign  hi_req[1] = hi_req_mask[1];
assign  hi_req[2] = la_hpri_req & hi_req_mask[2];
assign  as_is_tdata     = m_axis_tdata_reg;

	assign  as_is_tupsb     = m_axis_tupsb_reg;

assign  as_is_tstrb     = m_axis_tstrb_reg;
assign  as_is_tkeep     = m_axis_tkeep_reg; 
assign  as_is_tlast     = m_axis_tlast_reg;        
assign  as_is_tvalid    = m_axis_tvalid_reg;
assign  as_is_tuser     = m_axis_tuser_reg;   
assign  as_is_tid       = m_axis_tid_reg;
assign  as_up_tready = grant[0] && is_as_tready;    
assign  as_aa_tready = grant[1] && is_as_tready;
assign  as_la_tready = grant[2] && is_as_tready;    

 

always @(*) begin
  case (grant)
    3'b001: begin   					// For UP 
        m_axis_tdata_reg  = up_as_tdata;

        m_axis_tupsb_reg  = up_as_tupsb;

        m_axis_tstrb_reg  = up_as_tstrb;
        m_axis_tkeep_reg  = up_as_tkeep;
        m_axis_tvalid_reg = up_as_tvalid; 
        m_axis_tuser_reg  = up_as_tuser;
        m_axis_tid_reg    = 2'b00;  
        m_axis_tlast_reg  = up_as_tlast;  
    end
    3'b010: begin  						// For AA 
        m_axis_tdata_reg  = aa_as_tdata;

        m_axis_tupsb_reg  = 5'b0000_0;

        m_axis_tstrb_reg  = aa_as_tstrb;
        m_axis_tkeep_reg  = aa_as_tkeep;
        m_axis_tvalid_reg = aa_as_tvalid;   
        m_axis_tuser_reg  = aa_as_tuser;
        m_axis_tid_reg    = 2'b01; 
        m_axis_tlast_reg  = aa_as_tlast;              
    end	
    3'b100: begin  						// For LA 
        m_axis_tdata_reg  = la_as_tdata;

        m_axis_tupsb_reg  = 5'b0000_0;

        m_axis_tstrb_reg  = la_as_tstrb;
        m_axis_tkeep_reg  = la_as_tkeep;	
        m_axis_tvalid_reg = la_as_tvalid; 
        m_axis_tuser_reg  = la_as_tuser;
        m_axis_tid_reg    = 2'b10; 
        m_axis_tlast_reg  = la_as_tlast;    
    end
    default: begin
        m_axis_tdata_reg  = 32'h0000_0000;

        m_axis_tupsb_reg  = 5'b0000_0;

        m_axis_tstrb_reg  = 4'b0000;
        m_axis_tkeep_reg  = 4'b0000;
        m_axis_tvalid_reg = 1'b0;
        m_axis_tuser_reg  = 2'b00;
        m_axis_tid_reg    = 2'b00; 
        m_axis_tlast_reg  = 0;           
    end
  endcase  
end


reg [2:0] cnt;
//////////  counter for arbiter ack ///////////

always @(posedge axis_clk or negedge axi_reset_n)  begin
	if ( !axi_reset_n ) begin
	    cnt <= 3'b000;
	end
	else begin
		if ( grant!=3'b000 & (grant&hi_req)==3'b000 ) begin	// when grant is not in the hi_req state, after trransfer cnt+1.	
            if(as_is_tvalid & is_as_tready)  cnt<=cnt+1;
            else cnt<=cnt;      
		end
        else 
        cnt <= 3'b000;
	end
end

wire last;
assign last=(as_is_tvalid & is_as_tready & as_is_tlast)|cnt==3'b111;
reg [N:0]grant_next;
reg [N:0]grant_reg;
localparam WAIT_0 = 4'b0001, WAIT_1 = 4'b0010, WAIT_2 = 4'b0100, GRANT_0=4'b1001, GRANT_1=4'b1010, GRANT_2=4'b1100;

assign grant=(grant_reg[3])?grant_reg[2:0]:0;
always @* begin
    case(grant_reg)
    WAIT_0:begin 
        if(hi_req[1]) grant_next=GRANT_1;
        else if (hi_req[2]) grant_next=GRANT_2;
        else if (hi_req[0]) grant_next=GRANT_0;
        else if (req[1])grant_next=GRANT_1;
        else if (req[2])grant_next=GRANT_2;
        else if (req[0])grant_next=GRANT_0;
        else grant_next=grant_reg;
    end

    WAIT_1:begin 
        if(hi_req[2]) grant_next=GRANT_2;
        else if (hi_req[0]) grant_next=GRANT_0;
        else if (hi_req[1]) grant_next=GRANT_1;
        else if (req[2])grant_next=GRANT_2;
        else if (req[0])grant_next=GRANT_0;
        else if (req[1])grant_next=GRANT_1;
        else grant_next=grant_reg;
    end

    WAIT_2:begin 
        if(hi_req[0]) grant_next=GRANT_0;
        else if (hi_req[1]) grant_next=GRANT_1;
        else if (hi_req[2]) grant_next=GRANT_2;
        else if (req[0])grant_next=GRANT_0;
        else if (req[1])grant_next=GRANT_1;
        else if (req[2])grant_next=GRANT_2;
        else grant_next=grant_reg;
    end

    GRANT_0:begin
        if(last) grant_next=WAIT_0;
        else grant_next=grant_reg;
    end

    GRANT_1:begin
        if(last) grant_next=WAIT_1;
        else grant_next=grant_reg;
    end
    GRANT_2:begin
        if(last) grant_next=WAIT_2;
        else grant_next=grant_reg;
    end
    default: begin
             grant_next=grant_reg;
    end
    endcase
end

always @(posedge axis_clk or negedge axi_reset_n) begin
    if (!axi_reset_n)begin 
        grant_reg<=WAIT_0;
    end
    else begin
        grant_reg<=grant_next;
    end
end 



/////////////////////////////////// Downstream//////////////////////////////////////////////////
wire D_m_axis_tvalid; // Downstream master axis tvalid
wire D_m_axis_tready; // Downstream master axis tready
wire [WIDTH-1:0] s_axis; // slave from is.
wire [WIDTH-1:0] m_axis;
generate
    assign s_axis[pDATA_WIDTH-1:0]                  = is_as_tdata;

		assign s_axis[UPSB_OFFSET +: pUSER_PROJECT_SIDEBAND_WIDTH]     = is_as_tupsb;

    assign s_axis[STRB_OFFSET +: pDATA_WIDTH/8]     = is_as_tstrb;
    assign s_axis[KEEP_OFFSET +: pDATA_WIDTH/8]     = is_as_tkeep;
    assign s_axis[LAST_OFFSET]                      = is_as_tlast;
    assign s_axis[TID_OFFSET   +: TID_WIDTH]        = is_as_tid;
    assign s_axis[USER_OFFSET +: USER_WIDTH]        = is_as_tuser;
endgenerate




assign D_m_axis_tready=(as_up_tvalid && up_as_tready) | (as_aa_tvalid && aa_as_tready);

assign as_up_tvalid =(m_axis[TID_OFFSET +: TID_WIDTH]==2'b00) && D_m_axis_tvalid; 
assign as_up_tdata = (m_axis[TID_OFFSET +: TID_WIDTH]==2'b00) ? m_axis[pDATA_WIDTH - 1:0]: 0;

assign as_up_tupsb = (m_axis[TID_OFFSET +: TID_WIDTH]==2'b00) ? m_axis[UPSB_OFFSET +: pUSER_PROJECT_SIDEBAND_WIDTH]: 0;

assign as_up_tstrb = (m_axis[TID_OFFSET +: TID_WIDTH]==2'b00) ? m_axis[STRB_OFFSET +: pDATA_WIDTH/8]: 0;
assign as_up_tkeep = (m_axis[TID_OFFSET +: TID_WIDTH]==2'b00) ? m_axis[KEEP_OFFSET +: pDATA_WIDTH/8]: 0;
assign as_up_tlast = (m_axis[TID_OFFSET +: TID_WIDTH]==2'b00) ? m_axis[LAST_OFFSET]: 0;
assign as_up_tuser = (m_axis[TID_OFFSET +: TID_WIDTH]==2'b00) ? m_axis[USER_OFFSET +: USER_WIDTH]: 0;


assign as_aa_tvalid =(m_axis[TID_OFFSET +: TID_WIDTH]==2'b01) && D_m_axis_tvalid;
assign as_aa_tdata = (m_axis[TID_OFFSET +: TID_WIDTH]==2'b01) ? m_axis[pDATA_WIDTH-1:0]: 0;
assign as_aa_tstrb = (m_axis[TID_OFFSET +: TID_WIDTH]==2'b01) ? m_axis[STRB_OFFSET +: pDATA_WIDTH/8]: 0;
assign as_aa_tkeep = (m_axis[TID_OFFSET +: TID_WIDTH]==2'b01) ? m_axis[KEEP_OFFSET +: pDATA_WIDTH/8]: 0;
assign as_aa_tlast = (m_axis[TID_OFFSET +: TID_WIDTH]==2'b01) ? m_axis[LAST_OFFSET]: 0;
assign as_aa_tuser = (m_axis[TID_OFFSET +: TID_WIDTH]==2'b01) ? m_axis[USER_OFFSET +: USER_WIDTH]: 0;



    localparam fifo_depth=16;
    localparam sram_datawidth=100;

    wire sram_we;
    wire [$clog2(fifo_depth)-1:0] sram_addr;
    wire [sram_datawidth-1:0]sram_din;
    wire [sram_datawidth-1:0] sram_dout;

    fifo #(.WIDTH(WIDTH),.depth(fifo_depth),.sram_datawidth(sram_datawidth),.mode(1)) as_fifo
    (
        .axis_clk(axis_clk),
        .axi_reset_n(axi_reset_n),
        .w_vld(is_as_tvalid),
        .w_rdy(as_is_tready),
        .data_in(s_axis),
        .r_vld(D_m_axis_tvalid),
        .r_rdy(D_m_axis_tready),
        .data_out(m_axis),
        .TH_reg({4'd0,TH_reg}),
        .sram_we(sram_we),
        .sram_addr(sram_addr),
        .sram_din(sram_din),
        .sram_dout(sram_dout)
    );

    ra1shd16x100m4h3v2 AS_SRAM16x100(
        .CLK(axis_clk),
        .WEN(~sram_we),
        .OEN(1'b0),
        .CEN(1'b0),
        .A(sram_addr),
        .D(sram_din),
        .Q(sram_dout)
    );


endmodule
`timescale 1 ns / 1 ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/15/2023 10:02:45 AM
// Design Name: 
// Module Name: LOGIC_ANLZ
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// Function Description:
//   - Monitor signals provided by user project. Support up to 24 monitoring signals
//   - Support signal conditioning to trigger signal logging  (Currently, done by host program)
//   - Compress (Waveform compression, e.g. Run-Length-Encoding RLE) the logged signals and sent them to remote users using the Axis port. Waveform can be displayed in remote environments.
//   - Waveform log is designed to be saved in .vcd file format, it can be open by gtkwave.


module LOGIC_ANLZ #( parameter pADDR_WIDTH   = 15,
                     parameter pDATA_WIDTH   = 32
                   )
(
    //AxiLite
    output wire           axi_awready,
    output wire           axi_wready,
    output wire           axi_arready,
    output wire   [31: 0] axi_rdata,
    output wire           axi_rvalid,

    input  wire           axi_awvalid,
    input  wire   [14: 0] axi_awaddr,
    input  wire           axi_wvalid,
    input  wire   [31: 0] axi_wdata,
    input  wire   [3: 0]  axi_wstrb,
    input  wire           axi_arvalid,
    input  wire   [14: 0] axi_araddr,
    input  wire           axi_rready,
    input  wire           cc_la_enable,
    // input  wire           enable_la,     // Jiin : it is internal configuration register

    //AxiS  
    output wire   [31: 0] m_tdata,
    output wire   [3: 0]  m_tstrb,
    output wire   [3: 0]  m_tkeep,
    output wire           m_tlast,
    output wire           m_tvalid,
    output wire   [1: 0]  m_tuser,
    output wire           la_hpri_req,
    input  wire           m_tready,

    //User singals
    input  wire   [23: 0] up_la_data,

    //Generic
    input  wire           user_clock2,
    input  wire           axi_clk,
    input  wire           axi_reset_n,
    input  wire           axis_clk,
    input  wire           uck2_rst_n,
    input  wire           axis_rst_n
);
    localparam FIFO_DEPTH               = 32;  
    localparam AXIS_PKT_LEN             = 8; 
    localparam H_THRESH_DEFAULT         = 7'h40;
    localparam L_THRESH_DEFAULT         = 7'b10; 	

wire trace_push_ok;
reg [23:0] la_enable;
reg [6:0] h_thresh;
reg [6:0] l_thresh;
reg [6:0] pop_cond;
reg enable_la;              // Jiin configuratin register at 'h10  - it is used to reset enable_la
reg [7:0] rc_count;
reg [23:0] r_la_data;       // latched up_la_data;
wire la_change;             // la signal changed       
wire trace_push;            // trace is push into FIFO
wire fifo_full;
wire [31:0] trace_packet;
reg [7:0] fifo_count;       // Jiin: parameterize the size of fifo_count with FIFO_depth use $clog2
reg [7:0] tx_count;         // count # of transfer
reg la_hpri_req_o;


assign axi_awready  = axi_awvalid & axi_wvalid;
assign axi_wready   = axi_awvalid & axi_wvalid;

// axilite read - axi_rdata can be available when axi_arvalid (axi_araddr) is valid

assign axi_rvalid   = axi_arvalid;
assign axi_rdata    = (axi_araddr[11:2] == 10'h000) ? {8'b0, la_enable} :   
                      (axi_araddr[11:2] == 10'h001) ? {25'b0, h_thresh} :       // @'h4
                      (axi_araddr[11:2] == 10'h002) ? {25'b0, l_thresh} :       // @'h8
                      (axi_araddr[11:2] == 10'h003) ? {25'b0, pop_cond} :       // @'hc
                      (axi_araddr[11:2] == 10'h004) ? {31'b0, enable_la} : 32'hFFFFFFFF;  // Jiin @'h10
assign axi_arready  = axi_arvalid;

// Jiin : enable_la is the internal configuration register, we can not use enable_la to reset configuration register
//   use axi_reset_n instead
always @ ( posedge axi_clk or negedge axi_reset_n ) begin
    if( !axi_reset_n) begin
        la_enable   <= 24'h0;
        h_thresh    <= H_THRESH_DEFAULT;
        l_thresh    <= L_THRESH_DEFAULT;
        pop_cond    <= AXIS_PKT_LEN;
        enable_la   <= 1'b0;
    end 
    else if( cc_la_enable & axi_awvalid & axi_wvalid) begin
        if( axi_awaddr[11:2] == 10'h000) la_enable <= axi_wdata[23:0];
        if( axi_awaddr[11:2] == 10'h001) h_thresh  <= axi_wdata[6:0];
        if( axi_awaddr[11:2] == 10'h002) l_thresh  <= axi_wdata[6:0];
        if( axi_awaddr[11:2] == 10'h003) pop_cond  <= axi_wdata[6:0];
        if( axi_awaddr[11:2] == 10'h004) enable_la <= axi_wdata[0];         // Jiin: add configuration : enable_la
    end
end

assign la_change = |(la_enable & ( up_la_data != r_la_data)); 

// fifo full handling
//  - push null-packet all 0
//  - flush FIFO 
//  - restart - 
// issue: when fifo_full, do we still count rc?
// - rc continues count
// - signal waveform recovery
//   - when receive null-packet -> generate a cycle of 'x' signals
//   - generate signal waveforms with non-null packet with rc 


always @ ( posedge axi_clk or negedge enable_la) begin  // note: cc_la_enable to reset
    if( !enable_la ) begin
        rc_count  <= 8'h01;
        r_la_data <= 24'b0;
    end 
    else begin
        if( !la_change & rc_count != 8'hff)             // signal is not changed
            rc_count <= rc_count + 1;
        else begin
            r_la_data <= up_la_data;
            rc_count <= 8'h01;
        end
    end 
end


// trace_push : condition to push a trace into fifo
// 1. signal changes - la_change
// 2. rc_count reach 255
// 3. fifo_full -> push null packet (issue : use fifo_full - 1 or fifo_count == l_thread)

// --- FIFO Instance -----



    localparam sram_datawidth=64;

    wire sram_we;
    wire [$clog2(FIFO_DEPTH)-1:0] sram_addr;
    wire [sram_datawidth-1:0]sram_din;
    wire [sram_datawidth-1:0] sram_dout;

// --- FIFO Instance -----
fifo #(.WIDTH(32),.depth(FIFO_DEPTH),.sram_datawidth(sram_datawidth),.mode(0)) la_fifo
(
    .axis_clk (axis_clk) ,
    .axi_reset_n (enable_la),
    .w_vld (trace_push),          // fifo push
    .w_rdy (trace_push_ok),          // w_rdy
    .data_in (trace_packet),
    .r_rdy (m_tready),          // directly connect to axis r_ready
    .r_vld (m_tvalid),          // connect to axis r_valid
    .data_out (m_tdata),
    .TH_reg(8'd0),
    .sram_we(sram_we),
    .sram_addr(sram_addr),
    .sram_din(sram_din),
    .sram_dout(sram_dout)
);



    ra1shd32x64m4h3v2 la_SRAM32x64(
        .CLK(axis_clk),
        .WEN(~sram_we),// WEB =1 is read WEB=0 is w_vldite
        .OEN(1'b0),
        .CEN(1'b0),
        .A(sram_addr),
        .D(sram_din),
        .Q(sram_dout)
    );


// fifo pop & fifo push , m_tvalid is the fifo_empty , trace_push_ok is the fifo_full - JIANG
wire fifo_pop = m_tready & m_tvalid;
wire fifo_push = trace_push & trace_push_ok;

//  FIFO depth counter - it is used to asserts la_hpri_req
//  Jiin: explain the trace push logic
//  push condition
//  1. signal change: la_change
//  2. rc (repeat-count) reach maximum, i.e. rc = 8'hff
//  3. fifo_full_push - fifo_full & push (null_pakcet) - JIANG
//      r_block_push - block fifo push when fifo full
//      from fifo_full -> la_hpri_req_o (change to 1)
//      at the end of the r_block_push, push a null-packet (use la_hpri_req_o and r_block_push) - JIANG
//      from fifo_full -> la_hpri_req_o (change to 0)

reg r_block_push; 
wire fifo_full_push;

always @ ( posedge axi_clk or negedge enable_la )begin
      if(!enable_la) begin
        r_block_push <= 0;
      end 
      else if( trace_push_ok == 1'b0) r_block_push <= 1;
      else if( la_hpri_req_o == 1'b0) r_block_push <= 0; // delay one cycle(from fifo_count < l_thresh) - JIANG
    end

assign fifo_full_push = ((r_block_push == 1'b1) & (la_hpri_req_o == 1'b0)); // (fifo_full_push == 1'b0 & (la_hpri_req_o == 1'b1) the end of r_block_push
assign trace_push = ((la_change | (rc_count == 8'hff)) & !r_block_push)  | fifo_full_push; 

assign trace_packet = {32{!fifo_full_push}} & {rc_count, (r_la_data & la_enable)}; 

assign la_hpri_req = la_hpri_req_o;
  always @ ( posedge axi_clk or negedge enable_la ) begin
    if(!enable_la) begin
        fifo_count <= 8'b0;
        la_hpri_req_o <= 0; 
    end
    else begin
        // if(fifo_full) la_hpri_req_o <= 1 ;
        if(fifo_count >= h_thresh)  la_hpri_req_o <= 1;
        if(fifo_count < l_thresh) la_hpri_req_o <= 0;
        if( fifo_push & !fifo_pop) fifo_count <= fifo_count + 1;
        if(!fifo_push &  fifo_pop) fifo_count <= fifo_count - 1;
    end
  end
assign m_tuser = 2'b00;
assign m_tstrb = 4'b1111;
assign m_tkeep = 4'b1111;
assign m_tlast = (tx_count == pop_cond);
//assign m_tvalid = fifo_count > 0;

// m_tlast 
// 1. transfer count reaches AXIS_PKT_LEN - 1
// 2. reach repeat count = 255, then flush it out - this is to avoid staff un-issued traces
// 3. fifo empty 
// Check upstream Axi-switch will still transfer data when there is no tlast

  always @ ( posedge axi_clk or negedge enable_la ) begin 
    if( !enable_la ) 
        tx_count <= 1;
       else begin 
        if(tx_count == pop_cond)
            tx_count <= 1;
        else if(fifo_pop)
            tx_count <= tx_count + 1;
       end
    end
// ----    Jiin - comment out the following
endmodule
`timescale 1 ns / 1 ps

module CFG_CTRL #( parameter pADDR_WIDTH   = 12,
                   parameter pDATA_WIDTH   = 32
                 )
(
	//////////////////////////////////////
	// FPGA AXI-Lite, from Axis-Axilite //
	//////////////////////////////////////
	input  wire          aa_cfg_awvalid,
	input  wire  [31: 0] aa_cfg_awaddr,
	input  wire          aa_cfg_wvalid,
	input  wire  [31: 0] aa_cfg_wdata,
	input  wire   [3: 0] aa_cfg_wstrb,
	input  wire          aa_cfg_arvalid,
	input  wire  [31: 0] aa_cfg_araddr,
	input  wire          aa_cfg_rready,
	output wire  [31: 0] aa_cfg_rdata,
	output wire          aa_cfg_rvalid,
	output wire          aa_cfg_awready,
	output wire          aa_cfg_wready,
	output wire          aa_cfg_arready,
	
	/////////////////////
	// AXI-Lite Master //
	/////////////////////
	input  wire          axi_wready1,		//for AXIL_AXIS
	input  wire          axi_awready1,
	input  wire          axi_arready1,
	input  wire  [31: 0] axi_rdata1,
	input  wire          axi_rvalid1,
	input  wire          axi_awready4,		//for AXIL_SWITCH
	input  wire          axi_wready4,
	input  wire          axi_arready4,
	input  wire  [31: 0] axi_rdata4,
	input  wire          axi_rvalid4,
	input  wire          axi_awready3,		//for IO_SERDES
	input  wire          axi_wready3,
	input  wire          axi_arready3,
	input  wire  [31: 0] axi_rdata3,
	input  wire          axi_rvalid3,
	input  wire          axi_awready0,		//for LOGIC_ANLZ
	input  wire          axi_wready0,
	input  wire          axi_arready0,
	input  wire  [31: 0] axi_rdata0,
	input  wire          axi_rvalid0,
	input  wire          axi_awready2,		//for USERSUBSYS
	input  wire          axi_wready2,
	input  wire          axi_arready2,
	input  wire  [31: 0] axi_rdata2,
	input  wire          axi_rvalid2,
	output wire          axi_awvalid,
	output wire  [14: 0] axi_awaddr,
	output wire          axi_wvalid,
	output wire  [31: 0] axi_wdata,
	output wire   [3: 0] axi_wstrb,
	output wire          axi_arvalid,
	output wire  [14: 0] axi_araddr,
	output wire          axi_rready,	
	
	//////////////////////
	// Target Selection //
	//////////////////////
	output wire          cc_aa_enable,
	output wire          cc_as_enable,
	output wire          cc_is_enable,
	output wire          cc_la_enable,
	output wire          cc_up_enable,
	output wire   [4: 0] user_prj_sel,
	
	////////////////////////
	// Wishbone interface //
	////////////////////////	
	input  wire          wb_rst,
	input  wire          wb_clk,
	input  wire  [31: 0] wbs_adr,
	input  wire  [31: 0] wbs_wdata,
	input  wire   [3: 0] wbs_sel,
	input  wire          wbs_cyc,
	input  wire          wbs_stb,
	input  wire          wbs_we,
	output wire          wbs_ack,
	output wire  [31: 0] wbs_rdata,
	
	//////////////////////////
	// Top AXI-Lite Signals //
	//////////////////////////
	input  wire          user_clock2,
	input  wire          axi_clk,
	input  wire          axi_reset_n,
	input  wire          uck2_rst_n
);

	////////////////////////////
	// Internal Signals begin //
	////////////////////////////	
	reg wb_fsm_reg;
	reg wb_axi_request;
	reg wb_axi_request_rw;
	reg [3:0] wb_axi_wstrb;
	reg wb_axi_request_done;
	reg [31:0] wb_axi_request_add;
	reg [31:0] wb_axi_wdata;
	reg [31:0] wb_axi_rdata;
	
	reg [2:0] f_axi_fsm_reg;
	reg f_axi_request;
	reg f_axi_request_rw;
	reg [3:0] f_axi_wstrb;
	reg f_axi_request_done;
	reg [31:0] f_axi_request_add;
	reg [31:0] f_axi_wdata;
	reg [31:0] f_axi_rdata;
	
	reg [2:0] m_axi_fsm_reg;
	
	reg axi_grant_o_reg;
	wire m_axi_request;
	wire m_axi_request_rw;
	wire [3:0] m_axi_wstrb;
	wire m_axi_request_done;
	wire [31:0] m_axi_request_add;
	wire [31:0] m_axi_wdata;
	
	wire m_axi_awready;
	wire m_axi_wready;
	wire m_axi_arready;
	wire [31:0] m_axi_rdata;
	wire m_axi_rvalid;
	
	reg cc_enable;
	reg cc_sub_enable;

	wire cc_axi_awvalid;
	wire cc_axi_wvalid;

	reg [2:0] cc_s_fsm_reg;	
	reg [11:0] cc_s_addr;
	reg [31:0] cc_s_wdata;
	reg [31:0] cc_s_rdata;
	
	wire axi_awready5;
	wire axi_wready5;
	wire axi_arready5;
	wire [31: 0] axi_rdata5;
	wire axi_rvalid5;
	
	//////////////////////////////////////
	// Internal signals for Ports begin //
	//////////////////////////////////////
	reg [31:0] aa_cfg_rdata_o;
	reg aa_cfg_rvalid_o;
	reg aa_cfg_awready_o;
	reg aa_cfg_wready_o;
	reg aa_cfg_arready_o;
	
	reg axi_awvalid_o;
	reg [14:0] axi_awaddr_o;
	reg axi_wvalid_o;
	reg [31:0] axi_wdata_o;
	reg [3:0] axi_wstrb_o;
	reg axi_arvalid_o;
	reg [14:0] axi_araddr_o;
	reg axi_rready_o;

	reg cc_aa_enable_o;
	reg cc_as_enable_o;
	reg cc_is_enable_o;
	reg cc_la_enable_o;
	reg cc_up_enable_o;

	reg [4: 0] user_prj_sel_o;
	
	reg wbs_ack_o;
	reg [31: 0] wbs_rdata_o;
	
	///////////////////////////////////
	// Assignment for Internal begin //
	///////////////////////////////////
	assign m_axi_request = axi_grant_o_reg ? f_axi_request : wb_axi_request;
	assign m_axi_request_rw = axi_grant_o_reg ? f_axi_request_rw : wb_axi_request_rw;
	assign m_axi_wstrb = axi_grant_o_reg ? f_axi_wstrb : wb_axi_wstrb;
	assign m_axi_request_done = axi_grant_o_reg ? f_axi_request_done : wb_axi_request_done;
	assign m_axi_request_add = axi_grant_o_reg ? f_axi_request_add : wb_axi_request_add;
	assign m_axi_wdata = axi_grant_o_reg ? f_axi_wdata : wb_axi_wdata;

	/*
	In case of cc_sub_enable, read always return 0xFFFFFFFF, write always complete.
	({1{cc_sub_enable}} & axi_awvalid))
	({1{cc_sub_enable}} & axi_wvalid))
	({1{cc_sub_enable}} & axi_arvalid))
	({32{cc_sub_enable}} & 32'hFFFFFFFF))
	({1{cc_sub_enable}} & axi_arvalid))
	*/
	assign m_axi_awready = ((((((({1{cc_up_enable}} & axi_awready2) | ({1{cc_la_enable}} & axi_awready0)) | ({1{cc_aa_enable}} & axi_awready1)) | ({1{cc_is_enable}} & axi_awready3)) | ({1{cc_as_enable}} & axi_awready4)) | ({1{cc_enable}} & axi_awready5)) | ({1{cc_sub_enable}} & axi_awvalid));
	assign m_axi_wready = ((((((({1{cc_up_enable}} & axi_wready2) | ({1{cc_la_enable}} & axi_wready0)) | ({1{cc_aa_enable}} & axi_wready1)) | ({1{cc_is_enable}} & axi_wready3)) | ({1{cc_as_enable}} & axi_wready4)) | ({1{cc_enable}} & axi_wready5)) | ({1{cc_sub_enable}} & axi_wvalid));
	assign m_axi_arready = ((((((({1{cc_up_enable}} & axi_arready2) | ({1{cc_la_enable}} & axi_arready0)) | ({1{cc_aa_enable}} & axi_arready1)) | ({1{cc_is_enable}} & axi_arready3)) | ({1{cc_as_enable}} & axi_arready4)) | ({1{cc_enable}} & axi_arready5)) | ({1{cc_sub_enable}} & axi_arvalid));
	assign m_axi_rdata = ((((((({32{cc_up_enable}} & axi_rdata2) | ({32{cc_la_enable}} & axi_rdata0)) | ({32{cc_aa_enable}} & axi_rdata1)) | ({32{cc_is_enable}} & axi_rdata3)) | ({32{cc_as_enable}} & axi_rdata4)) | ({32{cc_enable}} & axi_rdata5)) | ({32{cc_sub_enable}} & 32'hFFFFFFFF));
	assign m_axi_rvalid = ((((((({1{cc_up_enable}} & axi_rvalid2) | ({1{cc_la_enable}} & axi_rvalid0)) | ({1{cc_aa_enable}} & axi_rvalid1)) | ({1{cc_is_enable}} & axi_rvalid3)) | ({1{cc_as_enable}} & axi_rvalid4)) | ({1{cc_enable}} & axi_rvalid5)) | ({1{cc_sub_enable}} & axi_arvalid));
	
	
	assign cc_axi_awvalid = axi_awvalid && cc_enable;
	assign cc_axi_wvalid = axi_wvalid && cc_enable;

	////////////////////////////////
	// Assignment for Ports begin //
	////////////////////////////////
	assign aa_cfg_rdata = aa_cfg_rdata_o;
	assign aa_cfg_rvalid = aa_cfg_rvalid_o;
	assign aa_cfg_awready = aa_cfg_awready_o;
	assign aa_cfg_wready = aa_cfg_wready_o;
	assign aa_cfg_arready = aa_cfg_arready_o;

	assign axi_awvalid = axi_awvalid_o;
	assign axi_awaddr = axi_awaddr_o;
	assign axi_wvalid = axi_wvalid_o;
	assign axi_wdata = axi_wdata_o;
	assign axi_wstrb = axi_wstrb_o;
	assign axi_arvalid = axi_arvalid_o;
	assign axi_araddr = axi_araddr_o;
	assign axi_rready = axi_rready_o;

	assign cc_aa_enable = cc_aa_enable_o;
	assign cc_as_enable = cc_as_enable_o;
	assign cc_is_enable = cc_is_enable_o;
	assign cc_la_enable = cc_la_enable_o;
	assign cc_up_enable = cc_up_enable_o;

	assign user_prj_sel = user_prj_sel_o;

	assign wbs_ack = wbs_ack_o;
	assign wbs_rdata = wbs_rdata_o;

	assign axi_awready5 = cc_axi_awvalid ? 1 : 0;
	assign axi_wready5 = cc_axi_wvalid ? 1 : 0;
	assign axi_arready5 = 1'b1;
	assign axi_rdata5 = { 27'b0, user_prj_sel_o };
	assign axi_rvalid5 = 1'b1;

	//////////////////////////// 
	// Local paramaters begin //
	////////////////////////////
	localparam wb_fsm_idle = 1'b0;
	localparam wb_fsm_inprogress = 1'b1;

	localparam axi_fsm_idle = 3'b000;
	localparam axi_fsm_read_data = 3'b001;
	localparam axi_fsm_read_complete = 3'b010;
	localparam axi_fsm_write_data = 3'b011;
	localparam axi_fsm_write_complete = 3'b100;
	
	/////////////////////////////////
	// Always for Target Selection //
	/////////////////////////////////
	always @ ( posedge axi_clk or negedge axi_reset_n)
	begin
		if ( !axi_reset_n )
		begin
			cc_aa_enable_o <= 1'b0;
			cc_as_enable_o <= 1'b0;
			cc_is_enable_o <= 1'b0;
			cc_la_enable_o <= 1'b0;
			cc_up_enable_o <= 1'b0;
			cc_enable <= 1'b0;
			cc_sub_enable <= 1'b0;
		end else
		begin
			cc_aa_enable_o <= ( m_axi_request_add[31:12] == 20'h30002 )? 1'b1 : 1'b0;
			cc_as_enable_o <= ( m_axi_request_add[31:12] == 20'h30004 )? 1'b1 : 1'b0;
			cc_is_enable_o <= ( m_axi_request_add[31:12] == 20'h30003 )? 1'b1 : 1'b0;
			cc_la_enable_o <= ( m_axi_request_add[31:12] == 20'h30001 )? 1'b1 : 1'b0;
			cc_up_enable_o <= ( m_axi_request_add[31:12] == 20'h30000 )? 1'b1 : 1'b0;
			cc_enable <= ( m_axi_request_add[31:12] == 20'h30005 )? 1'b1 : 1'b0;
			cc_sub_enable <= ( (m_axi_request_add[31:12] >= 20'h30006) && (m_axi_request_add[31:12] <= 20'h3FFFF ) )? 1'b1 : 1'b0;
		end
	end	
	////////////////////////////////////////////
	// Always for Wishbone Interface handling //
	////////////////////////////////////////////
	always @ ( posedge wb_clk or posedge wb_rst)
	begin
		if ( wb_rst ) 
		begin
			wb_fsm_reg <= wb_fsm_idle;
			wb_axi_request <= 1'b0;
			wb_axi_request_rw <= 1'b0;
			wb_axi_wstrb <= 4'b0;
			wb_axi_request_add <= 32'b0;
			wb_axi_wdata <= 32'b0;
			
			wbs_ack_o <= 1'b0;
			wbs_rdata_o <= 32'b0;						
		end else
		begin
			case (wb_fsm_reg) 
				wb_fsm_idle:
				begin
					wbs_ack_o <= 1'b0;
					wbs_rdata_o <= 32'h0;
					if ( !wbs_ack_o ) begin
						if ( wbs_cyc && wbs_stb ) begin
							wb_axi_request <= 1'b1;
							wb_axi_request_rw <= wbs_we;
							wb_axi_request_add <= wbs_adr;	//Latch wbs_adr
							if ( wbs_we ) begin
								wb_axi_wdata <= wbs_wdata;	//Latch wbs_wdata;
								wb_axi_wstrb <= wbs_sel;
							end
							wb_fsm_reg <= wb_fsm_inprogress;
						end
					end
				end
				wb_fsm_inprogress:
				begin
					if ( wb_axi_request_done )
					begin
						wbs_ack_o <= 1'b1;	
						if ( !wb_axi_request_rw )
							wbs_rdata_o <= wb_axi_rdata;	//Output wbs_rdata_o
						else
							wb_axi_wdata <= 32'h0;
						wb_axi_request <= 1'b0;
						wb_axi_request_add <= 32'b0;
						wb_fsm_reg <= wb_fsm_idle;						
					end
				end
			endcase
		end
	end	

	/////////////////////////////////////////////////
	// Always for FPGA-AXI-Lite Interface handling //
	/////////////////////////////////////////////////	
	always @ ( posedge axi_clk or negedge axi_reset_n)
	begin
		if ( !axi_reset_n )
		begin
			f_axi_fsm_reg <= axi_fsm_idle;
			f_axi_request <= 1'b0;
			f_axi_request_rw <= 1'b0;
			f_axi_wstrb <= 4'b0;
			f_axi_request_add <= 32'b0;
			f_axi_wdata <= 32'b0;
			
			aa_cfg_rdata_o <= 32'b0;
			aa_cfg_rvalid_o <= 1'b0;
			aa_cfg_awready_o <= 1'b0;
			aa_cfg_wready_o <= 1'b0;
			aa_cfg_arready_o <= 1'b0;			
		end else
		begin
			case ( f_axi_fsm_reg )
				axi_fsm_idle:
				begin			
					aa_cfg_wready_o <= 1'b0;
					if ( aa_cfg_awvalid ) begin
						aa_cfg_awready_o <= 1'b1;
						f_axi_request_add <= aa_cfg_awaddr;		//Latch awaddr
						f_axi_fsm_reg <= axi_fsm_write_data;
					end else if ( aa_cfg_arvalid ) begin
						aa_cfg_arready_o <= 1'b1;
						f_axi_request_add <= aa_cfg_araddr;		//Latch araddr
						f_axi_request_rw <= 1'b0;
						f_axi_request <= 1'b1;						
						f_axi_fsm_reg <= axi_fsm_read_data;
					end
				end
				axi_fsm_read_data:
				begin
					aa_cfg_arready_o <= 1'b0;
					if ( aa_cfg_rready && f_axi_request_done ) begin
						aa_cfg_rdata_o <= f_axi_rdata;			//Output aa_cfg_rdata_o
						aa_cfg_rvalid_o <= 1'b1;
						f_axi_request <= 1'b0;	
						f_axi_request_add <= 32'b0;
						f_axi_fsm_reg <= axi_fsm_read_complete;						
					end
				end
				axi_fsm_read_complete:
				begin
					if ( aa_cfg_rready ) begin
						aa_cfg_rdata_o <= 32'b0;
						aa_cfg_rvalid_o <= 1'b0;
						f_axi_fsm_reg <= axi_fsm_idle;		
					end					
				end
				axi_fsm_write_data:
				begin
					aa_cfg_awready_o <= 1'b0;
					if ( aa_cfg_wvalid ) begin
						f_axi_request <= 1'b1;
						f_axi_request_rw <= 1'b1;	
						f_axi_wdata <= aa_cfg_wdata;			//Latch wdata
						f_axi_wstrb <= aa_cfg_wstrb;						
						f_axi_fsm_reg <= axi_fsm_write_complete;		
					end
				end
				axi_fsm_write_complete:
				begin
					if ( f_axi_request_done ) begin
						aa_cfg_wready_o <= 1'b1;
						f_axi_request <= 1'b0;		
						f_axi_request_add <= 32'b0;
						f_axi_fsm_reg <= axi_fsm_idle;								
					end
				end
			endcase			
		end
	end
	
	/////////////////////////////////////////////////
	// Always for requests grant - axi_grant_o_reg //
	/////////////////////////////////////////////////
	always @( posedge wb_clk or posedge wb_rst )
	begin
		if ( wb_rst ) begin
			axi_grant_o_reg <= 1'b0;
		end else begin
			case (axi_grant_o_reg)
				1'b0: begin
					if ((~wb_axi_request)) begin
						if (f_axi_request) begin
							axi_grant_o_reg <= 1'b1;
						end
					end
				end
				1'b1: begin
					if ((~f_axi_request)) begin
						if (wb_axi_request) begin
							axi_grant_o_reg <= 1'b0;
						end
					end
				end			
			endcase
		end
	end		

	///////////////////////////////////////////////////
	// Always for AXI-Lite Master Interface handling //
	///////////////////////////////////////////////////
	always @ ( posedge axi_clk or negedge axi_reset_n )
	begin
		if ( !axi_reset_n ) begin
			wb_axi_rdata <= 32'b0;
			wb_axi_request_done <= 1'b0;
			
			f_axi_rdata <= 32'b0;
			f_axi_request_done <= 1'b0;
			
			axi_awvalid_o <= 1'b0;
			axi_awaddr_o <= 15'b0;
			axi_wvalid_o <= 1'b0;
			axi_wdata_o <= 32'b0;
			axi_wstrb_o <= 4'b0;
			axi_arvalid_o <= 1'b0;
			axi_araddr_o <= 15'b0;
			axi_rready_o <= 1'b0;			

			m_axi_fsm_reg <= axi_fsm_idle;
		end else begin
			case ( m_axi_fsm_reg )
				axi_fsm_idle:
				begin
					wb_axi_request_done <= 1'b0;
					f_axi_request_done <= 1'b0;			
					if ( m_axi_request && !m_axi_request_done ) begin
						if ( m_axi_request_rw ) begin
							axi_awvalid_o <= 1'b1;
							axi_awaddr_o <= m_axi_request_add[14:0];							
							axi_wvalid_o <= 1'b1;
							axi_wdata_o <= m_axi_wdata;
							axi_wstrb_o <= m_axi_wstrb;
							m_axi_fsm_reg <= axi_fsm_write_data;
						end else begin
							axi_arvalid_o <= 1'b1;							
							axi_araddr_o <= m_axi_request_add[14:0];
							axi_rready_o <= 1'b1;
							m_axi_fsm_reg <= axi_fsm_read_data;
						end
					end
				end
				axi_fsm_read_data:
				begin
					if ( m_axi_arready && m_axi_rvalid) begin
						axi_arvalid_o <= 1'b0;
						axi_araddr_o <= 15'b0;
						axi_rready_o <= 1'b0;
						if ( axi_grant_o_reg )
							f_axi_rdata <= m_axi_rdata;
						else 
							wb_axi_rdata <= m_axi_rdata;
						if ( axi_grant_o_reg )
							f_axi_request_done <= 1'b1;
						else 
							wb_axi_request_done <= 1'b1;
						m_axi_fsm_reg <= axi_fsm_idle;												
					end else if ( m_axi_arready ) begin
						axi_araddr_o <= 15'b0;
						axi_arvalid_o <= 1'b0;
						m_axi_fsm_reg <= axi_fsm_read_complete;	
					end
				end
				axi_fsm_read_complete:
				begin
					if ( m_axi_rvalid ) begin
						axi_rready_o <= 1'b0;
						if ( axi_grant_o_reg )
							f_axi_rdata <= m_axi_rdata;
						else 
							wb_axi_rdata <= m_axi_rdata;
						if ( axi_grant_o_reg )
							f_axi_request_done <= 1'b1;
						else 
							wb_axi_request_done <= 1'b1;
						m_axi_fsm_reg <= axi_fsm_idle;						
					end
				end
				axi_fsm_write_data:
				begin
					if ( m_axi_awready && m_axi_wready) begin
						axi_awvalid_o <= 1'b0;
						axi_awaddr_o <= 15'b0;
						axi_wvalid_o <= 1'b0;
						axi_wdata_o <= 32'b0;
						axi_wstrb_o <= 4'b0;
						if ( axi_grant_o_reg )
							f_axi_request_done <= 1'b1;
						else 
							wb_axi_request_done <= 1'b1;						
						m_axi_fsm_reg <= axi_fsm_idle;	
					end	else begin
						if ( m_axi_awready ) begin
							axi_awaddr_o <= 15'b0;
							axi_awvalid_o <= 1'b0;
							m_axi_fsm_reg <= axi_fsm_write_complete;								
						end
					end
				end
				axi_fsm_write_complete:
				begin
					if ( m_axi_wready) begin
						axi_wvalid_o <= 1'b0;
						axi_wdata_o <= 32'b0;
						axi_wstrb_o <= 4'b0;
						if ( axi_grant_o_reg )
							f_axi_request_done <= 1'b1;
						else 
							wb_axi_request_done <= 1'b1;					
						m_axi_fsm_reg <= axi_fsm_idle;	
					end
				end
			endcase
		end
	end

	///////////////////////////////////////////
	// Always for AXI-Lite CC Slave response //
	///////////////////////////////////////////	
	always @ ( posedge axi_clk or negedge axi_reset_n ) 
	begin	
		if ( !axi_reset_n ) begin
			user_prj_sel_o <= 5'b0;
		end else begin
			if ( cc_axi_awvalid && cc_axi_wvalid ) begin
				if (axi_awaddr[11:0] == 12'h000 && (axi_wstrb[0] == 1) ) begin //offset 0
					user_prj_sel_o <= axi_wdata[4:0];
				end
				else begin
					user_prj_sel_o <= user_prj_sel_o;
				end
			end
		end
	end	

endmodule
// AXIL-AXIS (AA module) - AXILite-AXIS Protcol Conversion
//  Specification: https://github.com/bol-edu/fsic_fpga/blob/main/fsic-spec-dev/modules/FSIC-AXIS%20interface%20specification.md
// 
// - Simplify the design, no fifo
//   Assuming there is no pipeline ss->lm transaction
//   Assuming there is no pipeline ls->sm tranaction 
//   Assuming there is no concurrent ss, ls transaction, i.e. either ss, or ls transaction is only, it will stall the other.
// 
// - Support 
//   Axis-slave to Axilite Master (ss->lm -> sm) read/write 
//   Axilite slave to Axis-master (ls -> sm -> ss) read/write
//   mailbox - support on 8 DW register (DW#0 - FSIC, DW#1 - FPGA)
// 

//reg [6:0] ss_lm_fsm;
`define SS_IDLE             7'b0_0_0_0_0_0_0
`define SS_RD               7'b0_1_0_0_0_0_0
`define SS_WR_S1            7'b0_1_1_0_0_0_0
`define SS_WR_S2            7'b0_1_1_0_0_1_0
`define SS_WR_LM            7'b0_0_1_1_0_0_0
`define SS_WR_LM_AW         7'b1_0_1_1_0_0_0
`define SS_RD_LM_AR         7'b0_0_0_1_0_0_0
`define SS_RD_LM_R          7'b0_0_0_1_0_1_0
`define SS_RD_SM_RS         7'b0_0_0_0_1_0_0
`define SS_DONE             7'b0_0_0_0_0_0_1


module AXIL_AXIS #( parameter pADDR_WIDTH   = 12,
                    parameter pDATA_WIDTH   = 32
                  )
(

//for post simulation signal in testbench
  output wire intr_enable_out,

// Clock & Reset - only use axis_clk, axis_rst_n
  input  wire          axi_clk,
  input  wire          axi_reset_n,
  input  wire          axis_clk,
  input  wire          axis_rst_n,

// LM - Axilite Master
// LM AW Channel
  output wire          m_awvalid,
  output wire  [31: 0] m_awaddr,
  input  wire          m_awready,

// LM  W Channel
  output wire          m_wvalid,
  output wire  [31: 0] m_wdata,
  output wire   [3: 0] m_wstrb,    // follow axis 2nd cycle ss_tdata[31:28]
  input  wire          m_wready,

/// LM AR Channel
  output wire          m_arvalid,
  output wire  [31: 0] m_araddr,
  input  wire          m_arready,

// LM R Channel
  output wire          m_rready,
  input  wire          m_rvalid,
  input  wire  [31: 0] m_rdata,


// LS - Axilite Slave
// LS AW Channel
  output wire          s_awready,
  input  wire          s_awvalid,
  input  wire  [14: 0] s_awaddr,

// LS W Channel
  output wire          s_wready,
  input  wire          s_wvalid,
  input  wire  [31: 0] s_wdata,  
  input  wire   [3: 0] s_wstrb,

// LS AR Channel
  output wire          s_arready,
  input  wire          s_arvalid,
  input  wire  [14: 0] s_araddr,

 // LS R Channel
  output wire  [31: 0] s_rdata,
  output wire          s_rvalid,
  input  wire          s_rready,

// -- Stream Interface with Axi-Switch (AS)

// SS - Stream Slave
  input  wire  [31: 0] as_aa_tdata,
  input  wire   [3: 0] as_aa_tstrb,
  input  wire   [3: 0] as_aa_tkeep,
  input  wire          as_aa_tlast,
  input  wire          as_aa_tvalid,
  input  wire   [1: 0] as_aa_tuser,
  output  wire         aa_as_tready,

// SM - Stream Master
  output wire  [31: 0] aa_as_tdata,
  output wire   [3: 0] aa_as_tstrb,
  output wire   [3: 0] aa_as_tkeep,
  output wire          aa_as_tlast,
  output wire          aa_as_tvalid,
  output wire   [1: 0] aa_as_tuser,
  input  wire          as_aa_tready,

// Misc
  input  wire          cc_aa_enable,   // all Axilite Slave transaction should be qualified by cc_aa_enable
  output wire          mb_irq          // Generate interrupt only when mailbox write by remote, i.e. from Axi-stream
 
);
  localparam TUSER_AXIS = 2'b00;
  localparam TUSER_AXILITE_WRITE = 2'b01;
  localparam TUSER_AXILITE_READ_REQ = 2'b10;
  localparam TUSER_AXILITE_READ_CPL = 2'b11;

  localparam TID_DN_UP = 2'b00;
  localparam TID_DN_AA = 2'b01;
  localparam TID_UP_UP = 2'b00;
  localparam TID_UP_AA = 2'b01;
  localparam TID_UP_LA = 2'b10;

// naming rule
// r_   : registered/latched
// _n   : active low
// _cyc : transaction cycle 
// interface ports:
// - ss (stream slave)
// - sm (stream master)
// - ls (axilite slave)
// - lm (axilite master)
// cycle type indicators:
// - wr : write transaction
// - rd : read transaction
// - rs : read response

// aa_reset_n - AA module reset, active low
// 1. system reset
// 2. cc_aa_enable = 0 : if AA is not enable, treated as reset
wire aa_reset_n = axis_rst_n;

// move here for early declaraion before use it to avoid error in simulation
wire ss_sm_cyc;
wire ss_t2;
reg [6:0] ss_lm_fsm;
wire ss_lm_enable;
//
//   SS Cycle type - decode from tuser, refer to fsic-axis specification
//   tuser = 2'b00    - axis cycle, ignored, we don't handle pure axi-stream transaction
//   tuser = 2'b01    - axilite write - 2T  T1:address, T2:data
//   tuser = 2'b10    - axilite read - address
//   tuser = 2'b11    - axilite read - data response
// Note: we should use latched tuser ----
wire ss_axis_cyc    = (as_aa_tuser == 2'b00);    // actually, we won't receive this cycle, as should filter it out
wire ss_wr_cyc      = (as_aa_tuser == 2'b01);    // tready is return as long as address/data latch is ok (ss_w_addr_data_ok)
wire ss_rd_cyc      = (as_aa_tuser == 2'b10);    // tready is return as long as ss_rw_addr latch is ok
wire ss_rs_cyc      = (as_aa_tuser == 2'b11); 


// --------------------------------
// Internal States
// --------------------------------
// Data/Address latches
// As a slave, we will latch (save) address and data used for the master transaction later, example
// SS -> LM  write : latch address (1st T) and data (2nd T)
// SS -> LM  read :  latch address (1st T)
// LS -> SS  write : latch address (@awvalid), data (@wvalid)
// LS -> SS  read : latch address (@arvalid), data @(rready) 
//

// ----------------------------
// cycle tracking  - ss_cyc, ls_cyc
// ----------------------------
// ------  SS -> LM  -----------
//reg  ss_wr;                  // status: latched ss transaction is read(0) or write(1)
//wire ss_rd = ~ss_wr;
wire ss_cyc;                    // indicate there is ss_cyc pending, set by ss, reset by axil transaction complete
//wire lm_ready;                // axil master transaction complete, m_wready(write), m_rvalid(read)
//wire lm_done = lm_ready;    // same as lm_ready
// reg r_ss_rresp;               // ss read data is complete, generate sm response data ??

// LS -> SM
wire ls_wr;                // indicate ls transaction is read(0), write(1)
wire ls_cyc;               // ls cycle is ongoing
                            //   write -> until sm send out stream write
                            //   read  -> until ss receive tuser= 2'b11, read response data
//reg r_sm_done;              // sm write transferred, or sm read address sent
// reg r_ss_axil_rresp;        // r_ss  ??

// ----------------------------------
//  Lached Input address / data from SS, LS, LM (response data)
// ----------------------------------
// --- SS ------------
reg [31:0] r_ss_rw_addr;            // ss-axil address latch for read and write - shared
reg [31:0] r_ss_wdata;             // ss-axil data latch for write, 
                                    //    also used for ss-axil read response data, guarantee exclusive ss w/rs by not responding ss_ready
                                    //    if ss_cyc is on-going, don't asserts ss_tready
                                    // TODO: what happend if ls and ss with valid signal at the same T? add arbitraion for it.
reg [3:0]  r_ss_wstrb;               // ss-axil wstb latch - from SS 1T tdata[31:28]
reg [1:0]  r_tuser;                 // tuser is encoded with cycle type            


// reg [31:0] ss_rs_data;         // ss data for tuser = 2'b11, used as ls respond data, i.e. s_rdata
wire [31:0] ss_rs_data = r_ss_wdata;  // shared, guarantee exclusive ss w/rs by not responding ss_ready, the code may be confusing


// ---  LS -----------  Axilite Slave
// ls side latched address, data, or read data to send
reg [31:0] r_ls_rw_addr;            // ls address

reg [31:0] r_ls_wdata;              // ls write data
reg [3:0]  r_ls_wstrb;              // ls wstrb

// --- LM  ------------ Axilite Master
// lm side - latch read response data
reg [31:0] r_lm_rs_data;            // lm read response data 


// ----------------------------------
//  Module Interface signals - Address/Data to LM, SM from internal latched registers
// ---------------------------------


// ----  LM - Adddress/Data   - from SS latched address/data
assign m_awaddr = r_ss_rw_addr;
assign m_araddr = r_ss_rw_addr;
assign m_wdata  = r_ss_wdata;
assign m_wstrb  = r_ss_wstrb;


// 
// aa_internal - address hit internal aa configuration or mailbox
// From SS
// AA  'h3000_2xxx   r_ss_rw_addr[27:0]
// aa_reg (internal) a[27:0] = 28'h000_21xx
// aa_mbox           a[27:0] = 28'h000_20xx
// From LS
// use r_ls_rw_addr[11:0]
//    aa_reg   12'h1xx
//    aa_mbox  12'h0xx
// 
// From LS
//   - read ( AA, MBOX), Write AA   => no need trigger LS state machine
// From SS
//   - write/read AA  => no need to trigger SS state machine
//   - write Mbox
wire ss_aa_reg  = ( as_aa_tdata[27:8] == 20'h000_21 );   // xxxx_3xxx, xxxx_2xxx only compare addr[11:8];
wire ss_aa_mbox = ( as_aa_tdata[27:8] == 20'h000_20 );  

wire ss_aa_reg_latch = ( r_ss_rw_addr[27:8] == 20'h000_21 );   // xxxx_3xxx, xxxx_2xxx only compare addr[11:8];
wire ss_aa_mbox_latch = ( r_ss_rw_addr[27:8] == 20'h000_20 );  

wire ls_aa_reg  = ( r_ls_rw_addr[14:12] == 3'b010 && r_ls_rw_addr[11:8] == 4'h1);
wire ls_aa_mbox = ( r_ls_rw_addr[14:12] == 3'b010 && r_ls_rw_addr[11:8] == 4'h0 );

wire ls_aa_reg_lw  = ( s_awaddr[14:12] == 3'b010 && s_awaddr[11:8] == 4'h1 );   //ls_aa_reg local write
wire ls_aa_mbox_lw = ( s_awaddr[14:12] == 3'b010 && s_awaddr[11:8] == 4'h0 );   //s_aa_mbox local write

wire ls_aa_reg_lr  = ( s_araddr[14:12] == 3'b010 && s_araddr[11:8] == 4'h1 );   //ls_aa_reg local read
wire ls_aa_mbox_lr = ( s_araddr[14:12] == 3'b010 && s_araddr[11:8] == 4'h0 );   //s_aa_mbox local read

// ---------------------------------------
// AA-register
// - Memory-mapped Address (32'h3000_2000 ~'h3000_2xxx) - cc_aa_enable
    //--------------------------------------------------
    // for AA_REG description
    // offset 0-3 (32bit):
    //   bit 0: Enable Interrupt
    //       0 = disable interrupt signal
    //       1 = enable interrupt signal
    // offset 4-7 (32bit):
    //   bit 0: Interrupt Status
    //       1: interrupt has occurred
    //       0: no interrupt
    //--------------------------------------------------
reg intr_enable;  // rw: offset:0, bit0  - use addr[2] to select
reg intr_status;  // ro: offset:4, bit0
assign intr_enable_out = intr_enable;
// ---------------------------------------
// Mailbox 
// - Memory-mapped address (32'h3000_2000~3000_201f)
//   Use address[4:2]  to index mb_regs
// ---------------------------------------
// parameter MBOX_BASE_  
reg [31:0] mb_regs[7:0];    // only support 8*DW to save space


/// wire [31:0] ss_aa_internal_data;        // ss won't read aa internal data

// for local read - r_ls_rw_addr is valid
wire [31:0] ls_aa_internal_data = ls_aa_reg ? (r_ls_rw_addr[2] ? {31'b0, intr_status}
                                                               : {31'b0, intr_enable})                                             
                                            : mb_regs[r_ls_rw_addr[4:2]];


// for SS read - not verify yet - 
// Question : how to read AA_reg target in remote side? - Limitation
// issue: local_ls read address in AA_reg range will cliam and return locally, do not send to remote side.
//   provide below solution
//   add a input signal named aa_type, AA in soc(0) or fpga(1)
//      for aa_type = soc(0)  then AA_reg in 15'h21xx 
//      for aa_type = fpga(1) then AA_reg in 15'h22xx 
//   for example : 
//         in fpga, ls addr = 15'h21xx for remote AA and send to remote side
//         in fpga, ls addr = 15'h22xx then cliam and return locally
//         in soc,  ls addr = 15'h21xx then cliam and return locally
//         in soc,  ls addr = 15'h22xx for remote AA and send to remote side
// note: mailbox do not support remote read, only support local write and send a mailbox message to remote side. no need different address in soc and fpga
//        mailbox address = 15'h20xx in both soc and fpga
wire [31:0] sm_aa_internal_data = ss_aa_reg ? (r_ss_rw_addr[2] ? {31'b0, intr_status}
                                                                : {31'b0, intr_enable})
                                            : mb_regs[r_ss_rw_addr[4:2]];
// ----- LS - Data Source
// 1. SS RS data  - ss_rs_data 
// 2. ls_aa_internal data
assign s_rdata  = (ls_aa_reg | ls_aa_mbox) ?  ls_aa_internal_data  // for local_ls read
                                              : ss_rs_data;        // from SS read-response tuser=11

// ----------------------------
// mb_regs, intr_status, inter_enalbe
// LS write - s_wready qualify by ls_aa_reg, ls_aa_mbox
// SS write - ss_t2 @ clk  qualify by ss_aa_reg ls_aa_mbox

reg r_ss_t2;   // one cycle after ss_t2 to ensure ss address/data is valid
always @(posedge axis_clk or negedge axis_rst_n) begin
    if(! axis_rst_n)  begin
        r_ss_t2 <= 0;
    end else begin
        r_ss_t2 <= ss_t2;
    end
end

// 
// intr_status
//  set by ss write to mbox
//  reset by ls write to status with 1  (write one to clear)
// 
wire s_rvalid_out;

always @(posedge axis_clk or negedge axis_rst_n) begin
    if( !axis_rst_n ) begin
        intr_status <= 0;
    end else begin
        // intr_staus
        if(s_rvalid_out & (ls_aa_mbox_lr|ls_aa_mbox)) //local read aa_mbox_lr to clear (youwei change)
            intr_status <= 1'b0;
        else if(s_wready & ls_aa_reg_lw & s_awaddr[2] & s_wdata[0] & & s_wstrb[0]) //local write one to clear
            intr_status <= 1'b0;    // write-one-to clear 
        else if( r_ss_t2  & ss_aa_mbox_latch & (|r_ss_wstrb) ) //Remote write any mbox register to set
            intr_status <= 1'b1;    // mbox write set status
        else     
            intr_status <= intr_status;

    end
end 

always @(posedge axis_clk or negedge axis_rst_n) begin
    if( !axis_rst_n ) begin
        intr_enable <= 0;
    end else begin

        // intr_enable
        if(s_wready & ls_aa_reg_lw & !s_awaddr[2] & s_wstrb[0])    //local access 
            intr_enable <= s_wdata[0];
        else if( r_ss_t2  & ss_aa_reg_latch & !r_ss_rw_addr[2] & r_ss_wstrb[0])  //Remote access 
            intr_enable  <= r_ss_wdata[0];
        else 
            intr_enable <= intr_enable ;

        // mbox
        if(s_wready & ls_aa_mbox_lw) begin 
            if ( s_wstrb[0] ) mb_regs[s_awaddr[4:2]][7:0] <= s_wdata[7:0];
            else              mb_regs[s_awaddr[4:2]][7:0] <= mb_regs[s_awaddr[4:2]][7:0];
            if ( s_wstrb[1] ) mb_regs[s_awaddr[4:2]][15:8] <= s_wdata[15:8];
            else              mb_regs[s_awaddr[4:2]][15:8] <= mb_regs[s_awaddr[4:2]][15:8];
            if ( s_wstrb[2] ) mb_regs[s_awaddr[4:2]][23:16] <= s_wdata[23:16];
            else              mb_regs[s_awaddr[4:2]][23:16] <= mb_regs[s_awaddr[4:2]][23:16];
            if ( s_wstrb[3] ) mb_regs[s_awaddr[4:2]][31:24] <= s_wdata[31:24];
            else              mb_regs[s_awaddr[4:2]][31:24] <= mb_regs[s_awaddr[4:2]][31:24];
        end    
        else if( r_ss_t2  & ss_aa_mbox_latch ) begin

            if ( r_ss_wstrb[0] ) mb_regs[r_ss_rw_addr[4:2]][7:0] <= r_ss_wdata[7:0];
            else              mb_regs[r_ss_rw_addr[4:2]][7:0] <= mb_regs[r_ss_rw_addr[4:2]][7:0];
            if ( r_ss_wstrb[1] ) mb_regs[r_ss_rw_addr[4:2]][15:8] <= r_ss_wdata[15:8];
            else              mb_regs[r_ss_rw_addr[4:2]][15:8] <= mb_regs[r_ss_rw_addr[4:2]][15:8];
            if ( r_ss_wstrb[2] ) mb_regs[r_ss_rw_addr[4:2]][23:16] <= r_ss_wdata[23:16];
            else              mb_regs[r_ss_rw_addr[4:2]][23:16] <= mb_regs[r_ss_rw_addr[4:2]][23:16];
            if ( r_ss_wstrb[3] ) mb_regs[r_ss_rw_addr[4:2]][31:24] <= r_ss_wdata[31:24];
            else              mb_regs[r_ss_rw_addr[4:2]][31:24] <= mb_regs[r_ss_rw_addr[4:2]][31:24];
        end    
    end
end

// --- mb_irq ---
// asserts mb_irq when  intr_status = 1 & intr_enable
//
assign mb_irq = intr_status & intr_enable; 

// -------------------------------------------------------
// LS State Machine - Tracking LS -> SM Conversion
// Note： LS State machine & SS State machine can not run currently
//  LS read AA reg + MBOX LS_RD -> LS_R_DONE
//  LS write AA_reg       LS_WR -> LS_W_DONE
//  LS write AA_MBOX   pass to FPGA -> LS_WR_SM1
// -------------------------------------------------------
reg [6:0] ls_sm_fsm;

//
// sm fsm state encoding is used to generate related control signal
//                         {rd_ss_wait_rs, mbox, ls_cyc, ls_wr, ls_sm_tvalid_cyc, w1/w2 or ss_read, done}
`define LS_IDLE             7'b0_0_0_0_0_0_0              
`define LS_RD               7'b0_0_1_0_0_0_0
`define LS_WR               7'b0_0_1_1_0_0_0
`define LS_WR_SM1           7'b0_0_1_1_1_0_0
`define LS_WR_SM2           7'b0_0_1_1_1_1_0
`define LS_RD_SM_REQ        7'b0_0_1_0_1_1_0
`define LS_RD_SS_WAIT_RS    7'b1_0_1_0_0_0_0
`define LS_R_DONE           7'b0_0_1_0_0_0_1
`define LS_W_DONE           7'b0_0_1_1_0_0_1
`define LS_MBOXW            7'b0_1_1_1_0_0_1
`define LS_MBOXW_SM1        7'b0_1_1_1_1_0_0
`define LS_MBOXW_SM2        7'b0_1_1_1_1_1_0

wire sm_tvalid;

// cycle indicator and control signal generaion
wire   ls_mbox = ls_sm_fsm[5];
assign ls_cyc = ls_sm_fsm[4];
wire   ls_only_cyc = ls_sm_fsm[4] & !ls_sm_fsm[2];  // LS_RD, LS_WR 
assign ls_wr  = ls_sm_fsm[3];
wire   ls_sm_tvalid_cyc = ls_sm_fsm[2];
wire   sm_wr_t1 = (ls_sm_fsm == `LS_WR_SM1) || (ls_sm_fsm == `LS_MBOXW_SM1);
wire   sm_wr_t2 = (ls_sm_fsm == `LS_WR_SM2) || (ls_sm_fsm == `LS_MBOXW_SM2);
wire   sm_read_t = (ls_sm_fsm == `LS_RD_SM_REQ);
wire   ls_r_done = (ls_sm_fsm == `LS_R_DONE);
wire   ls_done  = ls_sm_fsm[0];
wire   ls_rd_ss_wait_rs = (ls_sm_fsm == `LS_RD_SS_WAIT_RS);


// interface signals  - axilite slave
assign s_awready = ls_cyc & ls_wr & ls_done;
assign s_wready  = s_awready;
assign s_arready  = (ls_sm_fsm == `LS_RD);
assign s_rvalid_out=ls_cyc & !ls_wr & ls_done;
assign s_rvalid = s_rvalid_out;

// interface signals  - axis master
assign aa_as_tvalid = sm_tvalid;                           //sm_tvalid = ss_sm_cyc | ls_sm_tvalid_cyc

// ---- SM - data has several sources
// 1. LS write - 1st T = r_ls_wstrb + r_ls_rw_addr
//               2nd T = r_ls_wdata
// 2. LS read = 4'b0000 + r_ls_rw_addr
// 3. SS read response  : r_lm_rs_data
// 
assign aa_as_tdata =  ({32{sm_wr_t1}}  & {r_ls_wstrb, r_ls_rw_addr[27:0]} )     // from local to remote write(include mbox write), local_ls write t1 -> local_sm write 
                   |  ({32{sm_wr_t2}}  & r_ls_wdata )                           // from local to remote write(include mbox write), local_ls write t2 -> local_sm write 
                   |  ({32{sm_read_t}}  & {4'b0000, r_ls_rw_addr[27:0]} )       // from local to remote read, local_ls read -> local_sm read
                   |  ({32{ss_sm_cyc & !ss_aa_reg_latch}} & r_lm_rs_data )          // remote_ls read -> remote_sm read -> local_ss read -> local_lm read_resp -> local_sm read_resp
                   |  ({32{ss_sm_cyc  &  ss_aa_reg_latch}} & sm_aa_internal_data)   // remote_ls read -> remote_sm read -> local_ss read -> local_lm read_resp -> local_sm read_resp
                   ;

assign aa_as_tstrb = (ls_wr? r_ls_wstrb : 4'b1111);     //from local to remote write use r_ls_wstrb, local_ls write -> local_sm write 
                                                          //from local to remote read use 4'b1111 ? local_ls read -> local_sm read
                                                          //from remote remote_ls read  -> remote_sm read -> local_ss read -> local_lm read_resp -> local_sm read_resp use 4'b1111
assign aa_as_tkeep = 0;
assign aa_as_tlast = 1'b1;
assign aa_as_tuser = ls_wr? TUSER_AXILITE_WRITE : 
                              (sm_read_t? TUSER_AXILITE_READ_REQ : TUSER_AXILITE_READ_CPL) ;


// control signals
// {ls_sm_enable, ls_sm_wr, sm_ready, sm_rs_ready}
// Note: LS, SS State machine is exclusive - when ss_cyc is ongoing then pending ls_sm_enable until ss_cyc done.
// SS state machine with higher priority then LS State machine when both in IDLE state and try to move to next state.
wire ls_sm_enable = !((ss_lm_fsm == `SS_IDLE) & ss_lm_enable) & !ss_cyc & cc_aa_enable & ((s_awvalid & s_wvalid) | s_arvalid);   // axilite AW & W AR request asserts
wire ls_sm_wr = s_awvalid;                  // axilite AW - write transaction
wire sm_ready = as_aa_tready;               // sm bus ready if write 2 cycle
wire ss_rs_ready = as_aa_tvalid & ss_rs_cyc; // axis slave receives read completion
wire ls_ready  = ls_sm_wr ? ls_done : ls_done & s_rready;      // ls read need to wait s_rready

// State Machine - ls_sm_fsm
always @(posedge axis_clk or negedge axis_rst_n) begin   // asynchronous reset
    if( !axis_rst_n ) begin
        ls_sm_fsm <= `LS_IDLE;
    end else begin
        case(ls_sm_fsm) 
            `LS_IDLE : 
                if(ls_sm_enable) begin
                    if(ls_sm_wr) ls_sm_fsm <= `LS_WR;
                    else         ls_sm_fsm <= `LS_RD;
                end else begin
                                ls_sm_fsm <= `LS_IDLE;
                end
            `LS_WR:  
                if(ls_aa_reg_lw)          ls_sm_fsm <= `LS_W_DONE;    
                else if(ls_aa_mbox_lw)    ls_sm_fsm <= `LS_MBOXW;    
                else                      ls_sm_fsm <= `LS_WR_SM1;
            `LS_WR_SM1: 
                if(sm_ready)    ls_sm_fsm <= `LS_WR_SM2;
                else            ls_sm_fsm <= `LS_WR_SM1;
            `LS_WR_SM2:
                if(sm_ready)    ls_sm_fsm <= `LS_W_DONE;
                else            ls_sm_fsm <= `LS_WR_SM2;
            `LS_RD:             
                if( ls_aa_reg_lr || ls_aa_mbox_lr ) ls_sm_fsm <= `LS_R_DONE; 
                else                               ls_sm_fsm <= `LS_RD_SM_REQ;
            `LS_RD_SM_REQ:                  // send 1T read request
                if(sm_ready)    ls_sm_fsm <= `LS_RD_SS_WAIT_RS;
                else            ls_sm_fsm <= `LS_RD_SM_REQ;
            `LS_RD_SS_WAIT_RS:
                if(ss_rs_ready) ls_sm_fsm <= `LS_R_DONE;
                else            ls_sm_fsm <= `LS_RD_SS_WAIT_RS;
            `LS_R_DONE:           
                if(ls_ready)    ls_sm_fsm <= `LS_IDLE;
                else            ls_sm_fsm <= `LS_R_DONE;
            `LS_W_DONE:           
                if(ls_ready)    ls_sm_fsm <= `LS_IDLE;
                else            ls_sm_fsm <= `LS_W_DONE;
            `LS_MBOXW:           
                if(ls_ready)    ls_sm_fsm <= `LS_MBOXW_SM1;
                else            ls_sm_fsm <= `LS_MBOXW;
            `LS_MBOXW_SM1: 
                if(sm_ready)    ls_sm_fsm <= `LS_MBOXW_SM2;
                else            ls_sm_fsm <= `LS_MBOXW_SM1;
            `LS_MBOXW_SM2:
                if(sm_ready)    ls_sm_fsm <= `LS_IDLE;
                else            ls_sm_fsm <= `LS_MBOXW_SM2;
            default:            ls_sm_fsm <= `LS_IDLE;
        endcase
    end
end 



// ------------------------------------------------------
// SS State machine - tracking SS -> LM 
//reg [6:0] ss_lm_fsm;

//
// sm fsm state encoding is used to generate related control signal
//  SS read AA inernal  SS_RD     -> SS_RD_SM_RS
//  SS write AA internal SS_WR_S2 -> SS_DONE
// 
/*
                          {ss_only_cyc, ss_wr, lm_cyc, ss_sm_cyc, w1/w2 or RD_LM_AR/R, done}
`define SS_IDLE             7'b0_0_0_0_0_0_0
`define SS_RD               7'b0_1_0_0_0_0_0
`define SS_WR_S1            7'b0_1_1_0_0_0_0
`define SS_WR_S2            7'b0_1_1_0_0_1_0
`define SS_WR_LM            7'b0_0_1_1_0_0_0
`define SS_WR_LM_AW         7'b1_0_1_1_0_0_0
`define SS_RD_LM_AR         7'b0_0_0_1_0_0_0
`define SS_RD_LM_R          7'b0_0_0_1_0_1_0
`define SS_RD_SM_RS         7'b0_0_0_0_1_0_0
`define SS_DONE             7'b0_0_0_0_0_0_1
*/

// cycle indicator and control signal generaion
assign ss_cyc = ss_lm_fsm[5] | ss_lm_fsm[3] | ss_lm_fsm[2];   //ss_only_cyc + lm_cyc + ss_sm_cyc
wire ss_only_cyc = ss_lm_fsm[5];
wire ss_wr  = ss_lm_fsm[4];
wire lm_cyc = ss_lm_fsm[3];
wire   lm_ar_cyc = ( ss_lm_fsm == `SS_RD_LM_AR);
assign ss_sm_cyc = ss_lm_fsm[2];
wire ss_t1  = ss_wr & !ss_lm_fsm[1];
assign ss_t2  = ss_wr & ss_lm_fsm[1];
wire ss_done  = ss_lm_fsm[0];

//wire ss_rd = ~ss_wr;

// combine from lm->sm
assign sm_tvalid = ss_sm_cyc | ls_sm_tvalid_cyc;    //from ss_sm_cyc is from remote, ls_sm_tvalid_cyc is from local

// interface signals - axis slave
// 1. remote_sm to local_ss read req
// 2. remote_sm to local_ss write req (include remote to local mbox write)
// 3. remote_sm read_resp -> local_ss read_resp
//    - local_ls read -> loca_sm read -> remote_ss read -> remote_lm read_resp -> remote_sm read_resp -> local_ss read_resp
assign aa_as_tready = ss_only_cyc | ls_r_done;

// interface signal - axis master
//   assign aa_as_tdata 


reg r_m_arvalid;
// set by lm_cyc & !ss_wr;
// clear by m_arready
always @(posedge axis_clk or negedge axis_rst_n) begin   
    if( !axis_rst_n ) r_m_arvalid <= 1'b0;
    else if (r_m_arvalid == 1'b0 &&  lm_ar_cyc && !ss_wr )  r_m_arvalid <= 1'b1;
    else if ( (r_m_arvalid == 1'b1) && (m_arready == 1'b1) ) r_m_arvalid <= 1'b0;
    else r_m_arvalid <= r_m_arvalid;
end

reg r_m_rready;
// set by lm_cyc & !ss_wr;
// clear by m_rvalid
always @(posedge axis_clk or negedge axis_rst_n) begin   
    if( !axis_rst_n ) r_m_rready <= 1'b0;
    else if (r_m_rready == 1'b0 &&  lm_ar_cyc && !ss_wr )  r_m_rready <= 1'b1;
    else if ( (r_m_rready == 1'b1) && (m_rvalid == 1'b1) ) r_m_rready <= 1'b0;
    else r_m_rready <= r_m_rready;
end

// LM interface signal - lm master
//support slave device in lm interface assert m_awready then assert m_wready or at the same clock.
assign m_awvalid = lm_cyc & ss_wr & (ss_lm_fsm == `SS_WR_LM);
assign m_wvalid  = lm_cyc & ss_wr & ( (ss_lm_fsm == `SS_WR_LM) | (ss_lm_fsm == `SS_WR_LM_AW) );
assign m_arvalid = r_m_arvalid; // m_arvalid de-assert when detect m_arready assert
assign m_rready  = r_m_rready;  // m_rready de-assert when detect m_rvalid assert


// control signals
// Note:  1. LS, SS state mchine are exclusive
//        2. limitation: dead lock issue, if remote side send a read request and ss_aa_reg=1. current design do not assert tready in SS then dead lock.
//        3. dead lock issue - both side issue mailbox write
//            workaround - SS state mahcine from IDLE to next state when ss_wr_cyc=1

// ss_lm_enable in below conditions
// 1. no on going ls cycle and current request from remote sm to local ss read cycle address not in aa_reg range.
//    - for remote sm to local ss read_resp cycle (ss_rs_cyc) do not let ss_lm_enable=1
// 2. remote sm to local ss is write cycle 
//
// limitation : dead lock when both side issue cfg read to remote side at the same time
// - for example 
//    A. soc  issue cfg read request to fpga then the soc  ls_cyc=1 and isseu read req from soc's  SM to fpga's ss.
//    in soc's view point, the ls_sys=1 and ss_rd_cyc=1 then keep ss_lm_enable = 0
//    B. fpga issue cfg read request to soc  then the fpga ls_cyc=1 and isseu read req from fpga's SM to soc's ss.
//    in fpga's view point, the ls_sys=1 and ss_rd_cyc=1 then keep ss_lm_enable = 0
//    - dead lock in both side, the ss_lm_enable keep = 0.
// - usage : in most case only fpga need issue remote cfg read for debugging.
// - improve solution: use mailbox as a communication chaneel for sw to grant/release the remote cfg access right. The spec is defeined by software if need.(TBD)

assign ss_lm_enable = (!ls_cyc & ss_rd_cyc & !ss_aa_reg & as_aa_tvalid ) || (ss_wr_cyc & as_aa_tvalid );

        
// State Machine - ss_lm_fsm
always @(posedge axis_clk or negedge axis_rst_n) begin   // asynchronous reset
    if( !axis_rst_n ) begin
        ss_lm_fsm <= `SS_IDLE;
    end else begin
        case(ss_lm_fsm) 
            `SS_IDLE: 
                if(ss_lm_enable) begin
                    if(ss_wr_cyc)             ss_lm_fsm <=  `SS_WR_S1;
                    else if(ss_rd_cyc)        ss_lm_fsm <= `SS_RD;
                    else                      ss_lm_fsm <= `SS_IDLE;
                end 
                else begin
                    ss_lm_fsm <= `SS_IDLE;
                end
            `SS_WR_S1:  
                if(as_aa_tvalid)   ss_lm_fsm <= `SS_WR_S2;
                else               ss_lm_fsm <= `SS_WR_S1;
            `SS_WR_S2:
                if(as_aa_tvalid)   begin
                    if(ss_aa_reg_latch | ss_aa_mbox_latch)  ss_lm_fsm <= `SS_DONE;
                    else                        ss_lm_fsm <= `SS_WR_LM;
                end 
                else  begin 
                    ss_lm_fsm <= `SS_WR_S2;
                end
            `SS_WR_LM:
                if(m_awready && m_wready)       ss_lm_fsm <= `SS_DONE;      
                else if(m_awready)              ss_lm_fsm <= `SS_WR_LM_AW;
                else                            ss_lm_fsm <= `SS_WR_LM;
            `SS_WR_LM_AW:
                if(m_wready)        ss_lm_fsm <= `SS_DONE;
                else                ss_lm_fsm <= `SS_WR_LM_AW;
            `SS_RD:
                if(ss_aa_reg | ss_aa_mbox) ss_lm_fsm <= `SS_RD_SM_RS;
                else                      ss_lm_fsm <= `SS_RD_LM_AR;    //read cfg target not in AA
            `SS_RD_LM_AR:
                if( !m_arready )                ss_lm_fsm <= `SS_RD_LM_AR;
                else if( m_arready & !m_rvalid ) ss_lm_fsm <= `SS_RD_LM_R;
                else                            ss_lm_fsm <= `SS_RD_SM_RS;
            `SS_RD_LM_R:
                if( !m_rvalid )      ss_lm_fsm <= `SS_RD_LM_R;
                else                 ss_lm_fsm <= `SS_RD_SM_RS;
            `SS_RD_SM_RS:
                if( !as_aa_tready)   ss_lm_fsm <= `SS_RD_SM_RS;
                else                 ss_lm_fsm <= `SS_DONE;
            `SS_DONE:               ss_lm_fsm <= `SS_IDLE;
            default:            ss_lm_fsm <= `SS_IDLE;
        endcase
    end
end        


// ------------------------------------------------------
//  Address / Data Storage
// ------------------------------------------------------

// ---------   SS    ---------------
// SS - r_ss_rw_addr, r_ss_wdata, r_ss_wstrb, r_tuser
//  - ss side address/data latch
// Note: it does not need reset, why ? when it is used, the content will be valid anyway
// -------------------------

always @( posedge axis_clk ) begin              // T1 - address
    if( ss_only_cyc && (!ss_wr | ss_t1) ) begin     //ss_only_cyc = aa_as_tready
                                                        //latch addr, strb and user when read or ss_t1
        r_ss_rw_addr <= as_aa_tdata[27:0] | 32'h3000_0000;  //for received cfg R/W request in ss, update address bit[31:28]= 4'h3 in local for send to lm connect to config control.
        r_ss_wstrb <= as_aa_tdata[31:28];                          //how to use as_aa_tstrb?
        r_tuser <= as_aa_tuser;
    end else begin
        r_ss_rw_addr <= r_ss_rw_addr;
        r_ss_wstrb <= r_ss_wstrb;
        // r_tuser <= as_aa_tuser;
        r_tuser <= r_tuser;
    end
end

//r_ss_wdata come from below source
// 1. SS write - r_ss_wdata come from as_aa_tdata
//    when remote_ls write -> remote_sm write t2 -> local_ss write t2
// 2. SS read_resp r_ss_wdata come from as_aa_tdata
//    when local_ls read -> local_sm read -> remote_ss read -> remote_lm read_resp -> remote_sm read_resp -> local_ss read_resp

always @(posedge axis_clk) begin                // T2 - data
    if( ( ss_only_cyc && ss_t2 ) || (as_aa_tvalid && ls_rd_ss_wait_rs ) )     //ss_only_cyc = aa_as_tready
                                                                                  //early capture data when as_aa_tvalid
          r_ss_wdata <= as_aa_tdata;                      //ss_rs_data = r_ss_wdata, it is share. 
    else  r_ss_wdata <= r_ss_wdata;
end


// ----------  LS     ---------------------------
// r_ls_rw_addr   - LS address    @awvaid, arvalid
// r_ls_wdata       - LS write data @wvalid
// r_ls_wstrb      - ls write strb @awvalid
// 

always @( posedge axis_clk ) begin
    if( ls_only_cyc & (s_awvalid | s_arvalid))  begin   //use valid to latch addr.
        r_ls_rw_addr <= s_awvalid ? s_awaddr : s_araddr;   //r_ls_rw_addr[31:15] awlays = 0
    end else begin
        r_ls_rw_addr <= r_ls_rw_addr; 
    end
end

always @( posedge axis_clk ) begin
    if( ls_only_cyc & s_wvalid )  begin
        r_ls_wstrb <= s_wstrb;
        r_ls_wdata <= s_wdata;
    end else begin
        r_ls_wstrb <= r_ls_wstrb;
        r_ls_wdata <= r_ls_wdata;
    end
end


// ---------- LM   --------------------
//  r_lm_rs_data           // latch read response data in LM used for SM to return RS data
//
always @( posedge axis_clk ) begin
    if( m_rvalid && m_rready ) begin   
        r_lm_rs_data <= m_rdata;
    end else begin
        r_lm_rs_data <= r_lm_rs_data;
    end
end
 

endmodule // AXIL_AXIS







//////////////////////////////////////////////////////////////////////////////////
// Author : Tony Ho
//
// Create Date: 11/20/2023
// Design Name:
// Module Name: AXIL_SLAV
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module AXIL_SLAV #( parameter pADDR_WIDTH   = 12,
                    parameter pDATA_WIDTH   = 32
                  )
(
  input  wire                        awready_0,
  input  wire                        arready_0,
  input  wire                        wready_0,
  input  wire                        rvalid_0,
  input  wire  [(pDATA_WIDTH-1) : 0] rdata_0,
  input  wire                        awready_1,
  input  wire                        arready_1,
  input  wire                        wready_1,
  input  wire                        rvalid_1,
  input  wire  [(pDATA_WIDTH-1) : 0] rdata_1,
  input  wire                        awready_2,
  input  wire                        arready_2,
  input  wire                        wready_2,
  input  wire                        rvalid_2,
  input  wire  [(pDATA_WIDTH-1) : 0] rdata_2,
  input  wire                        awready_3,
  input  wire                        arready_3,
  input  wire                        wready_3,
  input  wire                        rvalid_3,
  input  wire  [(pDATA_WIDTH-1) : 0] rdata_3,
  output wire                        awvalid_0,
  output wire                [11: 0] awaddr,
  output wire                        arvalid_0,
  output wire                [11: 0] araddr,
  output wire                        wvalid_0,
  output wire                 [3: 0] wstrb_0,
  output wire  [(pDATA_WIDTH-1) : 0] wdata,
  output wire                        rready,
  output wire                        awvalid_1,
  output wire                        arvalid_1,
  output wire                        wvalid_1,
  output wire                 [3: 0] wstrb_1,
  output wire                        awvalid_2,
  output wire                        arvalid_2,
  output wire                        wvalid_2,
  output wire                 [3: 0] wstrb_2,
  output wire                        awvalid_3,
  output wire                        arvalid_3,
  output wire                        wvalid_3,
  output wire                 [3: 0] wstrb_3,
  input  wire                        axi_awvalid,
  input  wire                [14: 0] axi_awaddr,
  input  wire                        axi_arvalid,
  input  wire                [14: 0] axi_araddr,
  input  wire                        axi_wvalid,
  input  wire                 [3: 0] axi_wstrb,
  input  wire  [(pDATA_WIDTH-1) : 0] axi_wdata,
  input  wire                        axi_rready,
  input  wire                        cc_up_enable,
  output wire                        axi_awready,
  output wire                        axi_arready,
  output wire                        axi_wready,
  output wire                        axi_rvalid,
  output wire  [(pDATA_WIDTH-1) : 0] axi_rdata,
  input  wire                        axi_clk,
  input  wire                        axi_reset_n,
  input  wire                 [4: 0] user_prj_sel
);

wire  [3:0] axi_awready_bus;
assign axi_awready = |axi_awready_bus;

wire  [3:0] axi_wready_bus;
assign axi_wready = |axi_wready_bus;

wire  [3:0] axi_arready_bus;
assign axi_arready = |axi_arready_bus;

wire  [3:0] axi_rvalid_bus;
assign axi_rvalid = |axi_rvalid_bus;

wire  [(pDATA_WIDTH-1) : 0] axi_rdata_bus[3:0];
assign axi_rdata = axi_rdata_bus[0] | axi_rdata_bus[1] | axi_rdata_bus[2] | axi_rdata_bus[3];

//user project 0 
assign awvalid_0 = ( (user_prj_sel == 5'b00000) && cc_up_enable) ? axi_awvalid : 0;
assign axi_awready_bus[0] = ( (user_prj_sel == 5'b00000) && cc_up_enable) ? awready_0 : 0;
assign awaddr = axi_awaddr[11:0];
assign wstrb_0 = axi_wstrb;    //[TODO] share wstrb for all user projects.

assign wvalid_0 = ( (user_prj_sel == 5'b00000) && cc_up_enable) ? axi_wvalid : 0;
assign axi_wready_bus[0] = ( (user_prj_sel == 5'b00000) && cc_up_enable) ? wready_0 : 0;
assign wdata = axi_wdata;

assign arvalid_0 = ( (user_prj_sel == 5'b00000) && cc_up_enable) ? axi_arvalid : 0;
assign axi_arready_bus[0] = ( (user_prj_sel == 5'b00000) && cc_up_enable) ? arready_0 : 0;
assign araddr = axi_araddr;

assign axi_rvalid_bus[0] = ( (user_prj_sel == 5'b00000) && cc_up_enable) ? rvalid_0 : 0;
assign rready = axi_rready;
assign axi_rdata_bus[0] = ( (user_prj_sel == 5'b00000) && cc_up_enable) ? rdata_0 : 0;

//user project 1 
assign awvalid_1 = ( (user_prj_sel == 5'b00001) && cc_up_enable) ? axi_awvalid : 0;
assign axi_awready_bus[1] = ( (user_prj_sel == 5'b00001) && cc_up_enable) ? awready_1 : 0;
assign awaddr = axi_awaddr[11:0];
assign wstrb_1 = axi_wstrb;    //[TODO] share wstrb for all user projects.

assign wvalid_1 = ( (user_prj_sel == 5'b00001) && cc_up_enable) ? axi_wvalid : 0;
assign axi_wready_bus[1] = ( (user_prj_sel == 5'b00001) && cc_up_enable) ? wready_1 : 0;
assign wdata = axi_wdata;

assign arvalid_1 = ( (user_prj_sel == 5'b00001) && cc_up_enable) ? axi_arvalid : 0;
assign axi_arready_bus[1] = ( (user_prj_sel == 5'b00001) && cc_up_enable) ? arready_1 : 0;
assign araddr = axi_araddr;

assign axi_rvalid_bus[1] = ( (user_prj_sel == 5'b00001) && cc_up_enable) ? rvalid_1 : 0;
assign rready = axi_rready;
assign axi_rdata_bus[1] = ( (user_prj_sel == 5'b00001) && cc_up_enable) ? rdata_1 : 0;

//user project 2 
assign awvalid_2 = ( (user_prj_sel == 5'b00010) && cc_up_enable) ? axi_awvalid : 0;
assign axi_awready_bus[2] = ( (user_prj_sel == 5'b00010) && cc_up_enable) ? awready_2 : 0;
assign awaddr = axi_awaddr[11:0];
assign wstrb_2 = axi_wstrb;    //[TODO] share wstrb for all user projects.

assign wvalid_2 = ( (user_prj_sel == 5'b00010) && cc_up_enable) ? axi_wvalid : 0;
assign axi_wready_bus[2] = ( (user_prj_sel == 5'b00010) && cc_up_enable) ? wready_2 : 0;
assign wdata = axi_wdata;

assign arvalid_2 = ( (user_prj_sel == 5'b00010) && cc_up_enable) ? axi_arvalid : 0;
assign axi_arready_bus[2] = ( (user_prj_sel == 5'b00010) && cc_up_enable) ? arready_2 : 0;
assign araddr = axi_araddr;

assign axi_rvalid_bus[2] = ( (user_prj_sel == 5'b00010) && cc_up_enable) ? rvalid_2 : 0;
assign rready = axi_rready;
assign axi_rdata_bus[2] = ( (user_prj_sel == 5'b00010) && cc_up_enable) ? rdata_2 : 0;

//user project 3 
assign awvalid_3 = ( (user_prj_sel == 5'b00011) && cc_up_enable) ? axi_awvalid : 0;
assign axi_awready_bus[3] = ( (user_prj_sel == 5'b00011) && cc_up_enable) ? awready_3 : 0;
assign awaddr = axi_awaddr[11:0];
assign wstrb_3 = axi_wstrb;    //[TODO] share wstrb for all user projects.

assign wvalid_3 = ( (user_prj_sel == 5'b00011) && cc_up_enable) ? axi_wvalid : 0;
assign axi_wready_bus[3] = ( (user_prj_sel == 5'b00011) && cc_up_enable) ? wready_3 : 0;
assign wdata = axi_wdata;

assign arvalid_3 = ( (user_prj_sel == 5'b00011) && cc_up_enable) ? axi_arvalid : 0;
assign axi_arready_bus[3] = ( (user_prj_sel == 5'b00011) && cc_up_enable) ? arready_3 : 0;
assign araddr = axi_araddr;

assign axi_rvalid_bus[3] = ( (user_prj_sel == 5'b00011) && cc_up_enable) ? rvalid_3 : 0;
assign rready = axi_rready;
assign axi_rdata_bus[3] = ( (user_prj_sel == 5'b00011) && cc_up_enable) ? rdata_3 : 0;


endmodule // AXIL_SLAV

//////////////////////////////////////////////////////////////////////////////////
// Author : Tony Ho
//
// Create Date: 11/20/2023
// Design Name:
// Module Name: AXIS_MSTR
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module AXIS_MSTR #( parameter pUSER_PROJECT_SIDEBAND_WIDTH = 5,
          parameter pADDR_WIDTH   = 12,
                    parameter pDATA_WIDTH   = 32
                  )
(
  output wire                        sm_tready,
  input  wire                        sm_tvalid_0,
  input  wire  [(pDATA_WIDTH-1) : 0] sm_tdata_0,
  input  wire                 [2: 0] sm_tid_0,

  input  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] sm_tupsb_0,

  input  wire                 [3: 0] sm_tstrb_0,
  input  wire                 [3: 0] sm_tkeep_0,
  input  wire                        sm_tlast_0,
  input  wire                        sm_tvalid_1,
  input  wire  [(pDATA_WIDTH-1) : 0] sm_tdata_1,
  input  wire                 [2: 0] sm_tid_1,

  input  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] sm_tupsb_1,

  input  wire                 [3: 0] sm_tstrb_1,
  input  wire                 [3: 0] sm_tkeep_1,
  input  wire                        sm_tlast_1,
  input  wire                        sm_tvalid_2,
  input  wire  [(pDATA_WIDTH-1) : 0] sm_tdata_2,
  input  wire                 [2: 0] sm_tid_2,

  input  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] sm_tupsb_2,

  input  wire                 [3: 0] sm_tstrb_2,
  input  wire                 [3: 0] sm_tkeep_2,
  input  wire                        sm_tlast_2,
  input  wire                        sm_tvalid_3,
  input  wire  [(pDATA_WIDTH-1) : 0] sm_tdata_3,
  input  wire                 [2: 0] sm_tid_3,

  input  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] sm_tupsb_3,

  input  wire                 [3: 0] sm_tstrb_3,
  input  wire                 [3: 0] sm_tkeep_3,
  input  wire                        sm_tlast_3,
  input  wire                        m_tready,
  output wire                        m_tvalid,
  output wire  [(pDATA_WIDTH-1) : 0] m_tdata,
  output wire                 [1: 0] m_tuser,

   output  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] m_tupsb,

  output wire                 [3: 0] m_tstrb,
  output wire                 [3: 0] m_tkeep,
  output wire                        m_tlast,
  input  wire                        axis_clk,
  input  wire                        axi_reset_n,
  input  wire                        axis_rst_n,
  input  wire                 [4: 0] user_prj_sel
);

//common part
assign sm_tready =  m_tready;

//bus
wire [3:0] sm_tvalid_bus;
assign  m_tvalid = |sm_tvalid_bus;

wire [(pDATA_WIDTH-1) : 0] sm_tdata_bus[3:0];
assign  m_tdata = sm_tdata_bus[0] | sm_tdata_bus[1] | sm_tdata_bus[2] | sm_tdata_bus[3];

//wire [2: 0] sm_tid_bus;


  wire [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] sm_tupsb_bus[3:0];
  assign  m_tupsb = sm_tupsb_bus[0] | sm_tupsb_bus[1] | sm_tupsb_bus[2] | sm_tupsb_bus[3];


wire [3: 0] sm_tstrb_bus[3:0];
assign  m_tstrb = sm_tstrb_bus[0] | sm_tstrb_bus[1] | sm_tstrb_bus[2] | sm_tstrb_bus[3];

wire [3: 0] sm_tkeep_bus[3:0];
assign  m_tkeep = sm_tkeep_bus[0] | sm_tkeep_bus[1] | sm_tkeep_bus[2] | sm_tkeep_bus[3];

wire [3: 0] sm_tlast_bus[3:0];
assign  m_tlast = sm_tlast_bus[0] | sm_tlast_bus[1] | sm_tlast_bus[2] | sm_tlast_bus[3];

//user project 0 
assign sm_tvalid_bus[0] =  (user_prj_sel == 5'b00000)  ? sm_tvalid_0 : 0;
assign sm_tdata_bus[0] = (user_prj_sel == 5'b00000)  ? sm_tdata_0 : 0;

  assign sm_tupsb_bus[0] = (user_prj_sel == 5'b00000)  ? sm_tupsb_0 : 0;

assign sm_tstrb_bus[0] = (user_prj_sel == 5'b00000)  ? sm_tstrb_0 : 0;
assign sm_tkeep_bus[0] = (user_prj_sel == 5'b00000)  ? sm_tkeep_0 : 0;
assign sm_tlast_bus[0] = (user_prj_sel == 5'b00000)  ? sm_tlast_0 : 0;

//user project 1 
assign sm_tvalid_bus[1] =  (user_prj_sel == 5'b00001)  ? sm_tvalid_1 : 0;
assign sm_tdata_bus[1] = (user_prj_sel == 5'b00001)  ? sm_tdata_1 : 0;

  assign sm_tupsb_bus[1] = (user_prj_sel == 5'b00001)  ? sm_tupsb_1 : 0;

assign sm_tstrb_bus[1] = (user_prj_sel == 5'b00001)  ? sm_tstrb_1 : 0;
assign sm_tkeep_bus[1] = (user_prj_sel == 5'b00001)  ? sm_tkeep_1 : 0;
assign sm_tlast_bus[1] = (user_prj_sel == 5'b00001)  ? sm_tlast_1 : 0;

//user project 2 
assign sm_tvalid_bus[2] =  (user_prj_sel == 5'b00010)  ? sm_tvalid_2 : 0;
assign sm_tdata_bus[2] = (user_prj_sel == 5'b00010)  ? sm_tdata_2 : 0;

  assign sm_tupsb_bus[2] = (user_prj_sel == 5'b00010)  ? sm_tupsb_2 : 0;

assign sm_tstrb_bus[2] = (user_prj_sel == 5'b00010)  ? sm_tstrb_2 : 0;
assign sm_tkeep_bus[2] = (user_prj_sel == 5'b00010)  ? sm_tkeep_2 : 0;
assign sm_tlast_bus[2] = (user_prj_sel == 5'b00010)  ? sm_tlast_2 : 0;

//user project 3 
assign sm_tvalid_bus[3] =  (user_prj_sel == 5'b00011)  ? sm_tvalid_3 : 0;
assign sm_tdata_bus[3] = (user_prj_sel == 5'b00011)  ? sm_tdata_3 : 0;

  assign sm_tupsb_bus[3] = (user_prj_sel == 5'b00011)  ? sm_tupsb_3 : 0;

assign sm_tstrb_bus[3] = (user_prj_sel == 5'b00011)  ? sm_tstrb_3 : 0;
assign sm_tkeep_bus[3] = (user_prj_sel == 5'b00011)  ? sm_tkeep_3 : 0;
assign sm_tlast_bus[3] = (user_prj_sel == 5'b00011)  ? sm_tlast_3 : 0;

assign m_tuser       = 2'b00;    //MUST be 2'b00 for user project output axis from UP to AS.


endmodule // AXIS_MSTR

//////////////////////////////////////////////////////////////////////////////////
// Author : Tony Ho
//
// Create Date: 11/20/2023
// Design Name:
// Module Name: AXIS_SLAV
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module AXIS_SLAV #( parameter pUSER_PROJECT_SIDEBAND_WIDTH = 5,
          parameter pADDR_WIDTH   = 12,
                    parameter pDATA_WIDTH   = 32
                  )
(
  output wire                        ss_tvalid_0,
  output wire  [(pDATA_WIDTH-1) : 0] ss_tdata,
  output wire                 [1: 0] ss_tuser,

  output  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] ss_tupsb,

  output wire                 [3: 0] ss_tstrb,
  output wire                 [3: 0] ss_tkeep,
  output wire                        ss_tlast,
  output wire                        ss_tvalid_1,
  output wire                        ss_tvalid_2,
  output wire                        ss_tvalid_3,
  input  wire                        ss_tready_0,
  input  wire                        ss_tready_1,
  input  wire                        ss_tready_2,
  input  wire                        ss_tready_3,
  input  wire                        s_tvalid,
  input  wire  [(pDATA_WIDTH-1) : 0] s_tdata,
  input  wire                 [1: 0] s_tuser,

  input  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] s_tupsb,

  input  wire                 [3: 0] s_tstrb,
  input  wire                 [3: 0] s_tkeep,
  input  wire                        s_tlast,
  output wire                        s_tready,
  input  wire                        axis_clk,
  input  wire                        axi_reset_n,
  input  wire                        axis_rst_n,
  input  wire                 [4: 0] user_prj_sel
);

//common part
assign ss_tdata =  s_tdata;
assign ss_tuser =  2'b00;    //UP always received tuser = 2'b00, the tuser is used by AS, should not send to UP.

  assign ss_tupsb =  s_tupsb;

assign ss_tstrb =  s_tstrb;
assign ss_tkeep =  s_tkeep;
assign ss_tlast =  s_tlast;

wire [3:0] s_tready_bus;
assign  s_tready = |s_tready_bus;

//user project 0 
assign ss_tvalid_0 =  (user_prj_sel == 5'b00000)  ? s_tvalid : 0;
assign s_tready_bus[0] = (user_prj_sel == 5'b00000)  ? ss_tready_0 : 0;

//user project 1 
assign ss_tvalid_1 =  (user_prj_sel == 5'b00001)  ? s_tvalid : 0;
assign s_tready_bus[1] = (user_prj_sel == 5'b00001)  ? ss_tready_1 : 0;

//user project 2 
assign ss_tvalid_2 =  (user_prj_sel == 5'b00010)  ? s_tvalid : 0;
assign s_tready_bus[2] = (user_prj_sel == 5'b00010)  ? ss_tready_2 : 0;

//user project 3 
assign ss_tvalid_3 =  (user_prj_sel == 5'b00011)  ? s_tvalid : 0;
assign s_tready_bus[3] = (user_prj_sel == 5'b00011)  ? ss_tready_3 : 0;




endmodule // AXIS_SLAV

//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: nthuyouwei
// 
// Create Date: 09/06/2024 10:00:00 AM
// Design Name: 
// Module Name: fifo
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////




/*****************  how to use this fifo
This is a FIFO designed using a single port sram. Due to the nature of the single port sram, we cannot read and write simultaneously. 
To solve this prob, I used double data width to solve the problem by reading two data entries at once, aiming to maintain the latency the same as a normal FIFO under ideal conditions (i.e., 1T delay for reading). 
In the worst case, if write/read commands arrive simultaneously, we will first check if writing is possible before reading, which could cause a maximum delay of 3T for reads.

Additionally, this design has two modes:

- mode = 1: The read protocol uses the AXI-stream protocol, and the write protocol operates such that when `w_rdy` is 1, it indicates that the FIFO has at least the threshold space available for writing. 
When the other end receives `w_rdy` as 1, it can send `w_vld`, as the FIFO will write directly upon receiving `w_vld`.

- mode = 0: Both read and write protocols use the AXI-stream protocol. Note: `w_rdy` = !full.
***********************/


/********************setting
WIDTH is datawidth.
depth is fifo depth.
sram_datawidth is usually double of WIDTH(sram_datawidth>=2*WIDTH).
mode is 1/0
*******************/


module fifo
#( parameter WIDTH = 45,
   parameter depth= 64,
   parameter sram_datawidth= 128,
   parameter mode=1 // mode 1 is for as, 0 is for la
)
(
    input axis_clk ,
    input axi_reset_n ,
    // write protocol
    input   w_vld,
    output  w_rdy,
    input [WIDTH-1:0] data_in,
    // read protocol
    input r_rdy,
    output  r_vld,
    output [WIDTH-1:0] data_out,
    // use for above_TH 
    input [7:0] TH_reg,
    // external sram io
    output sram_we,
    output[$clog2(depth)-1:0] sram_addr,
    output[sram_datawidth-1:0]sram_din,
    input [sram_datawidth-1:0] sram_dout
    );   
    localparam IDLE = 2'd0, WAIT_SRAM_READ = 2'd1, WAIT_FIFO_READ = 2'd2, NORMAL = 2'd3; // state machine part
    localparam sram_addr_width=$clog2(depth);
    localparam ptr_width=sram_addr_width+2; // LSB note even/odd times, MSB to decide full or not 
    reg [1:0] state;
    reg [1:0] state_next;
    reg [ptr_width-1:0] w_ptr;
    reg [ptr_width-1:0] r_ptr;
    wire [ptr_width-1:0] w_ptr_next;
    wire [ptr_width-1:0] r_ptr_next;
    assign w_ptr_next=w_ptr+1'b1;
    assign r_ptr_next=r_ptr+1'b1;
    wire empty;
    ///////////////////  above TH part//////////////////

                                         
    wire above_TH;
    assign above_TH=({w_ptr[ptr_width-1]==~r_ptr[ptr_width-1],w_ptr[ptr_width-2:0]}-{1'b0,r_ptr[ptr_width-2:0]})>TH_reg;
    
    ///////////////////  state machine////////// 
    //If it may directly reads from data_l, we need to ensure that it doesn't skip some data when it needs to read from SRAM.
    //After reads from data_l, Since the normal condition should starts with r_ptr[0] == 0, we need to add this state machine to make it corretly exec in normal condition. 
    // w_ptr==r_ptr_next ie reads from data_l.
    always @(posedge axis_clk or negedge axi_reset_n) begin
        if (!axi_reset_n)begin 
            state<=2'd0;
        end
        else begin
            state<=state_next;
        end
    end 

    always @(*) begin
        case(state)
            IDLE: begin   
                if(!(w_ptr==r_ptr_next|empty))begin
                    if(r_ptr[0]) state_next=WAIT_SRAM_READ;
                    else state_next=NORMAL;
                end
                else state_next=state;
            end
            WAIT_SRAM_READ: begin
                if(~sram_we) state_next=WAIT_FIFO_READ;
                else state_next=state;
            end
            WAIT_FIFO_READ:begin
                if(r_rdy) state_next=NORMAL;
                else state_next=state;
            end
            NORMAL:begin
                if(w_ptr==r_ptr_next) state_next=IDLE;
                else state_next=state;
            end
        endcase
    end 

    /////////////////////////// ptr part ///////////////////////////////////////////////////////////////////////////

    wire w_rdy_mode;
    assign w_rdy_mode=mode|w_rdy;
    always @(posedge axis_clk or negedge axi_reset_n) begin
        if (!axi_reset_n)begin 
            w_ptr<=0;
        end
        else begin
            if(w_vld & w_rdy_mode )w_ptr<=w_ptr_next;
            else  w_ptr<=w_ptr;
        end
    end 
    always @(posedge axis_clk or negedge axi_reset_n) begin
        if (!axi_reset_n)begin 
            r_ptr<=0;
        end
        else begin
            if(r_rdy & r_vld)r_ptr<=r_ptr_next;
            else  r_ptr<=r_ptr;
        end
    end 

///////////////////////////////// Write part ////////////////////////////////////////////////////////////////
//the MSB is different while the other bits are the same, it indicates that w_ptr has already completed one full cycle ahead of r_ptr, meaning it is full.  
// above th can remove if you not use 
    assign w_rdy= (mode==1)? ~above_TH : ~((w_ptr[ptr_width-1]==~r_ptr[ptr_width-1])&(w_ptr[ptr_width-2:0]==r_ptr[ptr_width-2:0]));  // not use full and empty 
    reg [WIDTH-1:0]data_in_l;

    always @(posedge axis_clk or negedge axi_reset_n) begin
        if (!axi_reset_n)begin 
            data_in_l<=0;
        end
        else begin
            if(w_vld & w_rdy_mode)
            data_in_l<=data_in;
            else 
            data_in_l<=data_in_l;
        end
    end 
///////////////////////////////////////////////////////////////////////////////////////////////////////////////

    reg sram_read_flag;
    wire sram_read_flag_next;
    assign sram_read_flag_next=((state==WAIT_SRAM_READ)&(~sram_we))|((state==NORMAL) & ~(~r_ptr[0] & r_vld &r_rdy) & (~sram_we & !(r_ptr_next[ptr_width-2:1]==w_ptr[ptr_width-2:1])));
    always @(posedge axis_clk or negedge axi_reset_n) begin
        if (!axi_reset_n)
            sram_read_flag<=0;
        else 
            sram_read_flag<=sram_read_flag_next;
    end 


    assign sram_we= w_vld & w_ptr[0]; // only write in sram in w_ptr[0]==1 mean even times.
    // when we is w_ptr and ,re is r_ptr_next or r_ptr decided by state machine case.  
    assign sram_addr=(sram_we)?w_ptr[ptr_width-2:1]:(state==NORMAL)?r_ptr_next[ptr_width-2:1]:r_ptr[ptr_width-2:1];
    assign sram_din ={{{sram_datawidth-2*WIDTH}{1'b0}},data_in,data_in_l};//from latch and input data
    
    
    
    
    /////////////////// Read part ///////////////////////////
    wire [WIDTH-1:0] sram_out_even;
    wire [WIDTH-1:0] sram_out_odd;
    assign sram_out_even = sram_dout[WIDTH-1:0];
    assign sram_out_odd = sram_dout[2*WIDTH-1:WIDTH];



    reg [WIDTH-1:0] data_out_odd;
    reg [WIDTH-1:0] data_out_even;
       
    always @(posedge axis_clk or negedge axi_reset_n) begin
        if (!axi_reset_n)begin 
            data_out_odd<=0;
        end
        else begin
            if(sram_read_flag)
            data_out_odd<=sram_out_odd;
            else 
            data_out_odd<=data_out_odd;
        end
    end 
    always @(posedge axis_clk or negedge axi_reset_n) begin
        if (!axi_reset_n)begin 
            data_out_even<=0;
        end
        else begin
            if(sram_read_flag)
            data_out_even<=sram_out_even;
            else 
            data_out_even<=data_out_even;
        end
    end 
    reg [WIDTH-1:0] data_out_odd_l;
    always @(posedge axis_clk or negedge axi_reset_n) begin
        if (!axi_reset_n)begin 
            data_out_odd_l<=0;
        end
        else begin
            if(~r_ptr[0])begin
                if(sram_read_flag)
                data_out_odd_l<=sram_out_odd;
                else 
                data_out_odd_l<=data_out_odd;
            end
            else 
            data_out_odd_l<=data_out_odd_l;
        end
    end 

    reg r_vld_even;
    assign empty=(w_ptr==r_ptr);


    // there are three conidtion :1. when r_ptr_next=w_ptr is always 1 becuase data is from data_l. and 2. state if is normal can divide into two condition read even or odd times to decide.and contion isn't normal only when state==WAIT fifo read can be 1.
    assign r_vld=((r_ptr_next==w_ptr)?1'b1:(state==NORMAL)?((r_ptr[0])?1'b1:r_vld_even):state==WAIT_FIFO_READ)& !empty;
    assign data_out=(r_ptr_next==w_ptr)?data_in_l: (state==NORMAL)?((r_ptr[0])?data_out_odd_l:(sram_read_flag)?sram_out_even:data_out_even):(sram_read_flag)?sram_out_odd:data_out_odd;  

  

    always@(posedge axis_clk or negedge axi_reset_n) begin
        if (!axi_reset_n) begin 
            r_vld_even <= 1'b0;
        end
        else begin
            if(state==NORMAL)begin
                if(~r_ptr[0] & r_vld &r_rdy)
                    r_vld_even <= 1'b0;
                else if (~sram_we & !(r_ptr_next[ptr_width-2:1]==w_ptr[ptr_width-2:1]))  //r_ptr_next[ptr_width-2:1]==w_ptr[ptr_width-2:1] to avoid reading before writing.
                    r_vld_even <= 1'b1;
                else 
                    r_vld_even<=r_vld_even;
                end
            else r_vld_even<=1'b0;
        end
    end

endmodule



// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype wire
/*
 *-------------------------------------------------------------
 *
 * user_project_wrapper
 *
 * This wrapper enumerates all of the pins available to the
 * user for the user project.
 *
 * An example user project is provided in this wrapper.  The
 * example should be removed and replaced with the actual
 * user project.
 *
 *-------------------------------------------------------------
 */

module user_project_wrapper #(parameter BITS = 32)
(
    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // Analog (direct connection to GPIO pad---use with caution)
    // Note that analog I/O is not available on the 7 lowest-numbered
    // GPIO pads, and so the analog_io indexing is offset from the
    // GPIO indexing by 7 (also upper 2 GPIOs do not have analog_io).

    // Independent clock (on independent integer divider)
    input   user_clock2,

    // User maskable interrupt signals
    output [2:0] user_irq
);

/*
assign wbs_ack_o   = 1'b0;
assign wbs_dat_o   = 32'd0;
assign la_data_out = 128'd0;
assign io_out      = 38'd0;
assign io_oeb      = 38'd0;
assign user_irq    = 3'd0;
*/
FSIC #(.BITS( BITS )) u_fsic  (

                      // MGMT SoC Wishbone Slave
                      .wb_rst      (wb_rst_i),                // I
                      .wb_clk      (wb_clk_i),                // I

                      .wbs_adr     (wbs_adr_i),               // I  32
                      .wbs_wdata   (wbs_dat_i),               // I  32
                      .wbs_sel     (wbs_sel_i),               // I  4
                      .wbs_cyc     (wbs_cyc_i),               // I
                      .wbs_stb     (wbs_stb_i),               // I
                      .wbs_we      (wbs_we_i),                // I

                      .wbs_ack     (wbs_ack_o),               // O
                      .wbs_rdata   (wbs_dat_o),               // O  32

                      // Logic Analyzer
		      // Removed. fsic has no below la interfaces.
                      //.la_data_in  (la_data_in),              // I  128
                      //.la_oenb     (la_oenb),                 // I  128
                      //.la_data_out (la_data_out),             // O  128

                      // IO Pads
                      .io_in       (io_in),                   // I  38
                      .io_out      (io_out),                  // O  38
                      .io_oeb      (io_oeb),                  // O  38

                      // IRQ
                      .user_irq    (user_irq),                // O  3

                      // MISC (Independent clock, on independent integer divider)
                      .user_clock2 (user_clock2)              // I
                     );


endmodule	// user_project_wrapper

`default_nettype wire
//////////////////////////////////////////////////////////////////////////////////
// Author : Tony Ho
//
// Create Date: 11/20/2023
// Design Name:
// Module Name: USER_SUBSYS
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module USER_SUBSYS #( parameter pUSER_PROJECT_SIDEBAND_WIDTH = 5,
                      parameter pADDR_WIDTH   = 12,
                      parameter pDATA_WIDTH   = 32
                    )
(
  input  wire                        axi_awvalid,
  input  wire                [14: 0] axi_awaddr,
  input  wire                        axi_arvalid,
  input  wire                [14: 0] axi_araddr,
  input  wire                        axi_wvalid,
  input  wire                 [3: 0] axi_wstrb,
  input  wire  [(pDATA_WIDTH-1) : 0] axi_wdata,
  input  wire                        axi_rready,
  input  wire                        cc_up_enable,
  input  wire                        s_tvalid,
  input  wire  [(pDATA_WIDTH-1) : 0] s_tdata,
  input  wire                 [1: 0] s_tuser,
  input  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] s_tupsb,
  input  wire                 [3: 0] s_tstrb,
  input  wire                 [3: 0] s_tkeep,
  input  wire                        s_tlast,
  input  wire                        m_tready,
  output wire                        axi_awready,
  output wire                        axi_arready,
  output wire                        axi_wready,
  output wire                        axi_rvalid,
  output wire  [(pDATA_WIDTH-1) : 0] axi_rdata,
  output wire                        s_tready,
  output wire                        m_tvalid,
  output wire  [(pDATA_WIDTH-1) : 0] m_tdata,
  output wire                 [1: 0] m_tuser,
  output  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] m_tupsb,
  output wire                 [3: 0] m_tstrb,
  output wire                 [3: 0] m_tkeep,
  output wire                        m_tlast,
  output wire                        low__pri_irq,
  output wire                        high_pri_irq,
  output wire                [23: 0] up_la_data,
  input  wire                        axi_clk,
  input  wire                        axis_clk,
  input  wire                        axi_reset_n,
  input  wire                        axis_rst_n,
  input  wire                        user_clock2,
  input  wire                        uck2_rst_n,
  input  wire                 [4: 0] user_prj_sel
);


wire                         awready_0;
wire                         arready_0;
wire                         wready_0;
wire                         rvalid_0;
wire   [(pDATA_WIDTH-1) : 0] rdata_0;
wire                         awready_1;
wire                         arready_1;
wire                         wready_1;
wire                         rvalid_1;
wire   [(pDATA_WIDTH-1) : 0] rdata_1;
wire                         awready_2;
wire                         arready_2;
wire                         wready_2;
wire                         rvalid_2;
wire   [(pDATA_WIDTH-1) : 0] rdata_2;
wire                         awready_3;
wire                         arready_3;
wire                         wready_3;
wire                         rvalid_3;
wire   [(pDATA_WIDTH-1) : 0] rdata_3;
wire                         awvalid_0_awvalid;
wire                 [11: 0] awaddr;
wire                         arvalid_0_arvalid;
wire                 [11: 0] araddr;
wire                         wvalid_0_wvalid;
wire                  [3: 0] wstrb_0_wstrb;
wire   [(pDATA_WIDTH-1) : 0] wdata;
wire                         rready;
wire                         ss_tvalid_0_ss_tvalid;
wire   [(pDATA_WIDTH-1) : 0] ss_tdata;
wire                  [1: 0] ss_tuser;
wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] ss_tupsb;
wire                  [3: 0] ss_tstrb;
wire                  [3: 0] ss_tkeep;
wire                         ss_tlast;
wire                         sm_tready;
wire                         awvalid_1_awvalid;
wire                         arvalid_1_arvalid;
wire                         wvalid_1_wvalid;
wire                  [3: 0] wstrb_1_wstrb;
wire                         ss_tvalid_1_ss_tvalid;
wire                         awvalid_2_awvalid;
wire                         arvalid_2_arvalid;
wire                         wvalid_2_wvalid;
wire                  [3: 0] wstrb_2_wstrb;
wire                         ss_tvalid_2_ss_tvalid;
wire                         awvalid_3_awvalid;
wire                         arvalid_3_arvalid;
wire                         wvalid_3_wvalid;
wire                  [3: 0] wstrb_3_wstrb;
wire                         ss_tvalid_3_ss_tvalid;
wire                         ss_tready_0;
wire                         ss_tready_1;
wire                         ss_tready_2;
wire                         ss_tready_3;
wire                         sm_tvalid_0;
wire   [(pDATA_WIDTH-1) : 0] sm_tdata_0;
wire                  [2: 0] sm_tid_0;
wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] sm_tupsb_0;
wire                  [3: 0] sm_tstrb_0;
wire                  [3: 0] sm_tkeep_0;
wire                         sm_tlast_0;
wire                         sm_tvalid_1;
wire   [(pDATA_WIDTH-1) : 0] sm_tdata_1;
wire                  [2: 0] sm_tid_1;
wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] sm_tupsb_1;
wire                  [3: 0] sm_tstrb_1;
wire                  [3: 0] sm_tkeep_1;
wire                         sm_tlast_1;
wire                         sm_tvalid_2;
wire   [(pDATA_WIDTH-1) : 0] sm_tdata_2;
wire                  [2: 0] sm_tid_2;
wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] sm_tupsb_2;
wire                  [3: 0] sm_tstrb_2;
wire                  [3: 0] sm_tkeep_2;
wire                         sm_tlast_2;
wire                         sm_tvalid_3;
wire   [(pDATA_WIDTH-1) : 0] sm_tdata_3;
wire                  [2: 0] sm_tid_3;
wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] sm_tupsb_3;
wire                  [3: 0] sm_tstrb_3;
wire                  [3: 0] sm_tkeep_3;
wire                         sm_tlast_3;
wire                         low__pri_irq_0;
wire                         High_pri_req_0;
wire                         low__pri_irq_1;
wire                         High_pri_req_1;
wire                         low__pri_irq_2;
wire                         High_pri_req_2;
wire                         low__pri_irq_3;
wire                         High_pri_req_3;
wire                 [23: 0] la_data_o_la_data_0_0;
wire                 [23: 0] la_data_o_la_data_1_1;
wire                 [23: 0] la_data_o_la_data_2_2;
wire                 [23: 0] la_data_o_la_data_3_3;


// This code snippet was auto generated by xls2vlog.py from source file: ./user_project_wrapper.xlsx
// User: josh
// Date: Sep-22-23



AXIL_SLAV #(.pADDR_WIDTH( 12 ),
            .pDATA_WIDTH( 32 )) U_AXIL_SLAV0 (
                                              .awready_0    (awready_0),               // I  
                                              .arready_0    (arready_0),               // I  
                                              .wready_0     (wready_0),                // I  
                                              .rvalid_0     (rvalid_0),                // I  
                                              .rdata_0      (rdata_0),                 // I  pDATA_WIDTH
                                              .awready_1    (awready_1),               // I  
                                              .arready_1    (arready_1),               // I  
                                              .wready_1     (wready_1),                // I  
                                              .rvalid_1     (rvalid_1),                // I  
                                              .rdata_1      (rdata_1),                 // I  pDATA_WIDTH
                                              .awready_2    (awready_2),               // I  
                                              .arready_2    (arready_2),               // I  
                                              .wready_2     (wready_2),                // I  
                                              .rvalid_2     (rvalid_2),                // I  
                                              .rdata_2      (rdata_2),                 // I  pDATA_WIDTH
                                              .awready_3    (awready_3),               // I  
                                              .arready_3    (arready_3),               // I  
                                              .wready_3     (wready_3),                // I  
                                              .rvalid_3     (rvalid_3),                // I  
                                              .rdata_3      (rdata_3),                 // I  pDATA_WIDTH
                                              .awvalid_0    (awvalid_0_awvalid),       // O  
                                              .awaddr       (awaddr),                  // O  12
                                              .arvalid_0    (arvalid_0_arvalid),       // O  
                                              .araddr       (araddr),                  // O  12
                                              .wvalid_0     (wvalid_0_wvalid),         // O  
                                              .wstrb_0      (wstrb_0_wstrb),           // O  4
                                              .wdata        (wdata),                   // O  pDATA_WIDTH
                                              .rready       (rready),                  // O  
                                              .awvalid_1    (awvalid_1_awvalid),       // O  
                                              .arvalid_1    (arvalid_1_arvalid),       // O  
                                              .wvalid_1     (wvalid_1_wvalid),         // O  
                                              .wstrb_1      (wstrb_1_wstrb),           // O  4
                                              .awvalid_2    (awvalid_2_awvalid),       // O  
                                              .arvalid_2    (arvalid_2_arvalid),       // O  
                                              .wvalid_2     (wvalid_2_wvalid),         // O  
                                              .wstrb_2      (wstrb_2_wstrb),           // O  4
                                              .awvalid_3    (awvalid_3_awvalid),       // O  
                                              .arvalid_3    (arvalid_3_arvalid),       // O  
                                              .wvalid_3     (wvalid_3_wvalid),         // O  
                                              .wstrb_3      (wstrb_3_wstrb),           // O  4
                                              .axi_awvalid  (axi_awvalid),             // I  
                                              .axi_awaddr   (axi_awaddr),              // I  15
                                              .axi_arvalid  (axi_arvalid),             // I  
                                              .axi_araddr   (axi_araddr),              // I  15
                                              .axi_wvalid   (axi_wvalid),              // I  
                                              .axi_wstrb    (axi_wstrb),               // I  4
                                              .axi_wdata    (axi_wdata),               // I  pDATA_WIDTH
                                              .axi_rready   (axi_rready),              // I  
                                              .cc_up_enable (cc_up_enable),            // I  
                                              .axi_awready  (axi_awready),             // O  
                                              .axi_arready  (axi_arready),             // O  
                                              .axi_wready   (axi_wready),              // O  
                                              .axi_rvalid   (axi_rvalid),              // O  
                                              .axi_rdata    (axi_rdata),               // O  pDATA_WIDTH
                                              .axi_clk      (axi_clk),                 // I  
                                              .axi_reset_n  (axi_reset_n),             // I  
                                              .user_prj_sel (user_prj_sel)             // I  5
                                             );


// This code snippet was auto generated by xls2vlog.py from source file: ./user_project_wrapper.xlsx
// User: josh
// Date: Sep-22-23



USER_PRJ0 #(  .pUSER_PROJECT_SIDEBAND_WIDTH ( pUSER_PROJECT_SIDEBAND_WIDTH ), 
        .pADDR_WIDTH( 12 ),
        .pDATA_WIDTH( 32 )) U_USRPRJ0 (
                                          .awready      (awready_0),               // O  
                                          .arready      (arready_0),               // O  
                                          .wready       (wready_0),                // O  
                                          .rvalid       (rvalid_0),                // O  
                                          .rdata        (rdata_0),                 // O  pDATA_WIDTH
                                          .awvalid      (awvalid_0_awvalid),       // I  
                                          .awaddr       (awaddr),                  // I  12
                                          .arvalid      (arvalid_0_arvalid),       // I  
                                          .araddr       (araddr),                  // I  12
                                          .wvalid       (wvalid_0_wvalid),         // I  
                                          .wstrb        (wstrb_0_wstrb),           // I  4
                                          .wdata        (wdata),                   // I  pDATA_WIDTH
                                          .rready       (rready),                  // I  
                                          .ss_tvalid    (ss_tvalid_0_ss_tvalid),   // I  
                                          .ss_tdata     (ss_tdata),                // I  pDATA_WIDTH
                                          .ss_tuser     (ss_tuser),                // I  2

                       .ss_tupsb     (ss_tupsb),                // I  5    

                                          .ss_tstrb     (ss_tstrb),                // I  4
                                          .ss_tkeep     (ss_tkeep),                // I  4
                                          .ss_tlast     (ss_tlast),                // I  
                                          .sm_tready    (sm_tready),               // I  
                                          .ss_tready    (ss_tready_0),             // O  
                                          .sm_tvalid    (sm_tvalid_0),             // O  
                                          .sm_tdata     (sm_tdata_0),              // O  pDATA_WIDTH
                                          .sm_tid       (sm_tid_0),                // O  3

                       .sm_tupsb     (sm_tupsb_0),                // I  5    

                                          .sm_tstrb     (sm_tstrb_0),              // O  4
                                          .sm_tkeep     (sm_tkeep_0),              // O  4 
                                          .sm_tlast     (sm_tlast_0),              // O  
                                          .low__pri_irq (low__pri_irq_0),          // O  
                                          .High_pri_req (High_pri_req_0),          // O  
                                          .la_data_o    (la_data_o_la_data_0_0),   // O  24
                                          .axi_clk      (axi_clk),                 // I  
                                          .axis_clk     (axis_clk),                // I  
                                          .axi_reset_n  (axi_reset_n),             // I  
                                          .axis_rst_n   (axis_rst_n),              // I  
                                          .user_clock2  (user_clock2),             // I  
                                          .uck2_rst_n   (uck2_rst_n)               // I  
                                         );


// This code snippet was auto generated by xls2vlog.py from source file: ./user_project_wrapper.xlsx
// User: josh
// Date: Sep-22-23


USER_PRJ1 #(  .pUSER_PROJECT_SIDEBAND_WIDTH ( pUSER_PROJECT_SIDEBAND_WIDTH ), 
        .pADDR_WIDTH( 12 ),
        .pDATA_WIDTH( 32 )) U_USRPRJ1 (
                                          .awready      (awready_1),               // O  
                                          .arready      (arready_1),               // O  
                                          .wready       (wready_1),                // O  
                                          .rvalid       (rvalid_1),                // O  
                                          .rdata        (rdata_1),                 // O  pDATA_WIDTH
                                          .awvalid      (awvalid_1_awvalid),       // I  
                                          .awaddr       (awaddr),                  // I  12
                                          .arvalid      (arvalid_1_arvalid),       // I  
                                          .araddr       (araddr),                  // I  12
                                          .wvalid       (wvalid_1_wvalid),         // I  
                                          .wstrb        (wstrb_1_wstrb),           // I  4
                                          .wdata        (wdata),                   // I  pDATA_WIDTH
                                          .rready       (rready),                  // I  
                                          .ss_tvalid    (ss_tvalid_1_ss_tvalid),   // I  
                                          .ss_tdata     (ss_tdata),                // I  pDATA_WIDTH
                                          .ss_tuser     (ss_tuser),                // I  2

                       .ss_tupsb     (ss_tupsb),                // I  5    

                                          .ss_tstrb     (ss_tstrb),                // I  4
                                          .ss_tkeep     (ss_tkeep),                // I  4
                                          .ss_tlast     (ss_tlast),                // I  
                                          .sm_tready    (sm_tready),               // I  
                                          .ss_tready    (ss_tready_1),             // O  
                                          .sm_tvalid    (sm_tvalid_1),             // O  
                                          .sm_tdata     (sm_tdata_1),              // O  pDATA_WIDTH
                                          .sm_tid       (sm_tid_1),                // O  3

                       .sm_tupsb     (sm_tupsb_1),                // I  5    

                                          .sm_tstrb     (sm_tstrb_1),              // O  4
                                          .sm_tkeep     (sm_tkeep_1),              // O  4
                                          .sm_tlast     (sm_tlast_1),              // O  
                                          .low__pri_irq (low__pri_irq_1),          // O  
                                          .High_pri_req (High_pri_req_1),          // O  
                                          .la_data_o    (la_data_o_la_data_1_1),   // O  24
                                          .axi_clk      (axi_clk),                 // I  
                                          .axis_clk     (axis_clk),                // I  
                                          .axi_reset_n  (axi_reset_n),             // I  
                                          .axis_rst_n   (axis_rst_n),              // I  
                                          .user_clock2  (user_clock2),             // I  
                                          .uck2_rst_n   (uck2_rst_n)               // I  
                                         );


// This code snippet was auto generated by xls2vlog.py from source file: ./user_project_wrapper.xlsx
// User: josh
// Date: Sep-22-23



USER_PRJ2 #(  .pUSER_PROJECT_SIDEBAND_WIDTH ( pUSER_PROJECT_SIDEBAND_WIDTH ), 
        .pADDR_WIDTH( 12 ),
        .pDATA_WIDTH( 32 )) U_USRPRJ2 (
                                          .awready      (awready_2),               // O  
                                          .arready      (arready_2),               // O  
                                          .wready       (wready_2),                // O  
                                          .rvalid       (rvalid_2),                // O  
                                          .rdata        (rdata_2),                 // O  pDATA_WIDTH
                                          .awvalid      (awvalid_2_awvalid),       // I  
                                          .awaddr       (awaddr),                  // I  12
                                          .arvalid      (arvalid_2_arvalid),       // I  
                                          .araddr       (araddr),                  // I  12
                                          .wvalid       (wvalid_2_wvalid),         // I  
                                          .wstrb        (wstrb_2_wstrb),           // I  4
                                          .wdata        (wdata),                   // I  pDATA_WIDTH
                                          .rready       (rready),                  // I  
                                          .ss_tvalid    (ss_tvalid_2_ss_tvalid),   // I  
                                          .ss_tdata     (ss_tdata),                // I  pDATA_WIDTH
                                          .ss_tuser     (ss_tuser),                // I  2

                       .ss_tupsb     (ss_tupsb),                // I  5    

                                          .ss_tstrb     (ss_tstrb),                // I  4
                                          .ss_tkeep     (ss_tkeep),                // I  4
                                          .ss_tlast     (ss_tlast),                // I  
                                          .sm_tready    (sm_tready),               // I  
                                          .ss_tready    (ss_tready_2),             // O  
                                          .sm_tvalid    (sm_tvalid_2),             // O  
                                          .sm_tdata     (sm_tdata_2),              // O  pDATA_WIDTH
                                          .sm_tid       (sm_tid_2),                // O  3

                       .sm_tupsb     (sm_tupsb_2),                // I  5    

                                          .sm_tstrb     (sm_tstrb_2),              // O  4
                                          .sm_tkeep     (sm_tkeep_2),              // O  4
                                          .sm_tlast     (sm_tlast_2),              // O  
                                          .low__pri_irq (low__pri_irq_2),          // O  
                                          .High_pri_req (High_pri_req_2),          // O  
                                          .la_data_o    (la_data_o_la_data_2_2),   // O  24
                                          .axi_clk      (axi_clk),                 // I  
                                          .axis_clk     (axis_clk),                // I  
                                          .axi_reset_n  (axi_reset_n),             // I  
                                          .axis_rst_n   (axis_rst_n),              // I  
                                          .user_clock2  (user_clock2),             // I  
                                          .uck2_rst_n   (uck2_rst_n)               // I  
                                         );


// This code snippet was auto generated by xls2vlog.py from source file: ./user_project_wrapper.xlsx
// User: josh
// Date: Sep-22-23



USER_PRJ3 #(  .pUSER_PROJECT_SIDEBAND_WIDTH ( pUSER_PROJECT_SIDEBAND_WIDTH ), 
        .pADDR_WIDTH( 12 ),
        .pDATA_WIDTH( 32 )) U_USRPRJ3 (
                                          .awready      (awready_3),               // O  
                                          .arready      (arready_3),               // O  
                                          .wready       (wready_3),                // O  
                                          .rvalid       (rvalid_3),                // O  
                                          .rdata        (rdata_3),                 // O  pDATA_WIDTH
                                          .awvalid      (awvalid_3_awvalid),       // I  
                                          .awaddr       (awaddr),                  // I  12
                                          .arvalid      (arvalid_3_arvalid),       // I  
                                          .araddr       (araddr),                  // I  12
                                          .wvalid       (wvalid_3_wvalid),         // I  
                                          .wstrb        (wstrb_3_wstrb),           // I  4
                                          .wdata        (wdata),                   // I  pDATA_WIDTH
                                          .rready       (rready),                  // I  
                                          .ss_tvalid    (ss_tvalid_3_ss_tvalid),   // I  
                                          .ss_tdata     (ss_tdata),                // I  pDATA_WIDTH
                                          .ss_tuser     (ss_tuser),                // I  2

                       .ss_tupsb     (ss_tupsb),                // I  5    

                                          .ss_tstrb     (ss_tstrb),                // I  4
                                          .ss_tkeep     (ss_tkeep),                // I  4
                                          .ss_tlast     (ss_tlast),                // I  
                                          .sm_tready    (sm_tready),               // I  
                                          .ss_tready    (ss_tready_3),             // O  
                                          .sm_tvalid    (sm_tvalid_3),             // O  
                                          .sm_tdata     (sm_tdata_3),              // O  pDATA_WIDTH
                                          .sm_tid       (sm_tid_3),                // O  3

                       .sm_tupsb     (sm_tupsb_3),                // I  5    

                                          .sm_tstrb     (sm_tstrb_3),              // O  4
                                          .sm_tkeep     (sm_tkeep_3),              // O  4
                                          .sm_tlast     (sm_tlast_3),              // O  
                                          .low__pri_irq (low__pri_irq_3),          // O  
                                          .High_pri_req (High_pri_req_3),          // O  
                                          .la_data_o    (la_data_o_la_data_3_3),   // O  24
                                          .axi_clk      (axi_clk),                 // I  
                                          .axis_clk     (axis_clk),                // I  
                                          .axi_reset_n  (axi_reset_n),             // I  
                                          .axis_rst_n   (axis_rst_n),              // I  
                                          .user_clock2  (user_clock2),             // I  
                                          .uck2_rst_n   (uck2_rst_n)               // I  
                                         );


// This code snippet was auto generated by xls2vlog.py from source file: ./user_project_wrapper.xlsx
// User: josh
// Date: Sep-22-23



AXIS_SLAV #(.pUSER_PROJECT_SIDEBAND_WIDTH ( pUSER_PROJECT_SIDEBAND_WIDTH ), 
      .pADDR_WIDTH( 12 ),
            .pDATA_WIDTH( 32 )) U_AXIS_SLAV0 (
                                              .ss_tvalid_0  (ss_tvalid_0_ss_tvalid),   // O  
                                              .ss_tdata     (ss_tdata),                // O  pDATA_WIDTH
                                              .ss_tuser     (ss_tuser),                // O  2

                          .ss_tupsb     (ss_tupsb),                // O  5    

                                              .ss_tstrb     (ss_tstrb),                // O  4
                                              .ss_tkeep     (ss_tkeep),                // O  4
                                              .ss_tlast     (ss_tlast),                // O  
                                              .ss_tvalid_1  (ss_tvalid_1_ss_tvalid),   // O  
                                              .ss_tvalid_2  (ss_tvalid_2_ss_tvalid),   // O  
                                              .ss_tvalid_3  (ss_tvalid_3_ss_tvalid),   // O  
                                              .ss_tready_0  (ss_tready_0),             // I  
                                              .ss_tready_1  (ss_tready_1),             // I  
                                              .ss_tready_2  (ss_tready_2),             // I  
                                              .ss_tready_3  (ss_tready_3),             // I  
                                              .s_tvalid     (s_tvalid),                // I  
                                              .s_tdata      (s_tdata),                 // I  pDATA_WIDTH
                                              .s_tuser      (s_tuser),                 // I  2

                        .s_tupsb      (s_tupsb),                 // I  4

                                              .s_tstrb      (s_tstrb),                 // I  4
                                              .s_tkeep      (s_tkeep),                 // I  4
                                              .s_tlast      (s_tlast),                 // I  
                                              .s_tready     (s_tready),                // O  
                                              .axis_clk     (axis_clk),                // I  
                                              .axi_reset_n  (axi_reset_n),             // I  
                                              .axis_rst_n   (axis_rst_n),              // I  
                                              .user_prj_sel (user_prj_sel)             // I  5
                                             );


// This code snippet was auto generated by xls2vlog.py from source file: ./user_project_wrapper.xlsx
// User: josh
// Date: Sep-22-23



AXIS_MSTR #(.pUSER_PROJECT_SIDEBAND_WIDTH ( pUSER_PROJECT_SIDEBAND_WIDTH ), 
      .pADDR_WIDTH( 12 ),
            .pDATA_WIDTH( 32 )) U_AXIS_MSTR0 (
                                              .sm_tready    (sm_tready),               // O  
                                              .sm_tvalid_0  (sm_tvalid_0),             // I  
                                              .sm_tdata_0   (sm_tdata_0),              // I  pDATA_WIDTH
                                              .sm_tid_0     (sm_tid_0),                // I  3

                          .sm_tupsb_0     (sm_tupsb_0),                // I  5    

                                              .sm_tstrb_0   (sm_tstrb_0),              // I  4
                                              .sm_tkeep_0   (sm_tkeep_0),              // I  4
                                              .sm_tlast_0   (sm_tlast_0),              // I  
                                              .sm_tvalid_1  (sm_tvalid_1),             // I  
                                              .sm_tdata_1   (sm_tdata_1),              // I  pDATA_WIDTH
                                              .sm_tid_1     (sm_tid_1),                // I  3

                          .sm_tupsb_1     (sm_tupsb_1),                // I  5    

                                              .sm_tstrb_1   (sm_tstrb_1),              // I  4
                                              .sm_tkeep_1   (sm_tkeep_1),              // I  4
                                              .sm_tlast_1   (sm_tlast_1),              // I  
                                              .sm_tvalid_2  (sm_tvalid_2),             // I  
                                              .sm_tdata_2   (sm_tdata_2),              // I  pDATA_WIDTH
                                              .sm_tid_2     (sm_tid_2),                // I  3

                          .sm_tupsb_2     (sm_tupsb_2),                // I  5    

                                              .sm_tstrb_2   (sm_tstrb_2),              // I  4
                                              .sm_tkeep_2   (sm_tkeep_2),              // I  4
                                              .sm_tlast_2   (sm_tlast_2),              // I  
                                              .sm_tvalid_3  (sm_tvalid_3),             // I  
                                              .sm_tdata_3   (sm_tdata_3),              // I  pDATA_WIDTH
                                              .sm_tid_3     (sm_tid_3),                // I  3

                          .sm_tupsb_3     (sm_tupsb_3),                // I  5    

                                              .sm_tstrb_3   (sm_tstrb_3),              // I  4
                                              .sm_tkeep_3   (sm_tkeep_3),              // I  4
                                              .sm_tlast_3   (sm_tlast_3),              // I  
                                              .m_tready     (m_tready),                // I  
                                              .m_tvalid     (m_tvalid),                // O  
                                              .m_tdata      (m_tdata),                 // O  pDATA_WIDTH
                                              .m_tuser      (m_tuser),                 // O  2

                        .m_tupsb      (m_tupsb),                 // O  5

                                              .m_tstrb      (m_tstrb),                 // O  4
                                              .m_tkeep      (m_tkeep),                 // O  4
                                              .m_tlast      (m_tlast),                 // O  
                                              .axis_clk     (axis_clk),                // I  
                                              .axi_reset_n  (axi_reset_n),             // I  
                                              .axis_rst_n   (axis_rst_n),              // I  
                                              .user_prj_sel (user_prj_sel)             // I  5
                                             );


// This code snippet was auto generated by xls2vlog.py from source file: ./user_project_wrapper.xlsx
// User: josh
// Date: Sep-22-23



IRQ_MUX #(.pADDR_WIDTH( 10 )) U_IRQ_MUX0 (
                                          .low__pri_irq_0 (low__pri_irq_0),          // I  
                                          .High_pri_req_0 (High_pri_req_0),          // I  
                                          .low__pri_irq_1 (low__pri_irq_1),          // I  
                                          .High_pri_req_1 (High_pri_req_1),          // I  
                                          .low__pri_irq_2 (low__pri_irq_2),          // I  
                                          .High_pri_req_2 (High_pri_req_2),          // I  
                                          .low__pri_irq_3 (low__pri_irq_3),          // I  
                                          .High_pri_req_3 (High_pri_req_3),          // I  
                                          .low__pri_irq   (low__pri_irq),            // O  
                                          .high_pri_irq   (high_pri_irq),            // O  
                                          .axi_clk        (axi_clk),                 // I  
                                          .axi_reset_n    (axi_reset_n),             // I  
                                          .axis_rst_n     (axis_rst_n),              // I  
                                          .user_prj_sel   (user_prj_sel)             // I  5
                                         );


// This code snippet was auto generated by xls2vlog.py from source file: ./user_project_wrapper.xlsx
// User: josh
// Date: Sep-22-23



LA_MUX #(.pADDR_WIDTH( 12 ),
         .pDATA_WIDTH( 32 )) U_LA_MUX0 (
                                        .la_data_0    (la_data_o_la_data_0_0),   // I  24
                                        .la_data_1    (la_data_o_la_data_1_1),   // I  24
                                        .la_data_2    (la_data_o_la_data_2_2),   // I  24
                                        .la_data_3    (la_data_o_la_data_3_3),   // I  24
                                        .up_la_data   (up_la_data),              // O  24
                                        .axi_clk      (axi_clk),                 // I  
                                        .axis_clk     (axis_clk),                // I  
                                        .axi_reset_n  (axi_reset_n),             // I  
                                        .axis_rst_n   (axis_rst_n),              // I  
                                        .user_prj_sel (user_prj_sel)             // I  5
                                       );




endmodule // USER_SUBSYS


// This code snippet was auto generated by xls2vlog.py from source file: ./user_project_wrapper.xlsx
// User: josh
// Date: Sep-22-23

//`define USE_EDGEDETECT_IP

`timescale 1ns / 10ps

module USER_PRJ0 #(parameter pUSER_PROJECT_SIDEBAND_WIDTH   = 5,
                   parameter pADDR_WIDTH   = 12,
                   parameter pDATA_WIDTH   = 32
                 )
(
  output wire                        awready,
  output wire                        arready,
  output wire                        wready,
  output wire                        rvalid,
  output wire  [(pDATA_WIDTH-1) : 0] rdata,
  input  wire                        awvalid,
  input  wire                [11: 0] awaddr,
  input  wire                        arvalid,
  input  wire                [11: 0] araddr,
  input  wire                        wvalid,
  input  wire                 [3: 0] wstrb,
  input  wire  [(pDATA_WIDTH-1) : 0] wdata,
  input  wire                        rready,
  input  wire                        ss_tvalid,
  input  wire  [(pDATA_WIDTH-1) : 0] ss_tdata,
  input  wire                 [1: 0] ss_tuser,
  input  wire  [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] ss_tupsb,
  input  wire                 [3: 0] ss_tstrb,
  input  wire                 [3: 0] ss_tkeep,
  input  wire                        ss_tlast,
  input  wire                        sm_tready,
  output wire                        ss_tready,
  output wire                        sm_tvalid,
  output wire  [(pDATA_WIDTH-1) : 0] sm_tdata,
  output wire                 [2: 0] sm_tid,
  output  wire [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] sm_tupsb,
  output wire                 [3: 0] sm_tstrb,
  output wire                 [3: 0] sm_tkeep,
  output wire                        sm_tlast,
  output wire                        low__pri_irq,
  output wire                        High_pri_req,
  output wire                [23: 0] la_data_o,
  input  wire                        axi_clk,
  input  wire                        axis_clk,
  input  wire                        axi_reset_n,
  input  wire                        axis_rst_n,
  input  wire                        user_clock2,
  input  wire                        uck2_rst_n
  );

  localparam	RD_IDLE = 1'b0;
  localparam	RD_ADDR_DONE = 1'b1;
   wire sm_tvalid_out;
   assign sm_tvalid=sm_tvalid_out;
  //[TODO] does tlast from FPGA to SOC need send to UP? or use upsb as UP's tlast?
  localparam	FIFO_WIDTH = (pUSER_PROJECT_SIDEBAND_WIDTH + 4 + 4 + 1 + pDATA_WIDTH);		//upsb, tstrb, tkeep, tlast, tdata  

  wire [33:0] dat_in_rsc_dat = {ss_tupsb[1:0], ss_tdata[31:0]};

  wire [33:0] dat_out_rsc_dat;

  wire        ram0_en;
  wire [63:0] ram0_q;
  wire        ram0_we;
  wire [63:0] ram0_d;
  wire [6:0]  ram0_adr;
  wire        ram1_en;
  wire [63:0] ram1_q;
  wire        ram1_we;
  wire [63:0] ram1_d;
  wire [6:0]  ram1_adr;

  reg  [9:0]  reg_widthIn;
  reg  [8:0]  reg_heightIn;
  reg         reg_sw_in;
  reg         reg_rst;
  wire [31:0] crc32_stream_in;
  wire [31:0] crc32_stream_out;
  wire        edgedetect_done;
  reg  [31:0] reg_crc32_stream_in;
  reg  [31:0] reg_crc32_stream_out;
  reg         reg_edgedetect_done;

  wire awvalid_in;
  wire wvalid_in;

  reg [31:0] RegisterData;

  //write addr channel
  assign 	awvalid_in	= awvalid; 
  wire awready_out;
  assign awready = awready_out;

  //write data channel
  assign 	wvalid_in	= wvalid;
  wire wready_out;
  assign wready = wready_out;

  // if both awvalid_in=1 and wvalid_in=1 then output awready_out = 1 and wready_out = 1
  assign awready_out = (awvalid_in && wvalid_in) ? 1 : 0;
  assign wready_out = (awvalid_in && wvalid_in) ? 1 : 0;


  //write register
  always @(posedge axi_clk or negedge axi_reset_n)  begin
    if ( !axi_reset_n ) begin
      reg_widthIn         <= 640;
      reg_heightIn        <= 480;
      reg_sw_in           <= 1;
      reg_rst             <= 0;
    end else begin
      if ( awvalid_in && wvalid_in ) begin		//when awvalid_in=1 and wvalid_in=1 means awready_out=1 and wready_out=1
        if          (awaddr[11:2] == 10'h000 ) begin //offset 0
          if ( wstrb[0] == 1) reg_rst           <= wdata[0];
        end else if (awaddr[11:2] == 10'h001 ) begin //offset 1
          if ( wstrb[0] == 1) reg_widthIn[7:0]  <= wdata[7:0];
          if ( wstrb[1] == 1) reg_widthIn[9:8]  <= wdata[9:8];
        end else if (awaddr[11:2] == 10'h002 ) begin //offset 2
          if ( wstrb[0] == 1) reg_heightIn[7:0] <= wdata[7:0];
          if ( wstrb[1] == 1) reg_heightIn[8]   <= wdata[8];
        end else if (awaddr[11:2] == 10'h003 ) begin //offset 3
          if ( wstrb[0] == 1) reg_sw_in         <= wdata[0];
        end
      end
    end
  end

  always @(posedge axi_clk or negedge axi_reset_n)  begin
    if ( !axi_reset_n ) begin
        reg_edgedetect_done <= 0;
    end else begin
      if (edgedetect_done)
        reg_edgedetect_done <= 1;
      else if ( awvalid_in && wvalid_in ) begin        //when awvalid_in=1 and wvalid_in=1 means awready_out=1 and wready_out=1 
        if (awaddr[11:2] == 10'h006 ) begin //offset 6
          if ( wstrb[0] == 1) reg_edgedetect_done <= 0;
        end
      end
    end
  end


  //read register
  reg [(pDATA_WIDTH-1) : 0] rdata_tmp;
  assign arready = 1; //always assigned to 1, limitation: only support 1T in arvalid, if master issue 2T in arvalid then only 1st raddr is captured.
  reg rvalid_out ;
  assign rvalid = rvalid_out;
  assign rdata =  rdata_tmp;
  reg rd_state;
  reg rd_next_state;
  reg [pADDR_WIDTH-1:0] rd_addr;

  ////
  always @(posedge axi_clk or negedge axi_reset_n)  begin
    if ( !axi_reset_n ) 
      rd_state <= RD_IDLE;
    else
      rd_state <= rd_next_state;
  end

  always@(*)begin
    case(rd_state)
      RD_IDLE:
        if(arvalid && arready) rd_next_state = RD_ADDR_DONE;
        else      rd_next_state = RD_IDLE;
      RD_ADDR_DONE:
        if(rready && rvalid_out) rd_next_state = RD_IDLE;
        else    rd_next_state = RD_ADDR_DONE;
      default:rd_next_state = RD_IDLE;
    endcase
  end 

  always @(posedge axi_clk or negedge axi_reset_n)  begin
    if ( !axi_reset_n ) begin
      rd_addr <= 0;
    rvalid_out <= 0;
    end	
    else begin
      if (rd_state == RD_IDLE )
      if(arvalid && arready) begin
      rd_addr <= araddr;
      rvalid_out <= 1;
      end	
    if (rd_state == RD_ADDR_DONE ) 
      if(rready && rvalid_out)
      rvalid_out <= 0;
    end	
  end

  ////
  always @* begin
    if      (rd_addr[11:2] == 10'h000) rdata_tmp = reg_rst;
    else if (rd_addr[11:2] == 10'h001) rdata_tmp = reg_widthIn;
    else if (rd_addr[11:2] == 10'h002) rdata_tmp = reg_heightIn;
    else if (rd_addr[11:2] == 10'h003) rdata_tmp = reg_sw_in;
    else if (rd_addr[11:2] == 10'h004) rdata_tmp = reg_crc32_stream_in;
    else if (rd_addr[11:2] == 10'h005) rdata_tmp = reg_crc32_stream_out;
    else if (rd_addr[11:2] == 10'h006) rdata_tmp = reg_edgedetect_done;
    else                              rdata_tmp = 0;
  end

  //DUT
  assign sm_tdata  = dat_out_rsc_dat[31: 0]; 

  assign sm_tupsb = dat_out_rsc_dat[33:32];


  assign sm_tlast = dat_out_rsc_dat[33];
  assign {sm_tstrb, sm_tkeep} = 0;

  wire dat_in_rsc_rdy;

  assign ss_tready = dat_in_rsc_rdy;

  always @(posedge axi_clk or negedge axi_reset_n)  begin
    if ( !axi_reset_n ) begin
      reg_crc32_stream_in  <= 0;
      reg_crc32_stream_out <= 0;
    end else if (edgedetect_done) begin
      reg_crc32_stream_in  <= crc32_stream_in ;
      reg_crc32_stream_out <= crc32_stream_out;
    end
  end

  EdgeDetect_Top U_EdgeDetect (
  .clk                     (axi_clk           ), //user_clock2 ?
  .rst                     (reg_rst           ), 
  .arst_n                  (axi_reset_n       ), //~uck2_rst_n ? 
  .widthIn                 (reg_widthIn       ), //I 
  .heightIn                (reg_heightIn      ), //I
  .sw_in                   (reg_sw_in         ), //I
  .crc32_pix_in_rsc_dat    (crc32_stream_in   ), //O
  .crc32_pix_in_triosy_lz  (),                   //O, not useful
  .crc32_dat_out_rsc_dat   (crc32_stream_out  ), //O
  .crc32_dat_out_triosy_lz (edgedetect_done   ), //O
  .dat_in_rsc_dat          (dat_in_rsc_dat    ), //I
  .dat_in_rsc_vld          (ss_tvalid         ), //I
  .dat_in_rsc_rdy          (dat_in_rsc_rdy    ), //O
  .dat_out_rsc_dat         (dat_out_rsc_dat   ), //O
  .dat_out_rsc_vld         (sm_tvalid_out     ), //O
  .dat_out_rsc_rdy         (sm_tready         ), //I
  .line_buf0_rsc_en        (ram0_en           ), //O
  .line_buf0_rsc_q         (ram0_q            ), //I
  .line_buf0_rsc_we        (ram0_we           ), //O
  .line_buf0_rsc_d         (ram0_d            ), //O
  .line_buf0_rsc_adr       (ram0_adr          ), //O
  .line_buf1_rsc_en        (ram1_en           ), //O
  .line_buf1_rsc_q         (ram1_q            ), //I 
  .line_buf1_rsc_we        (ram1_we           ), //O 
  .line_buf1_rsc_d         (ram1_d            ), //O 
  .line_buf1_rsc_adr       (ram1_adr          )  //O
  );


  ra1shd80x64m4h3v2 U_SPRAM_0(
    .A   (ram0_adr ), 
    .D   (ram0_d   ), 
    .CEN (~ram0_en  ), 
    .WEN (~ram0_we  ), 
    .OEN (1'b0     ), 
    .CLK (axi_clk  ), //user_clock2 ? 
    .Q   (ram0_q   )
    );


  ra1shd80x64m4h3v2 U_SPRAM_1(
    .A   (ram1_adr ), 
    .D   (ram1_d   ), 
    .CEN (~ram1_en  ), 
    .WEN (~ram1_we  ), 
    .OEN (1'b0     ), 
    .CLK (axi_clk  ), //user_clock2 ? 
    .Q   (ram1_q   )
    );
  //~

// 24 bit 
// [23:16] for axi-lite interface; [15:12] for axi-stream interface;
assign la_data_o[23:16] = {awvalid,awready_out,wvalid,wready_out,arvalid,1'b1,rready,rvalid_out};
assign la_data_o[15:12] = {ss_tvalid,dat_in_rsc_rdy,sm_tvalid_out,sm_tready};
assign la_data_o[11:8]=wdata[3:0];
assign la_data_o[7:4]=ss_tdata[3:0];
assign la_data_o[3:0]=dat_out_rsc_dat[3:0];


endmodule //USER_PRJ0





module USER_PRJ1 #( parameter pUSER_PROJECT_SIDEBAND_WIDTH   = 5,
          parameter pADDR_WIDTH   = 12,
                   parameter pDATA_WIDTH   = 32
                 )
(
  output wire                        awready,
  output wire                        arready,
  output wire                        wready,
  output wire                        rvalid,
  output wire  [(pDATA_WIDTH-1) : 0] rdata,
  input  wire                        awvalid,
  input  wire                [11: 0] awaddr,
  input  wire                        arvalid,
  input  wire                [11: 0] araddr,
  input  wire                        wvalid,
  input  wire                 [3: 0] wstrb,
  input  wire  [(pDATA_WIDTH-1) : 0] wdata,
  input  wire                        rready,
  input  wire                        ss_tvalid,
  input  wire  [(pDATA_WIDTH-1) : 0] ss_tdata,
  input  wire                 [1: 0] ss_tuser,
  input  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] ss_tupsb,
  input  wire                 [3: 0] ss_tstrb,
  input  wire                 [3: 0] ss_tkeep,
  input  wire                        ss_tlast,
  input  wire                        sm_tready,
  output wire                        ss_tready,
  output wire                        sm_tvalid,
  output wire  [(pDATA_WIDTH-1) : 0] sm_tdata,
  output wire                 [2: 0] sm_tid,
  output  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] sm_tupsb,
  output wire                 [3: 0] sm_tstrb,
  output wire                 [3: 0] sm_tkeep,
  output wire                        sm_tlast,
  output wire                        low__pri_irq,
  output wire                        High_pri_req,
  output wire                [23: 0] la_data_o,
  input  wire                        axi_clk,
  input  wire                        axis_clk,
  input  wire                        axi_reset_n,
  input  wire                        axis_rst_n,
  input  wire                        user_clock2,
  input  wire                        uck2_rst_n
);

////////////////////////// axi- lite part


wire awvalid_in;
wire wvalid_in;

//write addr channel
assign awvalid_in	= awvalid; 
wire awready_out;
assign awready = awready_out;

//write data channel
assign 	wvalid_in	= wvalid;
wire wready_out;
assign wready = wready_out;

// if both awvalid_in=1 and wvalid_in=1 then output awready_out = 1 and wready_out = 1
assign awready_out = (awvalid_in && wvalid_in) ? 1 : 0;
assign wready_out = (awvalid_in && wvalid_in) ? 1 : 0;

wire ss_tready_out;
assign ss_tready=ss_tready_out;


wire sm_tvalid_out;
assign sm_tvalid = sm_tvalid_out;

wire [31:0] sm_tdata_out;
assign sm_tdata  = sm_tdata_out;

//write register   // to let RESET State go back to Command state
/*always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) begin
    reg_ap_control         <= 0;

  end else begin
    if ( awvalid_in && wvalid_in ) begin		//when awvalid_in=1 and wvalid_in=1 means awready_out=1 and wready_out=1
       if  (awaddr[11:0] == 12'h000 ) begin //offset 0
      
       end 
       else begin
       end
    end
  end
end
*/
localparam	RD_IDLE = 1'b0;
localparam	RD_ADDR_DONE = 1'b1;
localparam	Command   = 4'd0;
localparam	IN_COPY   = 4'd1;
localparam	OUT_COPY  = 4'd2;
localparam	RESET     = 4'd3;
localparam	F_WAIT1    = 4'd1;
localparam	F_OUT1     = 4'd2;
localparam	F_OUT2     = 4'd3;
localparam	U_OUT      = 4'd4;
reg [3:0] state,next_state;
//read register
reg [(pDATA_WIDTH-1) : 0] rdata_tmp;
assign arready = 1; //always assigned to 1, limitation: only support 1T in arvalid, if master issue 2T in arvalid then only 1st raddr is captured.
reg rvalid_out ;
assign rvalid = rvalid_out;
assign rdata =  rdata_tmp;
reg rd_state;
reg rd_next_state;
reg [pADDR_WIDTH-1:0] rd_addr;
reg [3:0] Out_state,next_Out_state;
////
always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) 
    rd_state <= RD_IDLE;
  else
    rd_state <= rd_next_state;
end



always@(*)begin
  case(rd_state)
    RD_IDLE:
      if(arvalid && arready) rd_next_state = RD_ADDR_DONE;
      else      rd_next_state = RD_IDLE;
    RD_ADDR_DONE:
      if(rready && rvalid_out) rd_next_state = RD_IDLE;
      else    rd_next_state = RD_ADDR_DONE;
    default:rd_next_state = RD_IDLE;
  endcase
end 

always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) begin
        rd_addr <= 0;
	      rvalid_out <= 0;
  end	
  else begin
    if (rd_state == RD_IDLE )
	  if(arvalid && arready) begin
		rd_addr <= araddr;
		rvalid_out <= 1;
	  end	
	if (rd_state == RD_ADDR_DONE ) 
	  if(rready && rvalid_out)
		rvalid_out <= 0;
  end	
end

////
always @* begin
  if      (rd_addr[11:0] == 12'h000) rdata_tmp = (state==RESET);
  else                               rdata_tmp = 0;
end


assign sm_tid        = 3'b0;
assign sm_tupsb      = 5'b0;
assign sm_tstrb      = 4'b0;
assign sm_tkeep      = 1'b0;
assign low__pri_irq  = 1'b0;
assign High_pri_req  = 1'b0;

// 24 bit 
// [23:16] for axi-lite interface; [15:12] for axi-stream interface; [11:8] for state; [7:4] for Out_state; [3:0] for data;
assign la_data_o[23:16] = {awvalid,awready_out,wvalid,wready_out,arvalid,1'b1,rready,rvalid_out};
assign la_data_o[15:12] = {ss_tvalid,ss_tready_out,sm_tvalid_out,sm_tready};
assign la_data_o[11:8]=state;
assign la_data_o[7:4]=Out_state;
assign la_data_o[3:0]={wdata[0],ss_tdata[0],sm_tdata_out[0],1'b0};

wire        in_ramf_en;
wire [63:0] in_ramf_q;
wire        in_ramf_we;
wire [63:0] in_ramf_d;
wire [9:0]  in_ramf_adr;

wire        in_ramu_en;
wire [15:0] in_ramu_q;
wire        in_ramu_we;
wire [15:0] in_ramu_d;
wire [9:0]  in_ramu_adr;

wire        out_ramf_en;
wire [63:0] out_ramf_q;
wire        out_ramf_we;
wire [63:0] out_ramf_d;
wire [9:0]  out_ramf_adr;

wire        out_ramu_en;
wire [15:0] out_ramu_q;
wire        out_ramu_we;
wire [15:0] out_ramu_d;
wire [9:0]  out_ramu_adr;

wire        ram0_en;
wire [63:0] ram0_q;
wire        ram0_we;
wire [63:0] ram0_d;
wire [9:0]  ram0_adr;

wire        ram1_en;
wire [63:0] ram1_q;
wire        ram1_we;
wire [63:0] ram1_d;
wire [9:0]  ram1_adr;

wire [63:0] In_data;
wire In_vld;
wire In_rdy;	
wire [9:0] Inram_adr;
wire [63:0] Inram_d;
wire Inram_we;
reg reg_rst_incpopy;
reg reg_rst_out_stage;
reg [31:0]regx_data;
reg [31:0]regy_data;
reg [15:0]reg_mode1_in;

assign ss_tready_out=(state==Command)?1'b1:(state==IN_COPY)?In_rdy:1'b0;
assign In_vld=(state==IN_COPY)?ss_tvalid:1'b0;

In_copy In_copy (
  .clk(axi_clk), 
  .rst(reg_rst_incpopy), 
  .arst_n(axi_reset_n),
  .in_data_rsc_dat(ss_tdata),
  .in_data_rsc_vld(In_vld), //I
  .in_data_rsc_rdy(In_rdy), 
  .qin_rsc_adr(Inram_adr),
  .qin_rsc_d(Inram_d),
  .qin_rsc_we(Inram_we),
  .qin_rsc_q(),
  .qin_rsc_en(Inram_en),
  .qin_triosy_lz(),
  .ap_done_rsc_dat(), 
  .ap_done_rsc_vld(In_copy_done),
  .ap_done_rsc_rdy(1'b1),
  .ap_start_rsc_dat(1'b1),
  .ap_start_rsc_vld(state==IN_COPY),
  .ap_start_rsc_rdy(),
  .mode_rsc_dat(reg_mode1_in==2||reg_mode1_in==3)
);

wire ap_done_vld;     
wire ap_done_rdy;     

wire Out_vld;

always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) begin
    state <= 4'b0;
  end
  else begin
    state <= next_state;
  end
end

wire Out_copy_done;

always@(*)begin
  case(state)
    Command:   
    	if(ss_tvalid && ss_tdata[3:2]==2'b01) next_state = IN_COPY;
   		else next_state = Command;
    IN_COPY:   
    	if(In_copy_done) next_state = OUT_COPY;
   		else next_state = IN_COPY;
    OUT_COPY:  
    	if(Out_copy_done) next_state=RESET;
   		else next_state=OUT_COPY;
    RESET:
    	if(awvalid_in && wvalid_in &&(awaddr[11:0] == 12'h000)&&(wdata[0]==1)) next_state=Command;
     	else next_state = RESET;
    default:next_state = Command;
  endcase
end 

reg reg_rst;

always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) begin
    reg_mode1_in <= 16'b0;
  end
  else begin
    if(state==Command)begin
      reg_mode1_in <= {14'b0,ss_tdata[1:0]};
    end
    else begin
      reg_mode1_in <=reg_mode1_in;
    end
  end
end

always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) begin 
    Out_state <= 2'b0;
  end
  else begin
  	Out_state <= next_Out_state;
  end
end

always@(*)begin
  case(Out_state)
    Command: 
    	if(ss_tvalid && ss_tdata[3:2]==2'b01 && (ss_tdata[1:0]==2'd0 || ss_tdata[1:0]== 2'd1))  next_Out_state = F_WAIT1;
    	else if(ss_tvalid && ss_tdata[3:2]==2'b01 && (ss_tdata[1:0]==2'd2 || ss_tdata[1:0]==2'd3))  next_Out_state = U_OUT;
    	else next_Out_state=Command;
    	
    F_WAIT1:
    	if(Out_copy_done)next_Out_state = Command;
			else if(Out_vld)next_Out_state = F_OUT1;
    	else next_Out_state = F_WAIT1;
    	
    F_OUT1: 
    	if(sm_tready) next_Out_state = F_OUT2;
    	else next_Out_state = F_OUT1;
    	
    F_OUT2: 
    	if(sm_tready) next_Out_state = F_WAIT1;
    	else next_Out_state = F_OUT2;
    	
    U_OUT:    
    	if(Out_copy_done)next_Out_state = Command;
    	else next_Out_state = U_OUT;
    	
    default:next_Out_state=Command;
  endcase
end 

wire [79:0] Out_data;

always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) begin
		regx_data <= 32'b0;
		regy_data <= 32'b0;
  end
  else begin
  	if(Out_state==F_WAIT1 && Out_vld)begin
			regx_data <= Out_data[31:0];
			regy_data <= Out_data[63:32];
 	  end
 	  else begin
      regx_data <= regx_data;
			regy_data <= regy_data;
 	  end
  end
end

/********** sm_tlast ***********/

reg [11:0] last_cnt;
always @(posedge axi_clk or negedge axi_reset_n)  begin
  if ( !axi_reset_n ) begin
		last_cnt <= 12'b0;
  end
  else begin
    if(state==RESET) last_cnt <= 12'b0;
    else begin
      if(((Out_state==U_OUT) ? Out_vld : (Out_state==F_OUT1||Out_state==F_OUT2))&sm_tready) last_cnt<=last_cnt+12'b1;
      else last_cnt<=last_cnt;
 	  end
  end
end




assign sm_tlast  = (reg_mode1_in[1])  ? ((last_cnt==12'd1023) ? 1 : 0) : ((last_cnt==12'd2047) ? 1 : 0);
assign sm_tvalid_out=(Out_state==U_OUT) ? Out_vld : (Out_state==F_OUT1||Out_state==F_OUT2);
assign sm_tdata_out=(Out_state==U_OUT) ? {16'b0,Out_data[79:64]} : ((Out_state==F_OUT1)?regx_data:regy_data);
assign Out_rdy   = (Out_state==U_OUT||Out_state==F_OUT2) ? sm_tready : 0;




fiFFNTT fiFFNTT(
.clk(axi_clk),          // I
.rst(reg_rst),          // I
.arst_n(axi_reset_n),   // I
.ap_start_rsc_dat(1'b1),// I
.ap_start_rsc_vld(state==OUT_COPY),    // I
.ap_start_rsc_rdy(),    // O
.ap_done_rsc_dat(),     // O
.ap_done_rsc_vld(Out_copy_done), // O
.ap_done_rsc_rdy(1'b1),     // I
.mode1_rsc_dat(reg_mode1_in),  //I 16
.mode1_triosy_lz(), 
.in_f_d_rsc_adr(in_ramf_adr),  // O 10
.in_f_d_rsc_d(in_ramf_d),    // O 64
.in_f_d_rsc_we(in_ramf_we),   // O 1 
.in_f_d_rsc_q(in_ramf_q),    // I 64
.in_f_d_rsc_en(in_ramf_en),   // O 1
.in_f_d_triosy_lz(), 
.in_u_rsc_adr(in_ramu_adr), // O 10
.in_u_rsc_d(in_ramu_d),   // O 16
.in_u_rsc_we(in_ramu_we),  // O
.in_u_rsc_q(in_ramu_q),   // I 16
.in_u_rsc_en(in_ramu_en),  // O 
.in_u_triosy_lz(),
.out_f_d_rsc_adr(out_ramf_adr),
.out_f_d_rsc_d(out_ramf_d),
.out_f_d_rsc_we(out_ramf_we),
.out_f_d_rsc_q(out_ramf_q), 
.out_f_d_rsc_en(out_ramf_en),
.out_f_d_triosy_lz(),
.out_u_rsc_adr(out_ramu_adr), 
.out_u_rsc_d(out_ramu_d),
.out_u_rsc_we(out_ramu_we), 
.out_u_rsc_q(out_ramu_q),
.out_u_rsc_en(out_ramu_en),
.out_u_triosy_lz(),
.out1_rsc_dat(Out_data),//O,80 bit{16'b,64'b},
.out1_rsc_vld(Out_vld),//O;
.out1_rsc_rdy(Out_rdy)
);






wire mux_state;
assign mux_state=!(reg_mode1_in==2||reg_mode1_in==3);
assign ram0_en   = (state==IN_COPY)?Inram_en  : ((mux_state)? in_ramf_en:in_ramu_en);
assign ram0_we   = (state==IN_COPY)?Inram_we  : ((mux_state)? in_ramf_we:in_ramu_we);
assign ram0_adr  = (state==IN_COPY)?Inram_adr : ((mux_state)? in_ramf_adr:in_ramu_adr);
assign ram0_d    = (state==IN_COPY)?Inram_d   : ((mux_state)? in_ramf_d:{48'b0,in_ramu_d});
assign in_ramu_q = ram0_q[15:0];
assign in_ramf_q = ram0_q;


assign ram1_en  	= (mux_state) ? out_ramf_en  : out_ramu_en;
assign ram1_we  	= (mux_state) ? out_ramf_we  : out_ramu_we;
assign ram1_adr 	= (mux_state) ? out_ramf_adr : out_ramu_adr;
assign ram1_d   	= (mux_state) ? out_ramf_d   : {48'b0,out_ramu_d};
assign out_ramu_q = ram1_q[15:0];
assign out_ramf_q = ram1_q;


ra1shd1024x64m4h3v2 SRAM0(
  .CLK(axi_clk),
  .WEN(~ram0_we),
  .OEN(1'b0),
  .CEN(~ram0_en),
  .A(ram0_adr),
  .D(ram0_d),
  .Q(ram0_q)
);

ra1shd1024x64m4h3v2 SRAM1(
  .CLK(axi_clk),
  .WEN(~ram1_we),
  .OEN(1'b0),
  .CEN(~ram1_en),
  .A(ram1_adr),
  .D(ram1_d),
  .Q(ram1_q)
);


endmodule 


// This code snippet was auto generated by xls2vlog.py from source file: ./user_project_wrapper.xlsx
// User: josh
// Date: Sep-22-23



module USER_PRJ2 #( parameter pUSER_PROJECT_SIDEBAND_WIDTH   = 5,
          parameter pADDR_WIDTH   = 12,
                   parameter pDATA_WIDTH   = 32
                 )
(
  output wire                        awready,
  output wire                        arready,
  output wire                        wready,
  output wire                        rvalid,
  output wire  [(pDATA_WIDTH-1) : 0] rdata,
  input  wire                        awvalid,
  input  wire                [11: 0] awaddr,
  input  wire                        arvalid,
  input  wire                [11: 0] araddr,
  input  wire                        wvalid,
  input  wire                 [3: 0] wstrb,
  input  wire  [(pDATA_WIDTH-1) : 0] wdata,
  input  wire                        rready,
  input  wire                        ss_tvalid,
  input  wire  [(pDATA_WIDTH-1) : 0] ss_tdata,
  input  wire                 [1: 0] ss_tuser,
  input  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] ss_tupsb,
  input  wire                 [3: 0] ss_tstrb,
  input  wire                 [3: 0] ss_tkeep,
  input  wire                        ss_tlast,
  input  wire                        sm_tready,
  output wire                        ss_tready,
  output wire                        sm_tvalid,
  output wire  [(pDATA_WIDTH-1) : 0] sm_tdata,
  output wire                 [2: 0] sm_tid,
  output  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] sm_tupsb,
  output wire                 [3: 0] sm_tstrb,
  output wire                 [3: 0] sm_tkeep,
  output wire                        sm_tlast,
  output wire                        low__pri_irq,
  output wire                        High_pri_req,
  output wire                [23: 0] la_data_o,
  input  wire                        axi_clk,
  input  wire                        axis_clk,
  input  wire                        axi_reset_n,
  input  wire                        axis_rst_n,
  input  wire                        user_clock2,
  input  wire                        uck2_rst_n
);


assign awready       = 1'b0;
assign arready       = 1'b0;
assign wready        = 1'b0;
assign rvalid        = 1'b0;
assign rdata         = {pDATA_WIDTH{1'b0}};
assign ss_tready     = 1'b0;
assign sm_tvalid     = 1'b0;
assign sm_tdata      = {pDATA_WIDTH{1'b0}};
assign sm_tid        = 3'b0;
assign sm_tupsb      = 5'b0;
assign sm_tstrb      = 4'b0;
assign sm_tkeep      = 1'b0;
assign sm_tlast      = 1'b0;
assign low__pri_irq  = 1'b0;
assign High_pri_req  = 1'b0;
assign la_data_o     = 24'b0;


endmodule // USER_PRJ2
// This code snippet was auto generated by xls2vlog.py from source file: ./user_project_wrapper.xlsx
// User: josh
// Date: Sep-22-23



module USER_PRJ3 #( parameter pUSER_PROJECT_SIDEBAND_WIDTH   = 5,
          parameter pADDR_WIDTH   = 12,
                   parameter pDATA_WIDTH   = 32
                 )
(
  output wire                        awready,
  output wire                        arready,
  output wire                        wready,
  output wire                        rvalid,
  output wire  [(pDATA_WIDTH-1) : 0] rdata,
  input  wire                        awvalid,
  input  wire                [11: 0] awaddr,
  input  wire                        arvalid,
  input  wire                [11: 0] araddr,
  input  wire                        wvalid,
  input  wire                 [3: 0] wstrb,
  input  wire  [(pDATA_WIDTH-1) : 0] wdata,
  input  wire                        rready,
  input  wire                        ss_tvalid,
  input  wire  [(pDATA_WIDTH-1) : 0] ss_tdata,
  input  wire                 [1: 0] ss_tuser,
  input  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] ss_tupsb,
  input  wire                 [3: 0] ss_tstrb,
  input  wire                 [3: 0] ss_tkeep,
  input  wire                        ss_tlast,
  input  wire                        sm_tready,
  output wire                        ss_tready,
  output wire                        sm_tvalid,
  output wire  [(pDATA_WIDTH-1) : 0] sm_tdata,
  output wire                 [2: 0] sm_tid,
  output  wire                 [pUSER_PROJECT_SIDEBAND_WIDTH-1: 0] sm_tupsb,
  output wire                 [3: 0] sm_tstrb,
  output wire                 [3: 0] sm_tkeep,
  output wire                        sm_tlast,
  output wire                        low__pri_irq,
  output wire                        High_pri_req,
  output wire                [23: 0] la_data_o,
  input  wire                        axi_clk,
  input  wire                        axis_clk,
  input  wire                        axi_reset_n,
  input  wire                        axis_rst_n,
  input  wire                        user_clock2,
  input  wire                        uck2_rst_n
);


assign awready       = 1'b0;
assign arready       = 1'b0;
assign wready        = 1'b0;
assign rvalid        = 1'b0;
assign rdata         = {pDATA_WIDTH{1'b0}};
assign ss_tready     = 1'b0;
assign sm_tvalid     = 1'b0;
assign sm_tdata      = {pDATA_WIDTH{1'b0}};
assign sm_tid        = 3'b0;
assign sm_tupsb      = 5'b0;
assign sm_tstrb      = 4'b0;
assign sm_tkeep      = 1'b0;
assign sm_tlast      = 1'b0;
assign low__pri_irq  = 1'b0;
assign High_pri_req  = 1'b0;
assign la_data_o     = 24'b0;


endmodule // USER_PRJ3

//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_in_wait_coupled_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_coupled_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

// same as falcon
// module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

//   parameter integer rscid = 1;
//   parameter integer width = 8;

//   output [width-1:0] idat;
//   output             rdy;
//   output             ivld;
//   input  [width-1:0] dat;
//   input              irdy;
//   input              vld;

//   wire   [width-1:0] idat;
//   wire               rdy;
//   wire               ivld;

//   localparam stallOff = 0; 
//   wire                  stall_ctrl;
//   assign stall_ctrl = stallOff;

//   assign idat = dat;
//   assign rdy = irdy && !stall_ctrl;
//   assign ivld = vld && !stall_ctrl;

// endmodule


//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

// same as falcon
// module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

//   parameter integer rscid = 1;
//   parameter integer width = 8;

//   output [width-1:0] dat;
//   output             irdy;
//   output             vld;
//   input  [width-1:0] idat;
//   input              rdy;
//   input              ivld;

//   wire   [width-1:0] dat;
//   wire               irdy;
//   wire               vld;

//   localparam stallOff = 0; 
//   wire stall_ctrl;
//   assign stall_ctrl = stallOff;

//   assign dat = idat;
//   assign irdy = rdy && !stall_ctrl;
//   assign vld = ivld && !stall_ctrl;

// endmodule



//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

// same as falcon
// module mgc_io_sync_v2 (ld, lz);
//     parameter valid = 0;

//     input  ld;
//     output lz;

//     wire   lz;

//     assign lz = ld;

// endmodule


//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_genreg_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_genreg_v1 (clk, en, arst, srst, d, z);
    parameter integer width   = 1;
    parameter integer ph_clk  = 1;
    parameter integer ph_en   = 1;
    parameter integer ph_arst = 0;
    parameter integer ph_srst = 1;
    parameter         has_en  = 1'b1;

    input clk;
    input en;
    input arst;
    input srst;
    input      [width-1:0] d;
    output reg [width-1:0] z;

    //  Generate parameters
    //  ph_clk | ph_arst | has_en     Label:
    //    1        1          1       GEN_CLK1_ARST1_EN1
    //    1        1          0       GEN_CLK1_ARST1_EN0
    //    1        0          1       GEN_CLK1_ARST0_EN1
    //    1        0          0       GEN_CLK1_ARST0_EN0
    //    0        1          1       GEN_CLK0_ARST1_EN1
    //    0        1          0       GEN_CLK0_ARST1_EN0
    //    0        0          1       GEN_CLK0_ARST0_EN1
    //    0        0          0       GEN_CLK0_ARST0_EN0
    
    generate 
      // Pos edge clock, pos edge async reset, has enable
      if (ph_clk == 1 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK1_ARST1_EN1
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST1_EN1

      // Pos edge clock, pos edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK1_ARST1_EN0
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST1_EN0

      // Pos edge clock, neg edge async reset, has enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK1_ARST0_EN1
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST0_EN1

      // Pos edge clock, neg edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK1_ARST0_EN0
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST0_EN0


      // Neg edge clock, pos edge async reset, has enable
      if (ph_clk == 0 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK0_ARST1_EN1
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST1_EN1

      // Neg edge clock, pos edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK0_ARST1_EN0
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST1_EN0

      // Neg edge clock, neg edge async reset, has enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK0_ARST0_EN1
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST0_EN1

      // Neg edge clock, neg edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK0_ARST0_EN0
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST0_EN0
    endgenerate
endmodule


//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_fifo_wait_core_v5.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

/*
 *            _________________________________________________
 * WRITER    |                                                 |   READER
 *           |               ccs_fifo_wait_core                |
 *           |             _____________________               |
 *        --<|  din_rdy --<|  ---------------- <|--- dout_rdy <|---
 *           |             |       FIFO         |              |
 *        ---|> din_vld ---|> ----------------  |>-- dout_vld  |>--
 *        ---|>     din ---|> ----------------  |>-- dout      |>--
 *           |             |____________________|              |
 *           |_________________________________________________|
 *
 *    rdy    - can be considered as a notFULL signal
 *    vld    - can be considered as a notEMPTY signal
 *    is_idle - clk can be safely gated
 *
 * Change History:
 *    2019-01-24 - Add assertion to verify rdy signal behavior under reset.
 *                 Fix bug in that behavior.
 */

module ccs_fifo_wait_core_v5 (clk, en, arst, srst, din_vld, din_rdy, din, dout_vld, dout_rdy, dout, sd, is_idle);

    parameter integer rscid    = 0;     // resource ID
    parameter integer width    = 8;     // fifo width
    parameter integer sz_width = 8;     // size of port for elements in fifo
    parameter integer fifo_sz  = 8;     // fifo depth
    parameter integer ph_clk   = 1;     // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1;     // clock enable polarity
    parameter integer ph_arst  = 1;     // async reset polarity
    parameter integer ph_srst  = 1;     // sync reset polarity
    parameter integer ph_log2  = 3;     // log2(fifo_sz)

    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 din_vld;    // writer has valid data
    output                din_rdy;    // fifo ready for data (not full)
    input  [width-1:0]    din;
    output                dout_vld;   // fifo has valid data (not empty)
    input                 dout_rdy;   // reader ready for data
    output [width-1:0]    dout;
    output [sz_width-1:0] sd;
    output                is_idle;

    localparam integer fifo_b  = width * fifo_sz;
    localparam integer fifo_mx = (fifo_sz > 0) ? (fifo_sz-1) : 0 ;
    localparam integer fifo_mx_over_8 = fifo_mx / 8 ;

    reg      [fifo_mx:0] stat_pre;
    wire     [fifo_mx:0] stat;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    wire     [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    reg      [fifo_mx:0] en_l;
    reg      [fifo_mx_over_8:0] en_l_s;

    reg      [width-1:0] buff_nxt;

    reg                  stat_nxt;
    reg                  stat_behind;
    reg                  stat_ahead;
    reg                  stat_tail;
    reg                  en_l_var;

    integer              i;
    genvar               eni;

    wire [32:0]          size_t;
    reg  [31:0]          count;
    reg  [31:0]          count_t;
    reg  [32:0]          n_elem;
    wire                 din_rdy_drv;
    wire                 dout_vld_drv;
    wire                 din_vld_int;
    wire                 hs_init;
    wire                 active;
    wire                 is_idle_drv;

    // synopsys translate_off
    reg  [31:0]          peak;
    initial
    begin
      peak  = 32'b0;
    end
    // synopsys translate_on

    assign din_rdy = din_rdy_drv;
    assign dout_vld = dout_vld_drv;
    assign is_idle = is_idle_drv;

    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
      assign din_vld_int = din_vld & hs_init;
      assign din_rdy_drv = (dout_rdy | (~stat[0])) & hs_init;
      assign dout_vld_drv = din_vld_int | stat[fifo_sz-1];

      assign active = (din_vld_int & din_rdy_drv) | (dout_rdy & dout_vld_drv);
      assign is_idle_drv = (~active) & hs_init;

      assign size_t = (count - {31'b0, (dout_rdy & stat[fifo_sz-1])}) + {31'b0, din_vld_int};
      assign sd = size_t[sz_width-1:0];

      assign dout = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : din;

      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          stat_behind = (i != 0) ? stat[i-1] : 1'b0;
          stat_ahead  = (i != (fifo_sz-1)) ? stat[i+1] : 1'b1;

          // Determine if this buffer element will have data
          stat_nxt = stat_ahead &                       // valid element ahead of this one (or head)
                       (stat_behind                     // valid element behind this one
                         | (stat[i] & (~dout_rdy))      // valid element and output not ready (in use and not shifted)
                         | (stat[i] & din_vld_int)      // valid element and input has data
                         | (din_vld_int & (~dout_rdy))  // input has data and output not ready
                       );
          stat_pre[i] = stat_nxt;

          // First empty elem when not shifting or last valid elem after shifting (assumes stat_behind == 0)
          stat_tail = stat_ahead & (((~stat[i]) & (~dout_rdy)) | (stat[i] & dout_rdy));

          if (dout_rdy & stat_behind)
          begin
            // shift valid element
            buff_nxt[0+:width] = buff[width*(i-1)+:width];
            en_l_var = 1'b1;
          end
          else if (din_vld_int & stat_tail)
          begin
            // update tail with input data
            buff_nxt = din;
            en_l_var = 1'b1;
          end
          else
          begin
            // no-op, disable register
            buff_nxt = din; // Don't care input to disabled flop
            en_l_var = 1'b0;
          end
          buff_pre[width*i+:width] = buff_nxt[0+:width];

          if (ph_en != 0)
            en_l[i] = en & en_l_var;
          else
            en_l[i] = en | ~en_l_var;

          if ((stat_ahead == 1'b1) & (stat[i] == 1'b0))
            //found tail, update the number of elements for count
            n_elem = ($unsigned(fifo_sz) - 1) - $unsigned(i);
        end //for loop

        // Enable for stat registers (partitioned into banks of eight)
        // Take care of the head first
        if (ph_en != 0)
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en & active;
        else
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en | ~active;

        // Now every eight
        for (i = fifo_sz-1; i >= 7; i = i - 1)
        begin
          if (($unsigned(i) % 32'd8) == 0)
          begin
            if (ph_en != 0)
              en_l_s[(i/8)-1] = en & (stat[i]) & (active);
            else
              en_l_s[(i/8)-1] = (en) | (~stat[i]) | (~active);
          end
        end

        // Update count and peak
        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = fifo_sz;
        else
          count_t = n_elem[31:0];
        count = count_t;
        // synopsys translate_off
        peak = (peak < count) ? count : peak;
        // synopsys translate_on
      end //FIFOPROC

      // Handshake valid after reset
      ccs_genreg_v1
      #(
        .width   (1),
        .ph_clk  (ph_clk),
        .ph_en   (1),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .has_en  (1'b0)
      )
      HS_INIT_REG
      (
        .clk     (clk),
        .en      (1'b1),
        .arst    (arst),
        .srst    (srst),
        .d       (1'b1),
        .z       (hs_init)
      );

      // Buffer and status registers
      for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
      begin: GEN_REGS
        ccs_genreg_v1
        #(
          .width   (1),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        STATREG
        (
          .clk     (clk),
          .en      (en_l_s[eni/8]),
          .arst    (arst),
          .srst    (srst),
          .d       (stat_pre[eni]),
          .z       (stat[eni])
        );

        ccs_genreg_v1
        #(
          .width   (width),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        BUFREG
        (
          .clk     (clk),
          .en      (en_l[eni]),
          .arst    (arst),
          .srst    (srst),
          .d       (buff_pre[width*eni+:width]),
          .z       (buff[width*eni+:width])
        );
      end

    end
    else
    begin: FEED_THRU
      assign din_rdy_drv  = dout_rdy;
      assign dout_vld_drv = din_vld;
      assign dout     = din;
      // non-blocking is not II=1 when fifo_sz=0
      assign sd = {{(sz_width-1){1'b0}}, (din_vld & ~dout_rdy)};
      assign is_idle_drv = ~(din_vld & dout_rdy);
    end
    endgenerate



endmodule

//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_pipe_v6.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
/*
 *
 *            _______________________________________________
 * WRITER    |                                              |          READER
 *           |                 ccs_pipe                     |
 *           |            ______________________            |
 *        --<| din_rdy --<|  ---------------- <|---dout_rdy<|---
 *           |            |       FIFO         |            |
 *        ---|>din_vld ---|> ----------------  |>--dout_vld |>--
 *        ---|>din -------|> ----------------  |> -----dout |>--
 *           |            |____________________|            |
 *           |______________________________________________|
 *
 *    din_rdy     - can be considered as a notFULL signal
 *    dout_vld    - can be considered as a notEMPTY signal
 *    write_stall - an internal debug signal formed from din_vld & !din_rdy
 *    read_stall  - an internal debug signal formed from dout_rdy & !dout_vld
 *    is_idle     - indicates the clock can be safely gated
 *    stall_ctrl  - Stall the pipe(fifo).  Used by STALL_FLAG_SV directive
 */

module ccs_pipe_v6 (clk, en, arst, srst, din_rdy, din_vld, din, dout_rdy, dout_vld, dout, 
                    sz, sz_req, is_idle);

    parameter integer rscid    = 0; // resource ID
    parameter integer width    = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz  = 8; // fifo depth
    parameter integer log2_sz  = 3; // log2(fifo_sz)
    parameter integer ph_clk   = 1; // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1; // clock enable polarity
    parameter integer ph_arst  = 1; // async reset polarity
    parameter integer ph_srst  = 1; // sync reset polarity

    // clock 
    input              clk;
    input              en;
    input              arst;
    input              srst;

    // writer
    output             din_rdy;
    input              din_vld;
    input  [width-1:0] din;

    // reader
    input              dout_rdy;
    output             dout_vld;
    output [width-1:0] dout;

    // size
    output [sz_width-1:0] sz;
    input                 sz_req;
    output                is_idle;

    localparam stallOff = 0; 
    wire                  stall_ctrl;
    assign stall_ctrl = stallOff;
   
    // synopsys translate_off
    wire   write_stall;
    wire   read_stall;
    assign write_stall = (din_vld & !din_rdy) | stall_ctrl;
    assign read_stall  = (dout_rdy & !dout_vld) | stall_ctrl;
    // synopsys translate_on

    wire    tmp_din_rdy;
    assign  din_rdy = tmp_din_rdy & !stall_ctrl;
    wire    tmp_dout_vld;
    assign  dout_vld = tmp_dout_vld & !stall_ctrl;
   
    ccs_fifo_wait_core_v5
    #(
        .rscid    (rscid),
        .width    (width),
        .sz_width (sz_width),
        .fifo_sz  (fifo_sz),
        .ph_clk   (ph_clk),
        .ph_en    (ph_en),
        .ph_arst  (ph_arst),
        .ph_srst  (ph_srst),
        .ph_log2  (log2_sz)
    )
    FIFO
    (
        .clk      (clk),
        .en       (en),
        .arst     (arst),
        .srst     (srst),
        .din_vld  (din_vld & !stall_ctrl),
        .din_rdy  (tmp_din_rdy),
        .din      (din),
        .dout_vld (tmp_dout_vld),
        .dout_rdy (dout_rdy & !stall_ctrl),
        .dout     (dout),
        .sd       (sz),
        .is_idle  (is_idle)
    );

endmodule


//------> ./EdgeDetect_Top.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.2/1059873 Production Release
//  HLS Date:       Mon Aug  7 10:54:31 PDT 2023
// 
//  Generated by:   b0126168@cad27
//  Generated date: Thu Sep 28 15:59:38 2023
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_7_64_7_80_80_64_5_gen
// ------------------------------------------------------------------


module EdgeDetect_VerDer_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_7_64_7_80_80_64_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [6:0] adr;
  input [6:0] adr_d;
  input [63:0] d_d;
  input en_d;
  input we_d;
  output [63:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_6_64_7_80_80_64_5_gen
// ------------------------------------------------------------------


module EdgeDetect_VerDer_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_6_64_7_80_80_64_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [6:0] adr;
  input [6:0] adr_d;
  input [63:0] d_d;
  input en_d;
  input we_d;
  output [63:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module EdgeDetect_VerDer_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output, VROW_C_0_tr0
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;
  input VROW_C_0_tr0;


  // FSM State Type Declaration for EdgeDetect_VerDer_run_run_fsm_1
  parameter
    main_C_0 = 2'd0,
    VROW_C_0 = 2'd1,
    main_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : EdgeDetect_VerDer_run_run_fsm_1
    case (state_var)
      VROW_C_0 : begin
        fsm_output = 3'b010;
        if ( VROW_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = VROW_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = VROW_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= main_C_0;
    end
    else if ( rst ) begin
      state_var <= main_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_run_staller
// ------------------------------------------------------------------


module EdgeDetect_VerDer_run_staller (
  run_wen, dat_in_rsci_wen_comp, pix_out_rsci_wen_comp, dy_rsci_wen_comp
);
  output run_wen;
  input dat_in_rsci_wen_comp;
  input pix_out_rsci_wen_comp;
  input dy_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = dat_in_rsci_wen_comp & pix_out_rsci_wen_comp & dy_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_run_wait_dp
// ------------------------------------------------------------------


module EdgeDetect_VerDer_run_wait_dp (
  line_buf0_rsci_en_d, run_wen, line_buf0_rsci_cgo, line_buf0_rsci_cgo_ir_unreg
);
  output line_buf0_rsci_en_d;
  input run_wen;
  input line_buf0_rsci_cgo;
  input line_buf0_rsci_cgo_ir_unreg;



  // Interconnect Declarations for Component Instantiations 
  assign line_buf0_rsci_en_d = run_wen & (line_buf0_rsci_cgo | line_buf0_rsci_cgo_ir_unreg);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_run_dy_rsci_dy_wait_dp
// ------------------------------------------------------------------


module EdgeDetect_VerDer_run_dy_rsci_dy_wait_dp (
  clk, rst, arst_n, dy_rsci_oswt, dy_rsci_wen_comp, dy_rsci_biwt, dy_rsci_bdwt, dy_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input dy_rsci_oswt;
  output dy_rsci_wen_comp;
  input dy_rsci_biwt;
  input dy_rsci_bdwt;
  output dy_rsci_bcwt;
  reg dy_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dy_rsci_wen_comp = (~ dy_rsci_oswt) | dy_rsci_biwt | dy_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dy_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      dy_rsci_bcwt <= 1'b0;
    end
    else begin
      dy_rsci_bcwt <= ~((~(dy_rsci_bcwt | dy_rsci_biwt)) | dy_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_run_dy_rsci_dy_wait_ctrl
// ------------------------------------------------------------------


module EdgeDetect_VerDer_run_dy_rsci_dy_wait_ctrl (
  run_wen, dy_rsci_oswt, dy_rsci_biwt, dy_rsci_bdwt, dy_rsci_bcwt, dy_rsci_irdy,
      dy_rsci_ivld_run_sct
);
  input run_wen;
  input dy_rsci_oswt;
  output dy_rsci_biwt;
  output dy_rsci_bdwt;
  input dy_rsci_bcwt;
  input dy_rsci_irdy;
  output dy_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire dy_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dy_rsci_bdwt = dy_rsci_oswt & run_wen;
  assign dy_rsci_biwt = dy_rsci_ogwt & dy_rsci_irdy;
  assign dy_rsci_ogwt = dy_rsci_oswt & (~ dy_rsci_bcwt);
  assign dy_rsci_ivld_run_sct = dy_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_run_pix_out_rsci_pix_out_wait_dp
// ------------------------------------------------------------------


module EdgeDetect_VerDer_run_pix_out_rsci_pix_out_wait_dp (
  clk, rst, arst_n, pix_out_rsci_oswt, pix_out_rsci_wen_comp, pix_out_rsci_biwt,
      pix_out_rsci_bdwt, pix_out_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input pix_out_rsci_oswt;
  output pix_out_rsci_wen_comp;
  input pix_out_rsci_biwt;
  input pix_out_rsci_bdwt;
  output pix_out_rsci_bcwt;
  reg pix_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign pix_out_rsci_wen_comp = (~ pix_out_rsci_oswt) | pix_out_rsci_biwt | pix_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      pix_out_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      pix_out_rsci_bcwt <= 1'b0;
    end
    else begin
      pix_out_rsci_bcwt <= ~((~(pix_out_rsci_bcwt | pix_out_rsci_biwt)) | pix_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_run_pix_out_rsci_pix_out_wait_ctrl
// ------------------------------------------------------------------


module EdgeDetect_VerDer_run_pix_out_rsci_pix_out_wait_ctrl (
  run_wen, pix_out_rsci_oswt, pix_out_rsci_biwt, pix_out_rsci_bdwt, pix_out_rsci_bcwt,
      pix_out_rsci_irdy, pix_out_rsci_ivld_run_sct
);
  input run_wen;
  input pix_out_rsci_oswt;
  output pix_out_rsci_biwt;
  output pix_out_rsci_bdwt;
  input pix_out_rsci_bcwt;
  input pix_out_rsci_irdy;
  output pix_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire pix_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign pix_out_rsci_bdwt = pix_out_rsci_oswt & run_wen;
  assign pix_out_rsci_biwt = pix_out_rsci_ogwt & pix_out_rsci_irdy;
  assign pix_out_rsci_ogwt = pix_out_rsci_oswt & (~ pix_out_rsci_bcwt);
  assign pix_out_rsci_ivld_run_sct = pix_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_run_dat_in_rsci_dat_in_wait_dp
// ------------------------------------------------------------------


module EdgeDetect_VerDer_run_dat_in_rsci_dat_in_wait_dp (
  clk, rst, arst_n, dat_in_rsci_oswt, dat_in_rsci_wen_comp, dat_in_rsci_idat_mxwt,
      dat_in_rsci_biwt, dat_in_rsci_bdwt, dat_in_rsci_bcwt, dat_in_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  input dat_in_rsci_oswt;
  output dat_in_rsci_wen_comp;
  output [31:0] dat_in_rsci_idat_mxwt;
  input dat_in_rsci_biwt;
  input dat_in_rsci_bdwt;
  output dat_in_rsci_bcwt;
  reg dat_in_rsci_bcwt;
  input [33:0] dat_in_rsci_idat;


  // Interconnect Declarations
  reg [31:0] dat_in_rsci_idat_bfwt_31_0;


  // Interconnect Declarations for Component Instantiations 
  assign dat_in_rsci_wen_comp = (~ dat_in_rsci_oswt) | dat_in_rsci_biwt | dat_in_rsci_bcwt;
  assign dat_in_rsci_idat_mxwt = MUX_v_32_2_2((dat_in_rsci_idat[31:0]), dat_in_rsci_idat_bfwt_31_0,
      dat_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dat_in_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      dat_in_rsci_bcwt <= 1'b0;
    end
    else begin
      dat_in_rsci_bcwt <= ~((~(dat_in_rsci_bcwt | dat_in_rsci_biwt)) | dat_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dat_in_rsci_idat_bfwt_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      dat_in_rsci_idat_bfwt_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( dat_in_rsci_biwt ) begin
      dat_in_rsci_idat_bfwt_31_0 <= dat_in_rsci_idat[31:0];
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_run_dat_in_rsci_dat_in_wait_ctrl
// ------------------------------------------------------------------


module EdgeDetect_VerDer_run_dat_in_rsci_dat_in_wait_ctrl (
  run_wen, dat_in_rsci_oswt, dat_in_rsci_biwt, dat_in_rsci_bdwt, dat_in_rsci_bcwt,
      dat_in_rsci_irdy_run_sct, dat_in_rsci_ivld
);
  input run_wen;
  input dat_in_rsci_oswt;
  output dat_in_rsci_biwt;
  output dat_in_rsci_bdwt;
  input dat_in_rsci_bcwt;
  output dat_in_rsci_irdy_run_sct;
  input dat_in_rsci_ivld;


  // Interconnect Declarations
  wire dat_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dat_in_rsci_bdwt = dat_in_rsci_oswt & run_wen;
  assign dat_in_rsci_biwt = dat_in_rsci_ogwt & dat_in_rsci_ivld;
  assign dat_in_rsci_ogwt = dat_in_rsci_oswt & (~ dat_in_rsci_bcwt);
  assign dat_in_rsci_irdy_run_sct = dat_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_HorDer_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module EdgeDetect_HorDer_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output, HROW_C_0_tr0
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;
  input HROW_C_0_tr0;


  // FSM State Type Declaration for EdgeDetect_HorDer_run_run_fsm_1
  parameter
    main_C_0 = 2'd0,
    HROW_C_0 = 2'd1,
    main_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : EdgeDetect_HorDer_run_run_fsm_1
    case (state_var)
      HROW_C_0 : begin
        fsm_output = 3'b010;
        if ( HROW_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = HROW_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = HROW_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= main_C_0;
    end
    else if ( rst ) begin
      state_var <= main_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_HorDer_run_staller
// ------------------------------------------------------------------


module EdgeDetect_HorDer_run_staller (
  run_wen, pix_in_rsci_wen_comp, pix_out_rsci_wen_comp, dx_rsci_wen_comp
);
  output run_wen;
  input pix_in_rsci_wen_comp;
  input pix_out_rsci_wen_comp;
  input dx_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = pix_in_rsci_wen_comp & pix_out_rsci_wen_comp & dx_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_HorDer_run_dx_rsci_dx_wait_dp
// ------------------------------------------------------------------


module EdgeDetect_HorDer_run_dx_rsci_dx_wait_dp (
  clk, rst, arst_n, dx_rsci_oswt, dx_rsci_wen_comp, dx_rsci_biwt, dx_rsci_bdwt, dx_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input dx_rsci_oswt;
  output dx_rsci_wen_comp;
  input dx_rsci_biwt;
  input dx_rsci_bdwt;
  output dx_rsci_bcwt;
  reg dx_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dx_rsci_wen_comp = (~ dx_rsci_oswt) | dx_rsci_biwt | dx_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dx_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      dx_rsci_bcwt <= 1'b0;
    end
    else begin
      dx_rsci_bcwt <= ~((~(dx_rsci_bcwt | dx_rsci_biwt)) | dx_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_HorDer_run_dx_rsci_dx_wait_ctrl
// ------------------------------------------------------------------


module EdgeDetect_HorDer_run_dx_rsci_dx_wait_ctrl (
  run_wen, dx_rsci_oswt, dx_rsci_biwt, dx_rsci_bdwt, dx_rsci_bcwt, dx_rsci_irdy,
      dx_rsci_ivld_run_sct
);
  input run_wen;
  input dx_rsci_oswt;
  output dx_rsci_biwt;
  output dx_rsci_bdwt;
  input dx_rsci_bcwt;
  input dx_rsci_irdy;
  output dx_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire dx_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dx_rsci_bdwt = dx_rsci_oswt & run_wen;
  assign dx_rsci_biwt = dx_rsci_ogwt & dx_rsci_irdy;
  assign dx_rsci_ogwt = dx_rsci_oswt & (~ dx_rsci_bcwt);
  assign dx_rsci_ivld_run_sct = dx_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_HorDer_run_pix_out_rsci_pix_out_wait_dp
// ------------------------------------------------------------------


module EdgeDetect_HorDer_run_pix_out_rsci_pix_out_wait_dp (
  clk, rst, arst_n, pix_out_rsci_oswt, pix_out_rsci_wen_comp, pix_out_rsci_biwt,
      pix_out_rsci_bdwt, pix_out_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input pix_out_rsci_oswt;
  output pix_out_rsci_wen_comp;
  input pix_out_rsci_biwt;
  input pix_out_rsci_bdwt;
  output pix_out_rsci_bcwt;
  reg pix_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign pix_out_rsci_wen_comp = (~ pix_out_rsci_oswt) | pix_out_rsci_biwt | pix_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      pix_out_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      pix_out_rsci_bcwt <= 1'b0;
    end
    else begin
      pix_out_rsci_bcwt <= ~((~(pix_out_rsci_bcwt | pix_out_rsci_biwt)) | pix_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_HorDer_run_pix_out_rsci_pix_out_wait_ctrl
// ------------------------------------------------------------------


module EdgeDetect_HorDer_run_pix_out_rsci_pix_out_wait_ctrl (
  run_wen, pix_out_rsci_oswt, pix_out_rsci_biwt, pix_out_rsci_bdwt, pix_out_rsci_bcwt,
      pix_out_rsci_irdy, pix_out_rsci_ivld_run_sct
);
  input run_wen;
  input pix_out_rsci_oswt;
  output pix_out_rsci_biwt;
  output pix_out_rsci_bdwt;
  input pix_out_rsci_bcwt;
  input pix_out_rsci_irdy;
  output pix_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire pix_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign pix_out_rsci_bdwt = pix_out_rsci_oswt & run_wen;
  assign pix_out_rsci_biwt = pix_out_rsci_ogwt & pix_out_rsci_irdy;
  assign pix_out_rsci_ogwt = pix_out_rsci_oswt & (~ pix_out_rsci_bcwt);
  assign pix_out_rsci_ivld_run_sct = pix_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_HorDer_run_pix_in_rsci_pix_in_wait_ctrl
// ------------------------------------------------------------------


module EdgeDetect_HorDer_run_pix_in_rsci_pix_in_wait_ctrl (
  run_wen, pix_in_rsci_iswt0, pix_in_rsci_irdy_run_sct
);
  input run_wen;
  input pix_in_rsci_iswt0;
  output pix_in_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign pix_in_rsci_irdy_run_sct = pix_in_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output, MROW_C_0_tr0
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;
  input MROW_C_0_tr0;


  // FSM State Type Declaration for EdgeDetect_MagAng_run_run_fsm_1
  parameter
    main_C_0 = 2'd0,
    MROW_C_0 = 2'd1,
    main_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : EdgeDetect_MagAng_run_run_fsm_1
    case (state_var)
      MROW_C_0 : begin
        fsm_output = 3'b010;
        if ( MROW_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = MROW_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = MROW_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= main_C_0;
    end
    else if ( rst ) begin
      state_var <= main_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_staller
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_staller (
  clk, rst, arst_n, run_wen, run_wten, dx_in_rsci_wen_comp, dy_in_rsci_wen_comp,
      pix_in_rsci_wen_comp, dat_out_rsci_wen_comp
);
  input clk;
  input rst;
  input arst_n;
  output run_wen;
  output run_wten;
  reg run_wten;
  input dx_in_rsci_wen_comp;
  input dy_in_rsci_wen_comp;
  input pix_in_rsci_wen_comp;
  input dat_out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = dx_in_rsci_wen_comp & dy_in_rsci_wen_comp & pix_in_rsci_wen_comp
      & dat_out_rsci_wen_comp;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten <= 1'b0;
    end
    else if ( rst ) begin
      run_wten <= 1'b0;
    end
    else begin
      run_wten <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_crc32_dat_out_triosy_obj_crc32_dat_out_triosy_wait_ctrl
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_crc32_dat_out_triosy_obj_crc32_dat_out_triosy_wait_ctrl
    (
  run_wten, crc32_dat_out_triosy_obj_iswt0, crc32_dat_out_triosy_obj_biwt
);
  input run_wten;
  input crc32_dat_out_triosy_obj_iswt0;
  output crc32_dat_out_triosy_obj_biwt;



  // Interconnect Declarations for Component Instantiations 
  assign crc32_dat_out_triosy_obj_biwt = (~ run_wten) & crc32_dat_out_triosy_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_crc32_pix_in_triosy_obj_crc32_pix_in_triosy_wait_ctrl
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_crc32_pix_in_triosy_obj_crc32_pix_in_triosy_wait_ctrl
    (
  run_wten, crc32_pix_in_triosy_obj_iswt0, crc32_pix_in_triosy_obj_biwt
);
  input run_wten;
  input crc32_pix_in_triosy_obj_iswt0;
  output crc32_pix_in_triosy_obj_biwt;



  // Interconnect Declarations for Component Instantiations 
  assign crc32_pix_in_triosy_obj_biwt = (~ run_wten) & crc32_pix_in_triosy_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_dat_out_rsci_dat_out_wait_dp
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_dat_out_rsci_dat_out_wait_dp (
  clk, rst, arst_n, dat_out_rsci_oswt, dat_out_rsci_wen_comp, dat_out_rsci_biwt,
      dat_out_rsci_bdwt, dat_out_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input dat_out_rsci_oswt;
  output dat_out_rsci_wen_comp;
  input dat_out_rsci_biwt;
  input dat_out_rsci_bdwt;
  output dat_out_rsci_bcwt;
  reg dat_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dat_out_rsci_wen_comp = (~ dat_out_rsci_oswt) | dat_out_rsci_biwt | dat_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dat_out_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      dat_out_rsci_bcwt <= 1'b0;
    end
    else begin
      dat_out_rsci_bcwt <= ~((~(dat_out_rsci_bcwt | dat_out_rsci_biwt)) | dat_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_dat_out_rsci_dat_out_wait_ctrl
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_dat_out_rsci_dat_out_wait_ctrl (
  run_wen, dat_out_rsci_oswt, dat_out_rsci_biwt, dat_out_rsci_bdwt, dat_out_rsci_bcwt,
      dat_out_rsci_irdy, dat_out_rsci_ivld_run_sct
);
  input run_wen;
  input dat_out_rsci_oswt;
  output dat_out_rsci_biwt;
  output dat_out_rsci_bdwt;
  input dat_out_rsci_bcwt;
  input dat_out_rsci_irdy;
  output dat_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire dat_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dat_out_rsci_bdwt = dat_out_rsci_oswt & run_wen;
  assign dat_out_rsci_biwt = dat_out_rsci_ogwt & dat_out_rsci_irdy;
  assign dat_out_rsci_ogwt = dat_out_rsci_oswt & (~ dat_out_rsci_bcwt);
  assign dat_out_rsci_ivld_run_sct = dat_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_pix_in_rsci_pix_in_wait_dp
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_pix_in_rsci_pix_in_wait_dp (
  clk, rst, arst_n, pix_in_rsci_oswt, pix_in_rsci_wen_comp, pix_in_rsci_idat_mxwt,
      pix_in_rsci_biwt, pix_in_rsci_bdwt, pix_in_rsci_bcwt, pix_in_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  input pix_in_rsci_oswt;
  output pix_in_rsci_wen_comp;
  output [31:0] pix_in_rsci_idat_mxwt;
  input pix_in_rsci_biwt;
  input pix_in_rsci_bdwt;
  output pix_in_rsci_bcwt;
  reg pix_in_rsci_bcwt;
  input [31:0] pix_in_rsci_idat;


  // Interconnect Declarations
  reg [31:0] pix_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign pix_in_rsci_wen_comp = (~ pix_in_rsci_oswt) | pix_in_rsci_biwt | pix_in_rsci_bcwt;
  assign pix_in_rsci_idat_mxwt = MUX_v_32_2_2(pix_in_rsci_idat, pix_in_rsci_idat_bfwt,
      pix_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      pix_in_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      pix_in_rsci_bcwt <= 1'b0;
    end
    else begin
      pix_in_rsci_bcwt <= ~((~(pix_in_rsci_bcwt | pix_in_rsci_biwt)) | pix_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      pix_in_rsci_idat_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      pix_in_rsci_idat_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( pix_in_rsci_biwt ) begin
      pix_in_rsci_idat_bfwt <= pix_in_rsci_idat;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_pix_in_rsci_pix_in_wait_ctrl
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_pix_in_rsci_pix_in_wait_ctrl (
  run_wen, pix_in_rsci_oswt, pix_in_rsci_biwt, pix_in_rsci_bdwt, pix_in_rsci_bcwt,
      pix_in_rsci_irdy_run_sct, pix_in_rsci_ivld
);
  input run_wen;
  input pix_in_rsci_oswt;
  output pix_in_rsci_biwt;
  output pix_in_rsci_bdwt;
  input pix_in_rsci_bcwt;
  output pix_in_rsci_irdy_run_sct;
  input pix_in_rsci_ivld;


  // Interconnect Declarations
  wire pix_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign pix_in_rsci_bdwt = pix_in_rsci_oswt & run_wen;
  assign pix_in_rsci_biwt = pix_in_rsci_ogwt & pix_in_rsci_ivld;
  assign pix_in_rsci_ogwt = pix_in_rsci_oswt & (~ pix_in_rsci_bcwt);
  assign pix_in_rsci_irdy_run_sct = pix_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_dy_in_rsci_dy_in_wait_ctrl
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_dy_in_rsci_dy_in_wait_ctrl (
  run_wen, dy_in_rsci_iswt0, dy_in_rsci_irdy_run_sct
);
  input run_wen;
  input dy_in_rsci_iswt0;
  output dy_in_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dy_in_rsci_irdy_run_sct = dy_in_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_dx_in_rsci_dx_in_wait_ctrl
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_dx_in_rsci_dx_in_wait_ctrl (
  run_wen, dx_in_rsci_iswt0, dx_in_rsci_irdy_run_sct
);
  input run_wen;
  input dx_in_rsci_iswt0;
  output dx_in_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dx_in_rsci_irdy_run_sct = dx_in_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_run_dy_rsci
// ------------------------------------------------------------------


module EdgeDetect_VerDer_run_dy_rsci (
  clk, rst, arst_n, dy_rsc_dat, dy_rsc_vld, dy_rsc_rdy, run_wen, dy_rsci_oswt, dy_rsci_wen_comp,
      dy_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [35:0] dy_rsc_dat;
  output dy_rsc_vld;
  input dy_rsc_rdy;
  input run_wen;
  input dy_rsci_oswt;
  output dy_rsci_wen_comp;
  input [35:0] dy_rsci_idat;


  // Interconnect Declarations
  wire dy_rsci_biwt;
  wire dy_rsci_bdwt;
  wire dy_rsci_bcwt;
  wire dy_rsci_irdy;
  wire dy_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd5),
  .width(32'sd36)) dy_rsci (
      .irdy(dy_rsci_irdy),
      .ivld(dy_rsci_ivld_run_sct),
      .idat(dy_rsci_idat),
      .rdy(dy_rsc_rdy),
      .vld(dy_rsc_vld),
      .dat(dy_rsc_dat)
    );
  EdgeDetect_VerDer_run_dy_rsci_dy_wait_ctrl EdgeDetect_VerDer_run_dy_rsci_dy_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dy_rsci_oswt(dy_rsci_oswt),
      .dy_rsci_biwt(dy_rsci_biwt),
      .dy_rsci_bdwt(dy_rsci_bdwt),
      .dy_rsci_bcwt(dy_rsci_bcwt),
      .dy_rsci_irdy(dy_rsci_irdy),
      .dy_rsci_ivld_run_sct(dy_rsci_ivld_run_sct)
    );
  EdgeDetect_VerDer_run_dy_rsci_dy_wait_dp EdgeDetect_VerDer_run_dy_rsci_dy_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .dy_rsci_oswt(dy_rsci_oswt),
      .dy_rsci_wen_comp(dy_rsci_wen_comp),
      .dy_rsci_biwt(dy_rsci_biwt),
      .dy_rsci_bdwt(dy_rsci_bdwt),
      .dy_rsci_bcwt(dy_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_run_pix_out_rsci
// ------------------------------------------------------------------


module EdgeDetect_VerDer_run_pix_out_rsci (
  clk, rst, arst_n, pix_out_rsc_dat, pix_out_rsc_vld, pix_out_rsc_rdy, run_wen, pix_out_rsci_oswt,
      pix_out_rsci_wen_comp, pix_out_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [31:0] pix_out_rsc_dat;
  output pix_out_rsc_vld;
  input pix_out_rsc_rdy;
  input run_wen;
  input pix_out_rsci_oswt;
  output pix_out_rsci_wen_comp;
  input [31:0] pix_out_rsci_idat;


  // Interconnect Declarations
  wire pix_out_rsci_biwt;
  wire pix_out_rsci_bdwt;
  wire pix_out_rsci_bcwt;
  wire pix_out_rsci_irdy;
  wire pix_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd4),
  .width(32'sd32)) pix_out_rsci (
      .irdy(pix_out_rsci_irdy),
      .ivld(pix_out_rsci_ivld_run_sct),
      .idat(pix_out_rsci_idat),
      .rdy(pix_out_rsc_rdy),
      .vld(pix_out_rsc_vld),
      .dat(pix_out_rsc_dat)
    );
  EdgeDetect_VerDer_run_pix_out_rsci_pix_out_wait_ctrl EdgeDetect_VerDer_run_pix_out_rsci_pix_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .pix_out_rsci_oswt(pix_out_rsci_oswt),
      .pix_out_rsci_biwt(pix_out_rsci_biwt),
      .pix_out_rsci_bdwt(pix_out_rsci_bdwt),
      .pix_out_rsci_bcwt(pix_out_rsci_bcwt),
      .pix_out_rsci_irdy(pix_out_rsci_irdy),
      .pix_out_rsci_ivld_run_sct(pix_out_rsci_ivld_run_sct)
    );
  EdgeDetect_VerDer_run_pix_out_rsci_pix_out_wait_dp EdgeDetect_VerDer_run_pix_out_rsci_pix_out_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .pix_out_rsci_oswt(pix_out_rsci_oswt),
      .pix_out_rsci_wen_comp(pix_out_rsci_wen_comp),
      .pix_out_rsci_biwt(pix_out_rsci_biwt),
      .pix_out_rsci_bdwt(pix_out_rsci_bdwt),
      .pix_out_rsci_bcwt(pix_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_run_dat_in_rsci
// ------------------------------------------------------------------


module EdgeDetect_VerDer_run_dat_in_rsci (
  clk, rst, arst_n, dat_in_rsc_dat, dat_in_rsc_vld, dat_in_rsc_rdy, run_wen, dat_in_rsci_oswt,
      dat_in_rsci_wen_comp, dat_in_rsci_idat_mxwt
);
  input clk;
  input rst;
  input arst_n;
  input [33:0] dat_in_rsc_dat;
  input dat_in_rsc_vld;
  output dat_in_rsc_rdy;
  input run_wen;
  input dat_in_rsci_oswt;
  output dat_in_rsci_wen_comp;
  output [31:0] dat_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire dat_in_rsci_biwt;
  wire dat_in_rsci_bdwt;
  wire dat_in_rsci_bcwt;
  wire dat_in_rsci_irdy_run_sct;
  wire dat_in_rsci_ivld;
  wire [33:0] dat_in_rsci_idat;
  wire [31:0] dat_in_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd34)) dat_in_rsci (
      .rdy(dat_in_rsc_rdy),
      .vld(dat_in_rsc_vld),
      .dat(dat_in_rsc_dat),
      .irdy(dat_in_rsci_irdy_run_sct),
      .ivld(dat_in_rsci_ivld),
      .idat(dat_in_rsci_idat)
    );
  EdgeDetect_VerDer_run_dat_in_rsci_dat_in_wait_ctrl EdgeDetect_VerDer_run_dat_in_rsci_dat_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dat_in_rsci_oswt(dat_in_rsci_oswt),
      .dat_in_rsci_biwt(dat_in_rsci_biwt),
      .dat_in_rsci_bdwt(dat_in_rsci_bdwt),
      .dat_in_rsci_bcwt(dat_in_rsci_bcwt),
      .dat_in_rsci_irdy_run_sct(dat_in_rsci_irdy_run_sct),
      .dat_in_rsci_ivld(dat_in_rsci_ivld)
    );
  EdgeDetect_VerDer_run_dat_in_rsci_dat_in_wait_dp EdgeDetect_VerDer_run_dat_in_rsci_dat_in_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .dat_in_rsci_oswt(dat_in_rsci_oswt),
      .dat_in_rsci_wen_comp(dat_in_rsci_wen_comp),
      .dat_in_rsci_idat_mxwt(dat_in_rsci_idat_mxwt_pconst),
      .dat_in_rsci_biwt(dat_in_rsci_biwt),
      .dat_in_rsci_bdwt(dat_in_rsci_bdwt),
      .dat_in_rsci_bcwt(dat_in_rsci_bcwt),
      .dat_in_rsci_idat(dat_in_rsci_idat)
    );
  assign dat_in_rsci_idat_mxwt = dat_in_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_HorDer_run_dx_rsci
// ------------------------------------------------------------------


module EdgeDetect_HorDer_run_dx_rsci (
  clk, rst, arst_n, dx_rsc_dat, dx_rsc_vld, dx_rsc_rdy, run_wen, dx_rsci_oswt, dx_rsci_wen_comp,
      dx_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [35:0] dx_rsc_dat;
  output dx_rsc_vld;
  input dx_rsc_rdy;
  input run_wen;
  input dx_rsci_oswt;
  output dx_rsci_wen_comp;
  input [35:0] dx_rsci_idat;


  // Interconnect Declarations
  wire dx_rsci_biwt;
  wire dx_rsci_bdwt;
  wire dx_rsci_bcwt;
  wire dx_rsci_irdy;
  wire dx_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd12),
  .width(32'sd36)) dx_rsci (
      .irdy(dx_rsci_irdy),
      .ivld(dx_rsci_ivld_run_sct),
      .idat(dx_rsci_idat),
      .rdy(dx_rsc_rdy),
      .vld(dx_rsc_vld),
      .dat(dx_rsc_dat)
    );
  EdgeDetect_HorDer_run_dx_rsci_dx_wait_ctrl EdgeDetect_HorDer_run_dx_rsci_dx_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dx_rsci_oswt(dx_rsci_oswt),
      .dx_rsci_biwt(dx_rsci_biwt),
      .dx_rsci_bdwt(dx_rsci_bdwt),
      .dx_rsci_bcwt(dx_rsci_bcwt),
      .dx_rsci_irdy(dx_rsci_irdy),
      .dx_rsci_ivld_run_sct(dx_rsci_ivld_run_sct)
    );
  EdgeDetect_HorDer_run_dx_rsci_dx_wait_dp EdgeDetect_HorDer_run_dx_rsci_dx_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .dx_rsci_oswt(dx_rsci_oswt),
      .dx_rsci_wen_comp(dx_rsci_wen_comp),
      .dx_rsci_biwt(dx_rsci_biwt),
      .dx_rsci_bdwt(dx_rsci_bdwt),
      .dx_rsci_bcwt(dx_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_HorDer_run_pix_out_rsci
// ------------------------------------------------------------------


module EdgeDetect_HorDer_run_pix_out_rsci (
  clk, rst, arst_n, pix_out_rsc_dat, pix_out_rsc_vld, pix_out_rsc_rdy, run_wen, pix_out_rsci_oswt,
      pix_out_rsci_wen_comp, pix_out_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [31:0] pix_out_rsc_dat;
  output pix_out_rsc_vld;
  input pix_out_rsc_rdy;
  input run_wen;
  input pix_out_rsci_oswt;
  output pix_out_rsci_wen_comp;
  input [31:0] pix_out_rsci_idat;


  // Interconnect Declarations
  wire pix_out_rsci_biwt;
  wire pix_out_rsci_bdwt;
  wire pix_out_rsci_bcwt;
  wire pix_out_rsci_irdy;
  wire pix_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd11),
  .width(32'sd32)) pix_out_rsci (
      .irdy(pix_out_rsci_irdy),
      .ivld(pix_out_rsci_ivld_run_sct),
      .idat(pix_out_rsci_idat),
      .rdy(pix_out_rsc_rdy),
      .vld(pix_out_rsc_vld),
      .dat(pix_out_rsc_dat)
    );
  EdgeDetect_HorDer_run_pix_out_rsci_pix_out_wait_ctrl EdgeDetect_HorDer_run_pix_out_rsci_pix_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .pix_out_rsci_oswt(pix_out_rsci_oswt),
      .pix_out_rsci_biwt(pix_out_rsci_biwt),
      .pix_out_rsci_bdwt(pix_out_rsci_bdwt),
      .pix_out_rsci_bcwt(pix_out_rsci_bcwt),
      .pix_out_rsci_irdy(pix_out_rsci_irdy),
      .pix_out_rsci_ivld_run_sct(pix_out_rsci_ivld_run_sct)
    );
  EdgeDetect_HorDer_run_pix_out_rsci_pix_out_wait_dp EdgeDetect_HorDer_run_pix_out_rsci_pix_out_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .pix_out_rsci_oswt(pix_out_rsci_oswt),
      .pix_out_rsci_wen_comp(pix_out_rsci_wen_comp),
      .pix_out_rsci_biwt(pix_out_rsci_biwt),
      .pix_out_rsci_bdwt(pix_out_rsci_bdwt),
      .pix_out_rsci_bcwt(pix_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_HorDer_run_pix_in_rsci
// ------------------------------------------------------------------


module EdgeDetect_HorDer_run_pix_in_rsci (
  pix_in_rsc_dat, pix_in_rsc_vld, pix_in_rsc_rdy, run_wen, pix_in_rsci_oswt, pix_in_rsci_wen_comp,
      pix_in_rsci_idat_mxwt
);
  input [31:0] pix_in_rsc_dat;
  input pix_in_rsc_vld;
  output pix_in_rsc_rdy;
  input run_wen;
  input pix_in_rsci_oswt;
  output pix_in_rsci_wen_comp;
  output [31:0] pix_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire pix_in_rsci_irdy_run_sct;
  wire pix_in_rsci_ivld;
  wire [31:0] pix_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd8),
  .width(32'sd32)) pix_in_rsci (
      .rdy(pix_in_rsc_rdy),
      .vld(pix_in_rsc_vld),
      .dat(pix_in_rsc_dat),
      .irdy(pix_in_rsci_irdy_run_sct),
      .ivld(pix_in_rsci_ivld),
      .idat(pix_in_rsci_idat)
    );
  EdgeDetect_HorDer_run_pix_in_rsci_pix_in_wait_ctrl EdgeDetect_HorDer_run_pix_in_rsci_pix_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .pix_in_rsci_iswt0(pix_in_rsci_oswt),
      .pix_in_rsci_irdy_run_sct(pix_in_rsci_irdy_run_sct)
    );
  assign pix_in_rsci_idat_mxwt = pix_in_rsci_idat;
  assign pix_in_rsci_wen_comp = (~ pix_in_rsci_oswt) | pix_in_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_crc32_dat_out_triosy_obj
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_crc32_dat_out_triosy_obj (
  crc32_dat_out_triosy_lz, run_wten, crc32_dat_out_triosy_obj_iswt0
);
  output crc32_dat_out_triosy_lz;
  input run_wten;
  input crc32_dat_out_triosy_obj_iswt0;


  // Interconnect Declarations
  wire crc32_dat_out_triosy_obj_biwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) crc32_dat_out_triosy_obj (
      .ld(crc32_dat_out_triosy_obj_biwt),
      .lz(crc32_dat_out_triosy_lz)
    );
  EdgeDetect_MagAng_run_crc32_dat_out_triosy_obj_crc32_dat_out_triosy_wait_ctrl EdgeDetect_MagAng_run_crc32_dat_out_triosy_obj_crc32_dat_out_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .crc32_dat_out_triosy_obj_iswt0(crc32_dat_out_triosy_obj_iswt0),
      .crc32_dat_out_triosy_obj_biwt(crc32_dat_out_triosy_obj_biwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_crc32_pix_in_triosy_obj
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_crc32_pix_in_triosy_obj (
  crc32_pix_in_triosy_lz, run_wten, crc32_pix_in_triosy_obj_iswt0
);
  output crc32_pix_in_triosy_lz;
  input run_wten;
  input crc32_pix_in_triosy_obj_iswt0;


  // Interconnect Declarations
  wire crc32_pix_in_triosy_obj_biwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) crc32_pix_in_triosy_obj (
      .ld(crc32_pix_in_triosy_obj_biwt),
      .lz(crc32_pix_in_triosy_lz)
    );
  EdgeDetect_MagAng_run_crc32_pix_in_triosy_obj_crc32_pix_in_triosy_wait_ctrl EdgeDetect_MagAng_run_crc32_pix_in_triosy_obj_crc32_pix_in_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .crc32_pix_in_triosy_obj_iswt0(crc32_pix_in_triosy_obj_iswt0),
      .crc32_pix_in_triosy_obj_biwt(crc32_pix_in_triosy_obj_biwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_dat_out_rsci
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_dat_out_rsci (
  clk, rst, arst_n, dat_out_rsc_dat, dat_out_rsc_vld, dat_out_rsc_rdy, run_wen, dat_out_rsci_oswt,
      dat_out_rsci_wen_comp, dat_out_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [33:0] dat_out_rsc_dat;
  output dat_out_rsc_vld;
  input dat_out_rsc_rdy;
  input run_wen;
  input dat_out_rsci_oswt;
  output dat_out_rsci_wen_comp;
  input [33:0] dat_out_rsci_idat;


  // Interconnect Declarations
  wire dat_out_rsci_biwt;
  wire dat_out_rsci_bdwt;
  wire dat_out_rsci_bcwt;
  wire dat_out_rsci_irdy;
  wire dat_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd22),
  .width(32'sd34)) dat_out_rsci (
      .irdy(dat_out_rsci_irdy),
      .ivld(dat_out_rsci_ivld_run_sct),
      .idat(dat_out_rsci_idat),
      .rdy(dat_out_rsc_rdy),
      .vld(dat_out_rsc_vld),
      .dat(dat_out_rsc_dat)
    );
  EdgeDetect_MagAng_run_dat_out_rsci_dat_out_wait_ctrl EdgeDetect_MagAng_run_dat_out_rsci_dat_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dat_out_rsci_oswt(dat_out_rsci_oswt),
      .dat_out_rsci_biwt(dat_out_rsci_biwt),
      .dat_out_rsci_bdwt(dat_out_rsci_bdwt),
      .dat_out_rsci_bcwt(dat_out_rsci_bcwt),
      .dat_out_rsci_irdy(dat_out_rsci_irdy),
      .dat_out_rsci_ivld_run_sct(dat_out_rsci_ivld_run_sct)
    );
  EdgeDetect_MagAng_run_dat_out_rsci_dat_out_wait_dp EdgeDetect_MagAng_run_dat_out_rsci_dat_out_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .dat_out_rsci_oswt(dat_out_rsci_oswt),
      .dat_out_rsci_wen_comp(dat_out_rsci_wen_comp),
      .dat_out_rsci_biwt(dat_out_rsci_biwt),
      .dat_out_rsci_bdwt(dat_out_rsci_bdwt),
      .dat_out_rsci_bcwt(dat_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_pix_in_rsci
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_pix_in_rsci (
  clk, rst, arst_n, pix_in_rsc_dat, pix_in_rsc_vld, pix_in_rsc_rdy, run_wen, pix_in_rsci_oswt,
      pix_in_rsci_wen_comp, pix_in_rsci_idat_mxwt
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] pix_in_rsc_dat;
  input pix_in_rsc_vld;
  output pix_in_rsc_rdy;
  input run_wen;
  input pix_in_rsci_oswt;
  output pix_in_rsci_wen_comp;
  output [31:0] pix_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire pix_in_rsci_biwt;
  wire pix_in_rsci_bdwt;
  wire pix_in_rsci_bcwt;
  wire pix_in_rsci_irdy_run_sct;
  wire pix_in_rsci_ivld;
  wire [31:0] pix_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd16),
  .width(32'sd32)) pix_in_rsci (
      .rdy(pix_in_rsc_rdy),
      .vld(pix_in_rsc_vld),
      .dat(pix_in_rsc_dat),
      .irdy(pix_in_rsci_irdy_run_sct),
      .ivld(pix_in_rsci_ivld),
      .idat(pix_in_rsci_idat)
    );
  EdgeDetect_MagAng_run_pix_in_rsci_pix_in_wait_ctrl EdgeDetect_MagAng_run_pix_in_rsci_pix_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .pix_in_rsci_oswt(pix_in_rsci_oswt),
      .pix_in_rsci_biwt(pix_in_rsci_biwt),
      .pix_in_rsci_bdwt(pix_in_rsci_bdwt),
      .pix_in_rsci_bcwt(pix_in_rsci_bcwt),
      .pix_in_rsci_irdy_run_sct(pix_in_rsci_irdy_run_sct),
      .pix_in_rsci_ivld(pix_in_rsci_ivld)
    );
  EdgeDetect_MagAng_run_pix_in_rsci_pix_in_wait_dp EdgeDetect_MagAng_run_pix_in_rsci_pix_in_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .pix_in_rsci_oswt(pix_in_rsci_oswt),
      .pix_in_rsci_wen_comp(pix_in_rsci_wen_comp),
      .pix_in_rsci_idat_mxwt(pix_in_rsci_idat_mxwt),
      .pix_in_rsci_biwt(pix_in_rsci_biwt),
      .pix_in_rsci_bdwt(pix_in_rsci_bdwt),
      .pix_in_rsci_bcwt(pix_in_rsci_bcwt),
      .pix_in_rsci_idat(pix_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_dy_in_rsci
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_dy_in_rsci (
  dy_in_rsc_dat, dy_in_rsc_vld, dy_in_rsc_rdy, run_wen, dy_in_rsci_oswt, dy_in_rsci_wen_comp,
      dy_in_rsci_idat_mxwt
);
  input [35:0] dy_in_rsc_dat;
  input dy_in_rsc_vld;
  output dy_in_rsc_rdy;
  input run_wen;
  input dy_in_rsci_oswt;
  output dy_in_rsci_wen_comp;
  output [35:0] dy_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire dy_in_rsci_irdy_run_sct;
  wire dy_in_rsci_ivld;
  wire [35:0] dy_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd15),
  .width(32'sd36)) dy_in_rsci (
      .rdy(dy_in_rsc_rdy),
      .vld(dy_in_rsc_vld),
      .dat(dy_in_rsc_dat),
      .irdy(dy_in_rsci_irdy_run_sct),
      .ivld(dy_in_rsci_ivld),
      .idat(dy_in_rsci_idat)
    );
  EdgeDetect_MagAng_run_dy_in_rsci_dy_in_wait_ctrl EdgeDetect_MagAng_run_dy_in_rsci_dy_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dy_in_rsci_iswt0(dy_in_rsci_oswt),
      .dy_in_rsci_irdy_run_sct(dy_in_rsci_irdy_run_sct)
    );
  assign dy_in_rsci_idat_mxwt = dy_in_rsci_idat;
  assign dy_in_rsci_wen_comp = (~ dy_in_rsci_oswt) | dy_in_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run_dx_in_rsci
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run_dx_in_rsci (
  dx_in_rsc_dat, dx_in_rsc_vld, dx_in_rsc_rdy, run_wen, dx_in_rsci_oswt, dx_in_rsci_wen_comp,
      dx_in_rsci_idat_mxwt
);
  input [35:0] dx_in_rsc_dat;
  input dx_in_rsc_vld;
  output dx_in_rsc_rdy;
  input run_wen;
  input dx_in_rsci_oswt;
  output dx_in_rsci_wen_comp;
  output [35:0] dx_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire dx_in_rsci_irdy_run_sct;
  wire dx_in_rsci_ivld;
  wire [35:0] dx_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd14),
  .width(32'sd36)) dx_in_rsci (
      .rdy(dx_in_rsc_rdy),
      .vld(dx_in_rsc_vld),
      .dat(dx_in_rsc_dat),
      .irdy(dx_in_rsci_irdy_run_sct),
      .ivld(dx_in_rsci_ivld),
      .idat(dx_in_rsci_idat)
    );
  EdgeDetect_MagAng_run_dx_in_rsci_dx_in_wait_ctrl EdgeDetect_MagAng_run_dx_in_rsci_dx_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dx_in_rsci_iswt0(dx_in_rsci_oswt),
      .dx_in_rsci_irdy_run_sct(dx_in_rsci_irdy_run_sct)
    );
  assign dx_in_rsci_idat_mxwt = dx_in_rsci_idat;
  assign dx_in_rsci_wen_comp = (~ dx_in_rsci_oswt) | dx_in_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer_run
// ------------------------------------------------------------------


module EdgeDetect_VerDer_run (
  clk, rst, arst_n, dat_in_rsc_dat, dat_in_rsc_vld, dat_in_rsc_rdy, widthIn, heightIn,
      pix_out_rsc_dat, pix_out_rsc_vld, pix_out_rsc_rdy, dy_rsc_dat, dy_rsc_vld,
      dy_rsc_rdy, line_buf0_rsci_d_d, line_buf0_rsci_en_d, line_buf0_rsci_q_d, line_buf1_rsci_d_d,
      line_buf1_rsci_q_d, line_buf0_rsci_adr_d_pff, line_buf0_rsci_we_d_pff, line_buf0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_pff
);
  input clk;
  input rst;
  input arst_n;
  input [33:0] dat_in_rsc_dat;
  input dat_in_rsc_vld;
  output dat_in_rsc_rdy;
  input [9:0] widthIn;
  input [8:0] heightIn;
  output [31:0] pix_out_rsc_dat;
  output pix_out_rsc_vld;
  input pix_out_rsc_rdy;
  output [35:0] dy_rsc_dat;
  output dy_rsc_vld;
  input dy_rsc_rdy;
  output [63:0] line_buf0_rsci_d_d;
  output line_buf0_rsci_en_d;
  input [63:0] line_buf0_rsci_q_d;
  output [63:0] line_buf1_rsci_d_d;
  input [63:0] line_buf1_rsci_q_d;
  output [6:0] line_buf0_rsci_adr_d_pff;
  output line_buf0_rsci_we_d_pff;
  output line_buf0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire dat_in_rsci_wen_comp;
  wire [31:0] dat_in_rsci_idat_mxwt;
  wire pix_out_rsci_wen_comp;
  reg [31:0] pix_out_rsci_idat;
  wire dy_rsci_wen_comp;
  reg [8:0] dy_rsci_idat_35_27;
  wire [9:0] nl_dy_rsci_idat_35_27;
  reg [8:0] dy_rsci_idat_26_18;
  wire [9:0] nl_dy_rsci_idat_26_18;
  reg [8:0] dy_rsci_idat_17_9;
  wire [9:0] nl_dy_rsci_idat_17_9;
  reg [8:0] dy_rsci_idat_8_0;
  wire [9:0] nl_dy_rsci_idat_8_0;
  wire [2:0] fsm_output;
  wire [8:0] VCOL_if_6_mux_tmp;
  wire VCOL_VCOL_if_6_VCOL_if_6_nor_tmp;
  wire [7:0] operator_10_false_acc_tmp;
  wire [8:0] nl_operator_10_false_acc_tmp;
  wire or_dcpl_3;
  wire or_dcpl_4;
  wire or_dcpl_5;
  wire or_dcpl_7;
  wire or_dcpl_21;
  wire or_dcpl_39;
  wire or_dcpl_41;
  wire or_dcpl_43;
  reg VCOL_equal_cse_sva_1;
  wire [8:0] VROW_y_sva_mx1;
  reg [8:0] VROW_y_sva;
  reg VCOL_nor_1_itm_1;
  reg VROW_stage_0_2;
  reg [7:0] VCOL_x_9_2_sva;
  reg VROW_stage_0_1;
  reg VCOL_x_slc_VCOL_x_9_2_0_2_itm_1;
  reg VROW_stage_0_3;
  reg [8:0] VCOL_asn_itm_2;
  reg VCOL_if_slc_operator_9_false_acc_9_svs_1;
  reg VCOL_equal_cse_sva_2;
  wire VCOL_if_5_and_cse;
  reg reg_line_buf1_rsci_cgo_ir_cse;
  reg reg_dy_rsci_iswt0_cse;
  reg reg_dat_in_rsci_iswt0_cse;
  reg reg_VCOL_x_slc_VCOL_x_9_2_0_5_itm_1_cse;
  wire [31:0] VCOL_mux_4_cse;
  wire or_50_cse;
  wire and_59_rmff;
  reg [31:0] wrbuf0_pix_31_0_sva_1;
  wire [63:0] rdbuf0_pix_mux_itm;
  reg [63:0] rdbuf0_pix_sva;
  reg [31:0] pix0_sva;
  reg [31:0] pix0_sva_dfm_1;
  reg VCOL_VCOL_nand_tmp_1;
  reg VROW_asn_1_itm_1;
  reg [31:0] rdbuf1_pix_sva_63_32;
  wire pix_out_rsci_idat_mx0c1;
  wire VROW_stage_0_1_mx0w1;
  wire [7:0] VCOL_x_9_2_sva_mx1;
  wire [31:0] pix0_sva_mx0;
  wire [31:0] pix2_lpi_2_dfm_1;
  wire [31:0] pix0_sva_dfm_2_mx0;
  wire [31:0] VCOL_qr_1_lpi_2_dfm_mx0;
  wire [63:0] rdbuf0_pix_sva_dfm_mx0;
  wire [8:0] VROW_y_sva_2;
  wire [9:0] nl_VROW_y_sva_2;
  wire [8:0] operator_11_true_acc_psp_sva_1;
  wire [9:0] nl_operator_11_true_acc_psp_sva_1;
  wire VROW_and_cse;
  wire VCOL_if_4_and_cse;
  wire VCOL_if_6_unequal_tmp;
  wire operator_9_false_acc_itm_9;

  wire mux_1_nl;
  wire mux_nl;
  wire or_68_nl;
  wire nand_2_nl;
  wire mux_5_nl;
  wire and_70_nl;
  wire VROW_y_and_nl;
  wire[7:0] VCOL_VCOL_and_nl;
  wire VCOL_if_6_VCOL_if_6_or_nl;
  wire[9:0] operator_9_false_acc_nl;
  wire[10:0] nl_operator_9_false_acc_nl;
  wire VCOL_and_nl;
  wire VCOL_and_1_nl;
  wire VCOL_if_6_and_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [35:0] nl_EdgeDetect_VerDer_run_dy_rsci_inst_dy_rsci_idat;
  assign nl_EdgeDetect_VerDer_run_dy_rsci_inst_dy_rsci_idat = {dy_rsci_idat_35_27
      , dy_rsci_idat_26_18 , dy_rsci_idat_17_9 , dy_rsci_idat_8_0};
  wire  nl_EdgeDetect_VerDer_run_run_fsm_inst_VROW_C_0_tr0;
  assign nl_EdgeDetect_VerDer_run_run_fsm_inst_VROW_C_0_tr0 = ~(VROW_stage_0_1 |
      VROW_stage_0_2 | VROW_stage_0_3);
  EdgeDetect_VerDer_run_dat_in_rsci EdgeDetect_VerDer_run_dat_in_rsci_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .dat_in_rsc_dat(dat_in_rsc_dat),
      .dat_in_rsc_vld(dat_in_rsc_vld),
      .dat_in_rsc_rdy(dat_in_rsc_rdy),
      .run_wen(run_wen),
      .dat_in_rsci_oswt(reg_dat_in_rsci_iswt0_cse),
      .dat_in_rsci_wen_comp(dat_in_rsci_wen_comp),
      .dat_in_rsci_idat_mxwt(dat_in_rsci_idat_mxwt)
    );
  EdgeDetect_VerDer_run_pix_out_rsci EdgeDetect_VerDer_run_pix_out_rsci_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .pix_out_rsc_dat(pix_out_rsc_dat),
      .pix_out_rsc_vld(pix_out_rsc_vld),
      .pix_out_rsc_rdy(pix_out_rsc_rdy),
      .run_wen(run_wen),
      .pix_out_rsci_oswt(reg_dy_rsci_iswt0_cse),
      .pix_out_rsci_wen_comp(pix_out_rsci_wen_comp),
      .pix_out_rsci_idat(pix_out_rsci_idat)
    );
  EdgeDetect_VerDer_run_dy_rsci EdgeDetect_VerDer_run_dy_rsci_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .dy_rsc_dat(dy_rsc_dat),
      .dy_rsc_vld(dy_rsc_vld),
      .dy_rsc_rdy(dy_rsc_rdy),
      .run_wen(run_wen),
      .dy_rsci_oswt(reg_dy_rsci_iswt0_cse),
      .dy_rsci_wen_comp(dy_rsci_wen_comp),
      .dy_rsci_idat(nl_EdgeDetect_VerDer_run_dy_rsci_inst_dy_rsci_idat[35:0])
    );
  EdgeDetect_VerDer_run_wait_dp EdgeDetect_VerDer_run_wait_dp_inst (
      .line_buf0_rsci_en_d(line_buf0_rsci_en_d),
      .run_wen(run_wen),
      .line_buf0_rsci_cgo(reg_line_buf1_rsci_cgo_ir_cse),
      .line_buf0_rsci_cgo_ir_unreg(and_59_rmff)
    );
  EdgeDetect_VerDer_run_staller EdgeDetect_VerDer_run_staller_inst (
      .run_wen(run_wen),
      .dat_in_rsci_wen_comp(dat_in_rsci_wen_comp),
      .pix_out_rsci_wen_comp(pix_out_rsci_wen_comp),
      .dy_rsci_wen_comp(dy_rsci_wen_comp)
    );
  EdgeDetect_VerDer_run_run_fsm EdgeDetect_VerDer_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .VROW_C_0_tr0(nl_EdgeDetect_VerDer_run_run_fsm_inst_VROW_C_0_tr0)
    );
  assign VCOL_if_5_and_cse = run_wen & (~((VCOL_asn_itm_2==9'b000000000))) & VROW_stage_0_3
      & (fsm_output[1]);
  assign VROW_and_cse = run_wen & VROW_stage_0_2;
  assign VCOL_if_4_and_cse = run_wen & (or_dcpl_21 | (~ VROW_stage_0_2)) & VROW_stage_0_1;
  assign and_59_rmff = (VROW_stage_0_2 | VROW_stage_0_3) & (fsm_output[1]);
  assign or_50_cse = or_dcpl_43 | reg_VCOL_x_slc_VCOL_x_9_2_0_5_itm_1_cse;
  assign VCOL_mux_4_cse = MUX_v_32_2_2(dat_in_rsci_idat_mxwt, pix0_sva_mx0, VCOL_if_slc_operator_9_false_acc_9_svs_1);
  assign VROW_y_and_nl = VCOL_VCOL_if_6_VCOL_if_6_nor_tmp & VROW_stage_0_2;
  assign VROW_y_sva_mx1 = MUX_v_9_2_2(VROW_y_sva, VROW_y_sva_2, VROW_y_and_nl);
  assign VROW_stage_0_1_mx0w1 = VROW_stage_0_1 & or_dcpl_41;
  assign VCOL_if_6_VCOL_if_6_or_nl = VCOL_equal_cse_sva_1 | (~ VCOL_VCOL_if_6_VCOL_if_6_nor_tmp);
  assign VCOL_VCOL_and_nl = MUX_v_8_2_2(8'b00000000, operator_10_false_acc_tmp, VCOL_if_6_VCOL_if_6_or_nl);
  assign VCOL_x_9_2_sva_mx1 = MUX_v_8_2_2(VCOL_x_9_2_sva, VCOL_VCOL_and_nl, VROW_stage_0_2);
  assign rdbuf0_pix_mux_itm = MUX_v_64_2_2(line_buf0_rsci_q_d, rdbuf0_pix_sva, or_50_cse);
  assign pix0_sva_mx0 = MUX_v_32_2_2(pix0_sva_dfm_2_mx0, pix0_sva, or_dcpl_43);
  assign nl_operator_9_false_acc_nl = ({1'b1 , heightIn}) + conv_u2s_9_10(~ VROW_y_sva_mx1);
  assign operator_9_false_acc_nl = nl_operator_9_false_acc_nl[9:0];
  assign operator_9_false_acc_itm_9 = readslicef_10_1_9(operator_9_false_acc_nl);
  assign VCOL_and_nl = (~ reg_VCOL_x_slc_VCOL_x_9_2_0_5_itm_1_cse) & VCOL_VCOL_nand_tmp_1;
  assign VCOL_and_1_nl = reg_VCOL_x_slc_VCOL_x_9_2_0_5_itm_1_cse & VCOL_VCOL_nand_tmp_1;
  assign pix2_lpi_2_dfm_1 = MUX1HOT_v_32_3_2(VCOL_qr_1_lpi_2_dfm_mx0, (line_buf1_rsci_q_d[31:0]),
      rdbuf1_pix_sva_63_32, {(~ VCOL_VCOL_nand_tmp_1) , VCOL_and_nl , VCOL_and_1_nl});
  assign pix0_sva_dfm_2_mx0 = MUX_v_32_2_2(pix0_sva_dfm_1, VCOL_qr_1_lpi_2_dfm_mx0,
      VCOL_equal_cse_sva_2);
  assign VCOL_qr_1_lpi_2_dfm_mx0 = MUX_v_32_2_2((line_buf0_rsci_q_d[31:0]), (rdbuf0_pix_sva[63:32]),
      reg_VCOL_x_slc_VCOL_x_9_2_0_5_itm_1_cse);
  assign rdbuf0_pix_sva_dfm_mx0 = MUX_v_64_2_2(line_buf0_rsci_q_d, rdbuf0_pix_sva,
      reg_VCOL_x_slc_VCOL_x_9_2_0_5_itm_1_cse);
  assign nl_VROW_y_sva_2 = VROW_y_sva + 9'b000000001;
  assign VROW_y_sva_2 = nl_VROW_y_sva_2[8:0];
  assign VCOL_if_6_unequal_tmp = VCOL_x_9_2_sva != (operator_11_true_acc_psp_sva_1[7:0]);
  assign VCOL_VCOL_if_6_VCOL_if_6_nor_tmp = ~(VCOL_if_6_unequal_tmp | (operator_11_true_acc_psp_sva_1[8]));
  assign nl_operator_11_true_acc_psp_sva_1 = conv_u2s_8_9(widthIn[9:2]) + 9'b111111111;
  assign operator_11_true_acc_psp_sva_1 = nl_operator_11_true_acc_psp_sva_1[8:0];
  assign nl_operator_10_false_acc_tmp = VCOL_x_9_2_sva + 8'b00000001;
  assign operator_10_false_acc_tmp = nl_operator_10_false_acc_tmp[7:0];
  assign VCOL_if_6_and_nl = (~ VCOL_equal_cse_sva_1) & VCOL_VCOL_if_6_VCOL_if_6_nor_tmp;
  assign VCOL_if_6_mux_tmp = MUX_v_9_2_2(VROW_y_sva, VROW_y_sva_2, VCOL_if_6_and_nl);
  assign or_dcpl_3 = (VROW_y_sva[5:4]!=2'b00);
  assign or_dcpl_4 = (VROW_y_sva[8:7]!=2'b00);
  assign or_dcpl_5 = or_dcpl_4 | (VROW_y_sva[6]);
  assign or_dcpl_7 = or_dcpl_5 | or_dcpl_3 | (VROW_y_sva[3:0]!=4'b0000);
  assign or_dcpl_21 = ~(VCOL_VCOL_if_6_VCOL_if_6_nor_tmp & VCOL_equal_cse_sva_1);
  assign or_dcpl_39 = (VCOL_asn_itm_2!=9'b000000000);
  assign or_dcpl_41 = ~(VCOL_VCOL_if_6_VCOL_if_6_nor_tmp & VCOL_equal_cse_sva_1 &
      VROW_stage_0_2);
  assign or_dcpl_43 = (~ VROW_stage_0_3) | VROW_asn_1_itm_1;
  assign pix_out_rsci_idat_mx0c1 = or_dcpl_39 & VROW_stage_0_3 & (~ reg_VCOL_x_slc_VCOL_x_9_2_0_5_itm_1_cse)
      & (fsm_output[1]);
  assign line_buf0_rsci_adr_d_pff = VCOL_x_9_2_sva[7:1];
  assign line_buf0_rsci_d_d = {VCOL_mux_4_cse , wrbuf0_pix_31_0_sva_1};
  assign line_buf0_rsci_we_d_pff = VROW_stage_0_2 & VCOL_x_slc_VCOL_x_9_2_0_2_itm_1
      & (fsm_output[1]);
  assign line_buf0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_pff = VROW_stage_0_2
      & (~ VCOL_x_slc_VCOL_x_9_2_0_2_itm_1) & (fsm_output[1]);
  assign line_buf1_rsci_d_d = rdbuf0_pix_mux_itm;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dy_rsci_idat_35_27 <= 9'b000000000;
      dy_rsci_idat_8_0 <= 9'b000000000;
      dy_rsci_idat_26_18 <= 9'b000000000;
      dy_rsci_idat_17_9 <= 9'b000000000;
    end
    else if ( rst ) begin
      dy_rsci_idat_35_27 <= 9'b000000000;
      dy_rsci_idat_8_0 <= 9'b000000000;
      dy_rsci_idat_26_18 <= 9'b000000000;
      dy_rsci_idat_17_9 <= 9'b000000000;
    end
    else if ( VCOL_if_5_and_cse ) begin
      dy_rsci_idat_35_27 <= nl_dy_rsci_idat_35_27[8:0];
      dy_rsci_idat_8_0 <= nl_dy_rsci_idat_8_0[8:0];
      dy_rsci_idat_26_18 <= nl_dy_rsci_idat_26_18[8:0];
      dy_rsci_idat_17_9 <= nl_dy_rsci_idat_17_9[8:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      pix_out_rsci_idat <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      pix_out_rsci_idat <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & ((or_dcpl_39 & VROW_stage_0_3 & reg_VCOL_x_slc_VCOL_x_9_2_0_5_itm_1_cse
        & (fsm_output[1])) | pix_out_rsci_idat_mx0c1) ) begin
      pix_out_rsci_idat <= MUX_v_32_2_2((rdbuf0_pix_sva_dfm_mx0[63:32]), (rdbuf0_pix_sva_dfm_mx0[31:0]),
          pix_out_rsci_idat_mx0c1);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      VROW_asn_1_itm_1 <= 1'b0;
      VCOL_asn_itm_2 <= 9'b000000000;
    end
    else if ( rst ) begin
      VROW_asn_1_itm_1 <= 1'b0;
      VCOL_asn_itm_2 <= 9'b000000000;
    end
    else if ( VROW_and_cse ) begin
      VROW_asn_1_itm_1 <= VCOL_equal_cse_sva_1 & VCOL_VCOL_if_6_VCOL_if_6_nor_tmp;
      VCOL_asn_itm_2 <= VROW_y_sva;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      VROW_y_sva <= 9'b000000000;
    end
    else if ( rst ) begin
      VROW_y_sva <= 9'b000000000;
    end
    else if ( (~((~(VROW_stage_0_2 & (~ (operator_11_true_acc_psp_sva_1[8])) & (~
        VCOL_if_6_unequal_tmp))) & (fsm_output[1]))) & run_wen ) begin
      VROW_y_sva <= MUX_v_9_2_2(9'b000000000, VROW_y_sva_mx1, (fsm_output[1]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      VROW_stage_0_1 <= 1'b0;
      VROW_stage_0_2 <= 1'b0;
      VROW_stage_0_3 <= 1'b0;
      reg_line_buf1_rsci_cgo_ir_cse <= 1'b0;
      reg_dy_rsci_iswt0_cse <= 1'b0;
      reg_dat_in_rsci_iswt0_cse <= 1'b0;
    end
    else if ( rst ) begin
      VROW_stage_0_1 <= 1'b0;
      VROW_stage_0_2 <= 1'b0;
      VROW_stage_0_3 <= 1'b0;
      reg_line_buf1_rsci_cgo_ir_cse <= 1'b0;
      reg_dy_rsci_iswt0_cse <= 1'b0;
      reg_dat_in_rsci_iswt0_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      VROW_stage_0_1 <= VROW_stage_0_1_mx0w1 | (~ (fsm_output[1]));
      VROW_stage_0_2 <= VROW_stage_0_1_mx0w1 & (fsm_output[1]);
      VROW_stage_0_3 <= VROW_stage_0_2 & (fsm_output[1]);
      reg_line_buf1_rsci_cgo_ir_cse <= and_59_rmff;
      reg_dy_rsci_iswt0_cse <= or_dcpl_39 & VROW_stage_0_3 & (fsm_output[1]);
      reg_dat_in_rsci_iswt0_cse <= or_dcpl_41 & VROW_stage_0_1 & (~ operator_9_false_acc_itm_9)
          & (fsm_output[1]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      VCOL_x_9_2_sva <= 8'b00000000;
    end
    else if ( rst ) begin
      VCOL_x_9_2_sva <= 8'b00000000;
    end
    else if ( (VROW_stage_0_2 | (~ (fsm_output[1]))) & run_wen ) begin
      VCOL_x_9_2_sva <= MUX_v_8_2_2(8'b00000000, VCOL_x_9_2_sva_mx1, (fsm_output[1]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      VCOL_equal_cse_sva_1 <= 1'b0;
      VCOL_x_slc_VCOL_x_9_2_0_2_itm_1 <= 1'b0;
      VCOL_if_slc_operator_9_false_acc_9_svs_1 <= 1'b0;
    end
    else if ( rst ) begin
      VCOL_equal_cse_sva_1 <= 1'b0;
      VCOL_x_slc_VCOL_x_9_2_0_2_itm_1 <= 1'b0;
      VCOL_if_slc_operator_9_false_acc_9_svs_1 <= 1'b0;
    end
    else if ( VCOL_if_4_and_cse ) begin
      VCOL_equal_cse_sva_1 <= VROW_y_sva_mx1 == heightIn;
      VCOL_x_slc_VCOL_x_9_2_0_2_itm_1 <= VCOL_x_9_2_sva_mx1[0];
      VCOL_if_slc_operator_9_false_acc_9_svs_1 <= operator_9_false_acc_itm_9;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      pix0_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      pix0_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( VROW_stage_0_3 & (~ VROW_asn_1_itm_1) & (~ VROW_stage_0_2) & operator_9_false_acc_itm_9
        & run_wen & VROW_stage_0_1 ) begin
      pix0_sva <= pix0_sva_mx0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rdbuf0_pix_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      rdbuf0_pix_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( (~ VROW_asn_1_itm_1) & VROW_stage_0_3 & (~ reg_VCOL_x_slc_VCOL_x_9_2_0_5_itm_1_cse)
        & run_wen ) begin
      rdbuf0_pix_sva <= rdbuf0_pix_mux_itm;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      VCOL_VCOL_nand_tmp_1 <= 1'b0;
    end
    else if ( rst ) begin
      VCOL_VCOL_nand_tmp_1 <= 1'b0;
    end
    else if ( run_wen & or_dcpl_7 & VROW_stage_0_2 ) begin
      VCOL_VCOL_nand_tmp_1 <= ~((VROW_y_sva[0]) & VCOL_nor_1_itm_1);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rdbuf1_pix_sva_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      rdbuf1_pix_sva_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & mux_1_nl & (VCOL_x_9_2_sva[0]) & (~ or_50_cse) ) begin
      rdbuf1_pix_sva_63_32 <= line_buf1_rsci_q_d[63:32];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_VCOL_x_slc_VCOL_x_9_2_0_5_itm_1_cse <= 1'b0;
    end
    else if ( rst ) begin
      reg_VCOL_x_slc_VCOL_x_9_2_0_5_itm_1_cse <= 1'b0;
    end
    else if ( run_wen & (or_dcpl_4 | (VROW_y_sva[6:2]!=5'b00000) | (VROW_stage_0_1
        & (~ VCOL_VCOL_if_6_VCOL_if_6_nor_tmp) & (operator_10_false_acc_tmp[0]))
        | (VROW_y_sva[1]) | VCOL_equal_cse_sva_1 | (VROW_y_sva[0])) & VROW_stage_0_2
        ) begin
      reg_VCOL_x_slc_VCOL_x_9_2_0_5_itm_1_cse <= VCOL_x_9_2_sva[0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      pix0_sva_dfm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      pix0_sva_dfm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( (VCOL_equal_cse_sva_2 | VROW_asn_1_itm_1 | (~(VCOL_if_slc_operator_9_false_acc_9_svs_1
        & VROW_stage_0_3))) & run_wen ) begin
      pix0_sva_dfm_1 <= VCOL_mux_4_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      VCOL_equal_cse_sva_2 <= 1'b0;
    end
    else if ( rst ) begin
      VCOL_equal_cse_sva_2 <= 1'b0;
    end
    else if ( run_wen & ((VROW_stage_0_1 & operator_9_false_acc_itm_9 & or_dcpl_21)
        | or_dcpl_5 | or_dcpl_3 | (VROW_y_sva[3:0]!=4'b0000)) & VROW_stage_0_2 )
        begin
      VCOL_equal_cse_sva_2 <= VCOL_equal_cse_sva_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      wrbuf0_pix_31_0_sva_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      wrbuf0_pix_31_0_sva_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & (~((~ (operator_10_false_acc_tmp[0])) | VCOL_VCOL_if_6_VCOL_if_6_nor_tmp))
        & VROW_stage_0_2 & VROW_stage_0_1 & (~ (VCOL_x_9_2_sva[0])) ) begin
      wrbuf0_pix_31_0_sva_1 <= VCOL_mux_4_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      VCOL_nor_1_itm_1 <= 1'b0;
    end
    else if ( rst ) begin
      VCOL_nor_1_itm_1 <= 1'b0;
    end
    else if ( run_wen & mux_5_nl & VROW_stage_0_1 ) begin
      VCOL_nor_1_itm_1 <= ~((VROW_y_sva_mx1[8:1]!=8'b00000000));
    end
  end
  assign nl_dy_rsci_idat_35_27  = ({1'b1 , (pix2_lpi_2_dfm_1[31:24])}) + conv_u2s_8_9(~
      (pix0_sva_dfm_2_mx0[31:24])) + 9'b000000001;
  assign nl_dy_rsci_idat_8_0  = ({1'b1 , (pix2_lpi_2_dfm_1[7:0])}) + conv_u2s_8_9(~
      (pix0_sva_dfm_2_mx0[7:0])) + 9'b000000001;
  assign nl_dy_rsci_idat_26_18  = ({1'b1 , (pix2_lpi_2_dfm_1[23:16])}) + conv_u2s_8_9(~
      (pix0_sva_dfm_2_mx0[23:16])) + 9'b000000001;
  assign nl_dy_rsci_idat_17_9  = ({1'b1 , (pix2_lpi_2_dfm_1[15:8])}) + conv_u2s_8_9(~
      (pix0_sva_dfm_2_mx0[15:8])) + 9'b000000001;
  assign or_68_nl = (~((~ (operator_10_false_acc_tmp[0])) | VCOL_VCOL_if_6_VCOL_if_6_nor_tmp
      | (~ VROW_stage_0_1))) | (VROW_y_sva[8:1]!=8'b00000000);
  assign nand_2_nl = ~(VCOL_nor_1_itm_1 & ((~ (operator_10_false_acc_tmp[0])) | VCOL_VCOL_if_6_VCOL_if_6_nor_tmp
      | (~ VROW_stage_0_1)));
  assign mux_nl = MUX_s_1_2_2(or_68_nl, nand_2_nl, VROW_y_sva[0]);
  assign mux_1_nl = MUX_s_1_2_2(VROW_stage_0_1, mux_nl, VROW_stage_0_2);
  assign and_70_nl = ((VCOL_if_6_mux_tmp!=9'b000000000)) & or_dcpl_21;
  assign mux_5_nl = MUX_s_1_2_2(or_dcpl_7, and_70_nl, VROW_stage_0_2);

  function automatic [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | (input_1 & {32{sel[1]}});
    result = result | (input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_10 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_HorDer_run
// ------------------------------------------------------------------


module EdgeDetect_HorDer_run (
  clk, rst, arst_n, pix_in_rsc_dat, pix_in_rsc_vld, pix_in_rsc_rdy, widthIn, heightIn,
      pix_out_rsc_dat, pix_out_rsc_vld, pix_out_rsc_rdy, dx_rsc_dat, dx_rsc_vld,
      dx_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] pix_in_rsc_dat;
  input pix_in_rsc_vld;
  output pix_in_rsc_rdy;
  input [9:0] widthIn;
  input [8:0] heightIn;
  output [31:0] pix_out_rsc_dat;
  output pix_out_rsc_vld;
  input pix_out_rsc_rdy;
  output [35:0] dx_rsc_dat;
  output dx_rsc_vld;
  input dx_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire pix_in_rsci_wen_comp;
  wire [31:0] pix_in_rsci_idat_mxwt;
  wire pix_out_rsci_wen_comp;
  wire dx_rsci_wen_comp;
  reg [7:0] pix_out_rsci_idat_31_24;
  reg [7:0] pix_out_rsci_idat_23_16;
  reg [7:0] pix_out_rsci_idat_15_8;
  reg [7:0] pix_out_rsci_idat_7_0;
  reg [8:0] dx_rsci_idat_35_27;
  wire [9:0] nl_dx_rsci_idat_35_27;
  reg [8:0] dx_rsci_idat_26_18;
  reg [8:0] dx_rsci_idat_17_9;
  reg [8:0] dx_rsci_idat_8_0;
  wire [2:0] fsm_output;
  wire HROW_equal_tmp;
  wire [7:0] operator_10_false_acc_tmp;
  wire [8:0] nl_operator_10_false_acc_tmp;
  wire HCOL_else_1_HCOL_else_1_if_HCOL_else_1_if_equal_tmp;
  wire or_dcpl_1;
  wire and_dcpl;
  wire and_dcpl_9;
  wire or_dcpl_5;
  wire or_dcpl_10;
  wire mux_tmp_1;
  wire or_dcpl_14;
  wire [7:0] HCOL_x_9_2_sva_mx1;
  reg HROW_stage_0_2;
  reg HROW_stage_0_1;
  reg [7:0] HCOL_x_9_2_sva;
  reg HCOL_unequal_tmp_1;
  reg HCOL_if_slc_operator_11_true_acc_8_svs_1;
  wire HCOL_if_2_and_cse;
  reg reg_dx_rsci_iswt0_cse;
  reg reg_pix_in_rsci_iswt0_cse;
  wire [7:0] HCOL_if_1_for_1_mux_8_cse;
  wire or_29_tmp;
  wire [31:0] pix_sva_dfm_mx0;
  reg [31:0] pix_sva;
  reg [7:0] win_5_sva;
  reg [7:0] win_6_sva;
  reg [7:0] win_7_sva;
  reg [7:0] win_8_sva;
  reg [8:0] HROW_y_sva;
  reg [8:0] operator_8_false_2_acc_1_itm_1;
  wire [9:0] nl_operator_8_false_2_acc_1_itm_1;
  reg [8:0] operator_8_false_2_acc_2_itm_1;
  wire [9:0] nl_operator_8_false_2_acc_2_itm_1;
  reg [8:0] operator_8_false_2_acc_3_itm_1;
  wire [9:0] nl_operator_8_false_2_acc_3_itm_1;
  wire HROW_stage_0_1_mx0w1;
  wire [7:0] win_5_sva_mx0;
  wire HCOL_unequal_tmp_1_1;
  wire operator_8_false_2_and_cse;
  wire HCOL_and_5_cse;
  wire win_and_2_cse;
  wire nand_12_cse;
  wire operator_11_true_acc_itm_8_1;

  wire[7:0] win_mux_6_nl;
  wire nand_9_nl;
  wire[8:0] HROW_acc_nl;
  wire[9:0] nl_HROW_acc_nl;
  wire mux_2_nl;
  wire mux_nl;
  wire or_nl;
  wire nor_nl;
  wire[7:0] HCOL_HCOL_mux1h_nl;
  wire HCOL_and_nl;
  wire HCOL_and_4_nl;
  wire[7:0] HCOL_if_1_for_1_mux_6_nl;
  wire[7:0] HCOL_if_1_for_1_mux_4_nl;
  wire[7:0] HCOL_HCOL_and_nl;
  wire HCOL_if_3_HCOL_if_3_or_nl;
  wire win_and_nl;
  wire win_and_1_nl;
  wire[8:0] operator_11_true_acc_nl;
  wire[9:0] nl_operator_11_true_acc_nl;
  wire[8:0] operator_9_false_acc_nl;
  wire[9:0] nl_operator_9_false_acc_nl;
  wire nor_3_nl;
  wire or_16_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_EdgeDetect_HorDer_run_pix_out_rsci_inst_pix_out_rsci_idat;
  assign nl_EdgeDetect_HorDer_run_pix_out_rsci_inst_pix_out_rsci_idat = {pix_out_rsci_idat_31_24
      , pix_out_rsci_idat_23_16 , pix_out_rsci_idat_15_8 , pix_out_rsci_idat_7_0};
  wire [35:0] nl_EdgeDetect_HorDer_run_dx_rsci_inst_dx_rsci_idat;
  assign nl_EdgeDetect_HorDer_run_dx_rsci_inst_dx_rsci_idat = {dx_rsci_idat_35_27
      , dx_rsci_idat_26_18 , dx_rsci_idat_17_9 , dx_rsci_idat_8_0};
  wire  nl_EdgeDetect_HorDer_run_run_fsm_inst_HROW_C_0_tr0;
  assign nl_EdgeDetect_HorDer_run_run_fsm_inst_HROW_C_0_tr0 = ~(HROW_stage_0_2 |
      HROW_stage_0_1);
  EdgeDetect_HorDer_run_pix_in_rsci EdgeDetect_HorDer_run_pix_in_rsci_inst (
      .pix_in_rsc_dat(pix_in_rsc_dat),
      .pix_in_rsc_vld(pix_in_rsc_vld),
      .pix_in_rsc_rdy(pix_in_rsc_rdy),
      .run_wen(run_wen),
      .pix_in_rsci_oswt(reg_pix_in_rsci_iswt0_cse),
      .pix_in_rsci_wen_comp(pix_in_rsci_wen_comp),
      .pix_in_rsci_idat_mxwt(pix_in_rsci_idat_mxwt)
    );
  EdgeDetect_HorDer_run_pix_out_rsci EdgeDetect_HorDer_run_pix_out_rsci_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .pix_out_rsc_dat(pix_out_rsc_dat),
      .pix_out_rsc_vld(pix_out_rsc_vld),
      .pix_out_rsc_rdy(pix_out_rsc_rdy),
      .run_wen(run_wen),
      .pix_out_rsci_oswt(reg_dx_rsci_iswt0_cse),
      .pix_out_rsci_wen_comp(pix_out_rsci_wen_comp),
      .pix_out_rsci_idat(nl_EdgeDetect_HorDer_run_pix_out_rsci_inst_pix_out_rsci_idat[31:0])
    );
  EdgeDetect_HorDer_run_dx_rsci EdgeDetect_HorDer_run_dx_rsci_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .dx_rsc_dat(dx_rsc_dat),
      .dx_rsc_vld(dx_rsc_vld),
      .dx_rsc_rdy(dx_rsc_rdy),
      .run_wen(run_wen),
      .dx_rsci_oswt(reg_dx_rsci_iswt0_cse),
      .dx_rsci_wen_comp(dx_rsci_wen_comp),
      .dx_rsci_idat(nl_EdgeDetect_HorDer_run_dx_rsci_inst_dx_rsci_idat[35:0])
    );
  EdgeDetect_HorDer_run_staller EdgeDetect_HorDer_run_staller_inst (
      .run_wen(run_wen),
      .pix_in_rsci_wen_comp(pix_in_rsci_wen_comp),
      .pix_out_rsci_wen_comp(pix_out_rsci_wen_comp),
      .dx_rsci_wen_comp(dx_rsci_wen_comp)
    );
  EdgeDetect_HorDer_run_run_fsm EdgeDetect_HorDer_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .HROW_C_0_tr0(nl_EdgeDetect_HorDer_run_run_fsm_inst_HROW_C_0_tr0)
    );
  assign HCOL_if_2_and_cse = run_wen & (~(and_dcpl_9 & (HCOL_x_9_2_sva[5:0]==6'b000000)))
      & HROW_stage_0_2 & (fsm_output[1]);
  assign nand_12_cse = ~(HCOL_else_1_HCOL_else_1_if_HCOL_else_1_if_equal_tmp & HROW_stage_0_2);
  assign mux_2_nl = MUX_s_1_2_2(HCOL_else_1_HCOL_else_1_if_HCOL_else_1_if_equal_tmp,
      mux_tmp_1, HCOL_x_9_2_sva[0]);
  assign win_and_2_cse = run_wen & and_dcpl & (~(mux_2_nl & HCOL_unequal_tmp_1))
      & HROW_stage_0_2;
  assign HCOL_if_1_for_1_mux_8_cse = MUX_v_8_2_2((pix_sva_dfm_mx0[15:8]), win_6_sva,
      or_dcpl_14);
  assign or_nl = (HCOL_x_9_2_sva!=8'b00000000);
  assign nor_nl = ~((~((operator_10_false_acc_tmp!=8'b00000000))) | HCOL_else_1_HCOL_else_1_if_HCOL_else_1_if_equal_tmp);
  assign mux_nl = MUX_s_1_2_2(or_nl, nor_nl, HROW_stage_0_2);
  assign operator_8_false_2_and_cse = run_wen & mux_nl & HROW_stage_0_1;
  assign HCOL_and_5_cse = run_wen & and_dcpl;
  assign HCOL_if_3_HCOL_if_3_or_nl = HROW_equal_tmp | (~ HCOL_else_1_HCOL_else_1_if_HCOL_else_1_if_equal_tmp);
  assign HCOL_HCOL_and_nl = MUX_v_8_2_2(8'b00000000, operator_10_false_acc_tmp, HCOL_if_3_HCOL_if_3_or_nl);
  assign HCOL_x_9_2_sva_mx1 = MUX_v_8_2_2(HCOL_x_9_2_sva, HCOL_HCOL_and_nl, HROW_stage_0_2);
  assign HROW_stage_0_1_mx0w1 = HROW_stage_0_1 & or_dcpl_5;
  assign or_29_tmp = or_dcpl_10 | (HCOL_x_9_2_sva[5:1]!=5'b00000) | (~((HCOL_x_9_2_sva[0])
      & HCOL_unequal_tmp_1));
  assign win_and_nl = (~ or_29_tmp) & HROW_stage_0_2;
  assign win_and_1_nl = or_29_tmp & HROW_stage_0_2;
  assign win_5_sva_mx0 = MUX1HOT_v_8_3_2(win_5_sva, win_7_sva, (pix_sva_dfm_mx0[7:0]),
      {(~ HROW_stage_0_2) , win_and_nl , win_and_1_nl});
  assign HCOL_unequal_tmp_1_1 = ~((HCOL_x_9_2_sva_mx1==8'b00000001));
  assign nl_operator_11_true_acc_nl = ({1'b1 , (widthIn[9:2])}) + conv_u2s_8_9(~
      HCOL_x_9_2_sva_mx1);
  assign operator_11_true_acc_nl = nl_operator_11_true_acc_nl[8:0];
  assign operator_11_true_acc_itm_8_1 = readslicef_9_1_8(operator_11_true_acc_nl);
  assign pix_sva_dfm_mx0 = MUX_v_32_2_2(pix_in_rsci_idat_mxwt, pix_sva, HCOL_if_slc_operator_11_true_acc_8_svs_1);
  assign nl_operator_10_false_acc_tmp = HCOL_x_9_2_sva + 8'b00000001;
  assign operator_10_false_acc_tmp = nl_operator_10_false_acc_tmp[7:0];
  assign nl_operator_9_false_acc_nl = heightIn + 9'b111111111;
  assign operator_9_false_acc_nl = nl_operator_9_false_acc_nl[8:0];
  assign HROW_equal_tmp = HROW_y_sva == operator_9_false_acc_nl;
  assign HCOL_else_1_HCOL_else_1_if_HCOL_else_1_if_equal_tmp = HCOL_x_9_2_sva ==
      (widthIn[9:2]);
  assign or_dcpl_1 = ~(HCOL_else_1_HCOL_else_1_if_HCOL_else_1_if_equal_tmp & HROW_stage_0_2
      & HROW_equal_tmp);
  assign and_dcpl = or_dcpl_1 & HROW_stage_0_1;
  assign and_dcpl_9 = ~((HCOL_x_9_2_sva[7:6]!=2'b00));
  assign or_dcpl_5 = nand_12_cse | (~ HROW_equal_tmp);
  assign or_dcpl_10 = (HCOL_x_9_2_sva[7:6]!=2'b00);
  assign nor_3_nl = ~((HCOL_x_9_2_sva[7:1]!=7'b0000000));
  assign or_16_nl = (HCOL_x_9_2_sva[7:1]!=7'b0000000);
  assign mux_tmp_1 = MUX_s_1_2_2(nor_3_nl, or_16_nl, HCOL_else_1_HCOL_else_1_if_HCOL_else_1_if_equal_tmp);
  assign or_dcpl_14 = ~((~(and_dcpl_9 & (HCOL_x_9_2_sva[5:0]==6'b000001) & HCOL_unequal_tmp_1))
      & HROW_stage_0_2);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      HCOL_x_9_2_sva <= 8'b00000000;
    end
    else if ( rst ) begin
      HCOL_x_9_2_sva <= 8'b00000000;
    end
    else if ( (HROW_stage_0_2 | (~ (fsm_output[1]))) & run_wen ) begin
      HCOL_x_9_2_sva <= MUX_v_8_2_2(8'b00000000, HCOL_x_9_2_sva_mx1, (fsm_output[1]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dx_rsci_idat_35_27 <= 9'b000000000;
      dx_rsci_idat_8_0 <= 9'b000000000;
      dx_rsci_idat_26_18 <= 9'b000000000;
      dx_rsci_idat_17_9 <= 9'b000000000;
      pix_out_rsci_idat_31_24 <= 8'b00000000;
      pix_out_rsci_idat_7_0 <= 8'b00000000;
      pix_out_rsci_idat_23_16 <= 8'b00000000;
      pix_out_rsci_idat_15_8 <= 8'b00000000;
    end
    else if ( rst ) begin
      dx_rsci_idat_35_27 <= 9'b000000000;
      dx_rsci_idat_8_0 <= 9'b000000000;
      dx_rsci_idat_26_18 <= 9'b000000000;
      dx_rsci_idat_17_9 <= 9'b000000000;
      pix_out_rsci_idat_31_24 <= 8'b00000000;
      pix_out_rsci_idat_7_0 <= 8'b00000000;
      pix_out_rsci_idat_23_16 <= 8'b00000000;
      pix_out_rsci_idat_15_8 <= 8'b00000000;
    end
    else if ( HCOL_if_2_and_cse ) begin
      dx_rsci_idat_35_27 <= nl_dx_rsci_idat_35_27[8:0];
      dx_rsci_idat_8_0 <= operator_8_false_2_acc_3_itm_1;
      dx_rsci_idat_26_18 <= operator_8_false_2_acc_1_itm_1;
      dx_rsci_idat_17_9 <= operator_8_false_2_acc_2_itm_1;
      pix_out_rsci_idat_31_24 <= win_8_sva;
      pix_out_rsci_idat_7_0 <= win_5_sva;
      pix_out_rsci_idat_23_16 <= win_7_sva;
      pix_out_rsci_idat_15_8 <= win_6_sva;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      HROW_stage_0_1 <= 1'b0;
      HROW_stage_0_2 <= 1'b0;
      reg_dx_rsci_iswt0_cse <= 1'b0;
      reg_pix_in_rsci_iswt0_cse <= 1'b0;
    end
    else if ( rst ) begin
      HROW_stage_0_1 <= 1'b0;
      HROW_stage_0_2 <= 1'b0;
      reg_dx_rsci_iswt0_cse <= 1'b0;
      reg_pix_in_rsci_iswt0_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      HROW_stage_0_1 <= HROW_stage_0_1_mx0w1 | (~ (fsm_output[1]));
      HROW_stage_0_2 <= HROW_stage_0_1_mx0w1 & (fsm_output[1]);
      reg_dx_rsci_iswt0_cse <= (or_dcpl_10 | (HCOL_x_9_2_sva[5:0]!=6'b000000)) &
          HROW_stage_0_2 & (fsm_output[1]);
      reg_pix_in_rsci_iswt0_cse <= or_dcpl_5 & HROW_stage_0_1 & (~ operator_11_true_acc_itm_8_1)
          & (fsm_output[1]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      HROW_y_sva <= 9'b000000000;
    end
    else if ( rst ) begin
      HROW_y_sva <= 9'b000000000;
    end
    else if ( (~(nand_12_cse & (fsm_output[1]))) & run_wen ) begin
      HROW_y_sva <= MUX_v_9_2_2(9'b000000000, HROW_acc_nl, (fsm_output[1]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      win_7_sva <= 8'b00000000;
      win_8_sva <= 8'b00000000;
      win_6_sva <= 8'b00000000;
    end
    else if ( rst ) begin
      win_7_sva <= 8'b00000000;
      win_8_sva <= 8'b00000000;
      win_6_sva <= 8'b00000000;
    end
    else if ( win_and_2_cse ) begin
      win_7_sva <= pix_sva_dfm_mx0[23:16];
      win_8_sva <= pix_sva_dfm_mx0[31:24];
      win_6_sva <= pix_sva_dfm_mx0[15:8];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_8_false_2_acc_3_itm_1 <= 9'b000000000;
      operator_8_false_2_acc_1_itm_1 <= 9'b000000000;
      operator_8_false_2_acc_2_itm_1 <= 9'b000000000;
    end
    else if ( rst ) begin
      operator_8_false_2_acc_3_itm_1 <= 9'b000000000;
      operator_8_false_2_acc_1_itm_1 <= 9'b000000000;
      operator_8_false_2_acc_2_itm_1 <= 9'b000000000;
    end
    else if ( operator_8_false_2_and_cse ) begin
      operator_8_false_2_acc_3_itm_1 <= nl_operator_8_false_2_acc_3_itm_1[8:0];
      operator_8_false_2_acc_1_itm_1 <= nl_operator_8_false_2_acc_1_itm_1[8:0];
      operator_8_false_2_acc_2_itm_1 <= nl_operator_8_false_2_acc_2_itm_1[8:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      win_5_sva <= 8'b00000000;
    end
    else if ( rst ) begin
      win_5_sva <= 8'b00000000;
    end
    else if ( ((operator_10_false_acc_tmp!=8'b00000000)) & (~ HCOL_else_1_HCOL_else_1_if_HCOL_else_1_if_equal_tmp)
        & run_wen & HROW_stage_0_1 & HROW_stage_0_2 ) begin
      win_5_sva <= win_5_sva_mx0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      HCOL_unequal_tmp_1 <= 1'b0;
      HCOL_if_slc_operator_11_true_acc_8_svs_1 <= 1'b0;
    end
    else if ( rst ) begin
      HCOL_unequal_tmp_1 <= 1'b0;
      HCOL_if_slc_operator_11_true_acc_8_svs_1 <= 1'b0;
    end
    else if ( HCOL_and_5_cse ) begin
      HCOL_unequal_tmp_1 <= HCOL_unequal_tmp_1_1;
      HCOL_if_slc_operator_11_true_acc_8_svs_1 <= operator_11_true_acc_itm_8_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      pix_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      pix_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & or_dcpl_1 & HROW_stage_0_1 & operator_11_true_acc_itm_8_1
        & (~(HCOL_if_slc_operator_11_true_acc_8_svs_1 | (~ HROW_stage_0_2))) ) begin
      pix_sva <= pix_in_rsci_idat_mxwt;
    end
  end
  assign nand_9_nl = ~(mux_tmp_1 & HCOL_unequal_tmp_1);
  assign win_mux_6_nl = MUX_v_8_2_2(win_7_sva, (pix_sva_dfm_mx0[7:0]), nand_9_nl);
  assign nl_dx_rsci_idat_35_27  = ({1'b1 , win_7_sva}) + conv_u2s_8_9(~ win_mux_6_nl)
      + 9'b000000001;
  assign nl_HROW_acc_nl = HROW_y_sva + 9'b000000001;
  assign HROW_acc_nl = nl_HROW_acc_nl[8:0];
  assign HCOL_and_nl = (~ HROW_stage_0_2) & HCOL_unequal_tmp_1_1;
  assign HCOL_and_4_nl = HROW_stage_0_2 & HCOL_unequal_tmp_1_1;
  assign HCOL_HCOL_mux1h_nl = MUX1HOT_v_8_3_2(HCOL_if_1_for_1_mux_8_cse, pix_out_rsci_idat_31_24,
      win_8_sva, {(~ HCOL_unequal_tmp_1_1) , HCOL_and_nl , HCOL_and_4_nl});
  assign nl_operator_8_false_2_acc_3_itm_1  = ({1'b1 , HCOL_HCOL_mux1h_nl}) + conv_u2s_8_9(~
      HCOL_if_1_for_1_mux_8_cse) + 9'b000000001;
  assign HCOL_if_1_for_1_mux_6_nl = MUX_v_8_2_2((pix_sva_dfm_mx0[31:24]), win_8_sva,
      or_dcpl_14);
  assign nl_operator_8_false_2_acc_1_itm_1  = ({1'b1 , HCOL_if_1_for_1_mux_8_cse})
      + conv_u2s_8_9(~ HCOL_if_1_for_1_mux_6_nl) + 9'b000000001;
  assign HCOL_if_1_for_1_mux_4_nl = MUX_v_8_2_2((pix_sva_dfm_mx0[23:16]), win_7_sva,
      or_dcpl_14);
  assign nl_operator_8_false_2_acc_2_itm_1  = ({1'b1 , win_5_sva_mx0}) + conv_u2s_8_9(~
      HCOL_if_1_for_1_mux_4_nl) + 9'b000000001;

  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng_run
// ------------------------------------------------------------------


module EdgeDetect_MagAng_run (
  clk, rst, arst_n, dx_in_rsc_dat, dx_in_rsc_vld, dx_in_rsc_rdy, dy_in_rsc_dat, dy_in_rsc_vld,
      dy_in_rsc_rdy, pix_in_rsc_dat, pix_in_rsc_vld, pix_in_rsc_rdy, widthIn, heightIn,
      sw_in, crc32_pix_in_triosy_lz, crc32_dat_out_triosy_lz, dat_out_rsc_dat, dat_out_rsc_vld,
      dat_out_rsc_rdy, crc32_pix_in_rsci_idat, crc32_dat_out_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  input [35:0] dx_in_rsc_dat;
  input dx_in_rsc_vld;
  output dx_in_rsc_rdy;
  input [35:0] dy_in_rsc_dat;
  input dy_in_rsc_vld;
  output dy_in_rsc_rdy;
  input [31:0] pix_in_rsc_dat;
  input pix_in_rsc_vld;
  output pix_in_rsc_rdy;
  input [9:0] widthIn;
  input [8:0] heightIn;
  input sw_in;
  output crc32_pix_in_triosy_lz;
  output crc32_dat_out_triosy_lz;
  output [33:0] dat_out_rsc_dat;
  output dat_out_rsc_vld;
  input dat_out_rsc_rdy;
  output [31:0] crc32_pix_in_rsci_idat;
  output [31:0] crc32_dat_out_rsci_idat;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire dx_in_rsci_wen_comp;
  wire [35:0] dx_in_rsci_idat_mxwt;
  wire dy_in_rsci_wen_comp;
  wire [35:0] dy_in_rsci_idat_mxwt;
  wire pix_in_rsci_wen_comp;
  wire [31:0] pix_in_rsci_idat_mxwt;
  wire dat_out_rsci_wen_comp;
  reg dat_out_rsci_idat_33;
  reg dat_out_rsci_idat_32;
  reg [7:0] dat_out_rsci_idat_31_24;
  reg [7:0] dat_out_rsci_idat_23_16;
  reg [7:0] dat_out_rsci_idat_15_8;
  reg [7:0] dat_out_rsci_idat_7_0;
  reg not_64;
  reg not_65;
  reg not_66;
  reg not_67;
  reg not_68;
  reg not_69;
  reg not_70;
  reg not_71;
  reg not_72;
  reg not_73;
  reg not_74;
  reg not_75;
  reg not_76;
  reg not_77;
  reg not_78;
  reg not_79;
  reg not_80;
  reg not_81;
  reg not_82;
  reg not_83;
  reg not_84;
  reg not_85;
  reg not_86;
  reg not_87;
  reg not_88;
  reg not_89;
  reg not_90;
  reg not_91;
  reg not_92;
  reg not_93;
  reg not_94;
  reg not_95;
  reg not_96;
  reg not_97;
  reg not_98;
  reg not_99;
  reg not_100;
  reg not_101;
  reg not_102;
  reg not_103;
  reg not_104;
  reg not_105;
  reg not_106;
  reg not_107;
  reg not_108;
  reg not_109;
  reg not_110;
  reg not_111;
  reg not_112;
  reg not_113;
  reg not_114;
  reg not_115;
  reg not_116;
  reg not_117;
  reg not_118;
  reg not_119;
  reg not_120;
  reg not_121;
  reg not_122;
  reg not_123;
  reg not_124;
  reg not_125;
  reg not_126;
  reg not_127;
  wire [2:0] fsm_output;
  wire MROW_equal_tmp;
  wire and_dcpl_7;
  wire and_dcpl_9;
  wire or_tmp_2;
  wire [8:0] MCOL_for_abs_sum_clip_asn_sat_1_sva_1;
  wire [9:0] nl_MCOL_for_abs_sum_clip_asn_sat_1_sva_1;
  wire [8:0] MCOL_for_abs_sum_clip_asn_sat_2_sva_1;
  wire [9:0] nl_MCOL_for_abs_sum_clip_asn_sat_2_sva_1;
  wire [8:0] MCOL_for_abs_sum_clip_asn_sat_3_sva_1;
  wire [9:0] nl_MCOL_for_abs_sum_clip_asn_sat_3_sva_1;
  wire [8:0] MCOL_for_abs_sum_clip_asn_sat_sva_1;
  wire [9:0] nl_MCOL_for_abs_sum_clip_asn_sat_sva_1;
  reg MROW_stage_0;
  reg reg_pix_in_rsci_oswt_cse;
  wire MCOL_and_cse;
  wire MCOL_and_4_cse;
  reg reg_crc32_dat_out_triosy_obj_iswt0_cse;
  reg reg_dat_out_rsci_iswt0_cse;
  wire and_307_cse;
  wire MCOL_unequal_itm;
  wire [8:0] z_out;
  wire [9:0] nl_z_out;
  reg [8:0] MROW_y_sva;
  reg [7:0] MCOL_x_9_2_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_28_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_31_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_31_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_9_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_21_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_24_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_25_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_27_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_crc_tmp_30_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_28_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_31_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_31_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_9_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_21_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_24_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_25_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_27_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_sva;
  reg EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_30_sva;
  wire [7:0] magn_out_7_0_lpi_2_dfm_mx0w1;
  wire [7:0] magn_out_15_8_lpi_2_dfm_mx0w1;
  wire [7:0] magn_out_23_16_lpi_2_dfm_mx0w1;
  wire [7:0] magn_out_31_24_lpi_2_dfm_mx0w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva_1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_9_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_30_sva_mx1w0;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_27_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_sva_mx1w0;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva_mx1w0;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_25_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_24_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_21_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_31_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_28_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_31_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva_mx1w0;
  wire EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva_1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_9_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_30_sva_mx1w0;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_27_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_sva_mx1w0;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva_mx1w0;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_25_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_24_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_21_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_31_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_28_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_31_sva_mx1w1;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva_mx1w0;
  wire [7:0] magn_out_7_0_lpi_2_dfm_mx0;
  wire [7:0] magn_out_15_8_lpi_2_dfm_mx0;
  wire [7:0] magn_out_23_16_lpi_2_dfm_mx0;
  wire [7:0] magn_out_31_24_lpi_2_dfm_mx0;
  wire [8:0] operator_11_true_acc_psp_sva_1;
  wire [9:0] nl_operator_11_true_acc_psp_sva_1;
  wire xor_cse;
  wire xor_cse_3;
  wire xor_cse_6;
  wire xor_cse_9;
  wire xor_cse_12;
  wire xor_cse_15;
  wire xor_cse_18;
  wire xor_cse_20;
  wire xor_cse_22;
  wire xor_cse_24;
  wire xor_cse_28;
  wire xor_cse_31;
  wire xor_cse_35;
  wire xor_cse_37;
  wire xor_cse_42;
  wire xor_cse_43;
  wire xor_cse_45;
  wire xor_cse_48;
  wire xor_cse_50;
  wire xor_cse_52;
  wire xor_cse_58;
  wire xor_cse_60;
  wire xor_cse_62;
  wire xor_cse_65;
  wire xor_cse_66;
  wire xor_cse_69;
  wire xor_cse_71;
  wire xor_cse_73;
  wire xor_cse_74;
  wire xor_cse_76;
  wire xor_cse_79;
  wire xor_cse_84;
  wire xor_cse_85;
  wire xor_cse_86;
  wire xor_cse_87;
  wire xor_cse_88;
  wire xor_cse_91;
  wire xor_cse_92;
  wire xor_cse_93;
  wire xor_cse_95;
  wire xor_cse_98;
  wire xor_cse_99;
  wire xor_cse_100;
  wire xor_cse_102;
  wire xor_cse_110;
  wire xor_cse_118;
  wire xor_cse_119;
  wire xor_cse_123;
  wire xor_cse_125;
  wire xor_cse_128;
  wire xor_cse_146;
  wire xor_cse_149;
  wire xor_cse_152;
  wire xor_cse_155;
  wire xor_cse_158;
  wire xor_cse_161;
  wire xor_cse_164;
  wire xor_cse_166;
  wire xor_cse_168;
  wire xor_cse_170;
  wire xor_cse_174;
  wire xor_cse_177;
  wire xor_cse_181;
  wire xor_cse_183;
  wire xor_cse_188;
  wire xor_cse_189;
  wire xor_cse_191;
  wire xor_cse_194;
  wire xor_cse_196;
  wire xor_cse_198;
  wire xor_cse_204;
  wire xor_cse_206;
  wire xor_cse_208;
  wire xor_cse_211;
  wire xor_cse_212;
  wire xor_cse_215;
  wire xor_cse_217;
  wire xor_cse_219;
  wire xor_cse_220;
  wire xor_cse_222;
  wire xor_cse_225;
  wire xor_cse_230;
  wire xor_cse_231;
  wire xor_cse_232;
  wire xor_cse_233;
  wire xor_cse_234;
  wire xor_cse_237;
  wire xor_cse_238;
  wire xor_cse_239;
  wire xor_cse_241;
  wire xor_cse_244;
  wire xor_cse_245;
  wire xor_cse_246;
  wire xor_cse_248;
  wire xor_cse_256;
  wire xor_cse_264;
  wire xor_cse_265;
  wire xor_cse_269;
  wire xor_cse_271;
  wire xor_cse_274;
  wire nand_6_cse;
  wire nor_cse;
  wire nand_5_cse;
  wire and_373_itm;

  wire EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_mux1h_1_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_1_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_3_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_5_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_7_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_9_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_11_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_13_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_15_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_17_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_19_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_21_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_23_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_25_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_27_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_29_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_31_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_33_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_35_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_37_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_39_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_41_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_43_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_45_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_47_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_49_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_51_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_53_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_55_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_57_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_59_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_61_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_mux1h_1_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_1_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_3_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_5_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_7_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_9_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_11_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_13_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_15_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_17_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_19_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_21_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_23_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_25_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_27_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_29_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_31_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_33_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_35_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_37_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_39_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_41_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_43_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_45_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_47_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_49_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_51_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_53_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_55_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_57_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_59_nl;
  wire EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_61_nl;
  wire MCOL_if_1_MCOL_if_1_or_nl;
  wire[7:0] MCOL_for_1_ac_math_ac_abs_9_8_xabs_acc_nl;
  wire[8:0] nl_MCOL_for_1_ac_math_ac_abs_9_8_xabs_acc_nl;
  wire[7:0] MCOL_for_1_ac_math_ac_abs_9_8_xabs_xor_nl;
  wire[7:0] MCOL_for_1_ac_math_ac_abs_9_8_1_xabs_acc_nl;
  wire[8:0] nl_MCOL_for_1_ac_math_ac_abs_9_8_1_xabs_acc_nl;
  wire[7:0] MCOL_for_1_ac_math_ac_abs_9_8_1_xabs_xor_nl;
  wire[7:0] MCOL_for_2_ac_math_ac_abs_9_8_xabs_acc_nl;
  wire[8:0] nl_MCOL_for_2_ac_math_ac_abs_9_8_xabs_acc_nl;
  wire[7:0] MCOL_for_2_ac_math_ac_abs_9_8_xabs_xor_nl;
  wire[7:0] MCOL_for_2_ac_math_ac_abs_9_8_1_xabs_acc_nl;
  wire[8:0] nl_MCOL_for_2_ac_math_ac_abs_9_8_1_xabs_acc_nl;
  wire[7:0] MCOL_for_2_ac_math_ac_abs_9_8_1_xabs_xor_nl;
  wire[7:0] MCOL_for_3_ac_math_ac_abs_9_8_xabs_acc_nl;
  wire[8:0] nl_MCOL_for_3_ac_math_ac_abs_9_8_xabs_acc_nl;
  wire[7:0] MCOL_for_3_ac_math_ac_abs_9_8_xabs_xor_nl;
  wire[7:0] MCOL_for_3_ac_math_ac_abs_9_8_1_xabs_acc_nl;
  wire[8:0] nl_MCOL_for_3_ac_math_ac_abs_9_8_1_xabs_acc_nl;
  wire[7:0] MCOL_for_3_ac_math_ac_abs_9_8_1_xabs_xor_nl;
  wire[7:0] MCOL_for_4_ac_math_ac_abs_9_8_xabs_acc_nl;
  wire[8:0] nl_MCOL_for_4_ac_math_ac_abs_9_8_xabs_acc_nl;
  wire[7:0] MCOL_for_4_ac_math_ac_abs_9_8_xabs_xor_nl;
  wire[7:0] MCOL_for_4_ac_math_ac_abs_9_8_1_xabs_acc_nl;
  wire[8:0] nl_MCOL_for_4_ac_math_ac_abs_9_8_1_xabs_acc_nl;
  wire[7:0] MCOL_for_4_ac_math_ac_abs_9_8_1_xabs_xor_nl;
  wire[8:0] operator_9_false_acc_nl;
  wire[9:0] nl_operator_9_false_acc_nl;
  wire MROW_MROW_and_1_nl;
  wire[7:0] MROW_mux_2_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [33:0] nl_EdgeDetect_MagAng_run_dat_out_rsci_inst_dat_out_rsci_idat;
  assign nl_EdgeDetect_MagAng_run_dat_out_rsci_inst_dat_out_rsci_idat = {dat_out_rsci_idat_33
      , dat_out_rsci_idat_32 , dat_out_rsci_idat_31_24 , dat_out_rsci_idat_23_16
      , dat_out_rsci_idat_15_8 , dat_out_rsci_idat_7_0};
  wire  nl_EdgeDetect_MagAng_run_run_fsm_inst_MROW_C_0_tr0;
  assign nl_EdgeDetect_MagAng_run_run_fsm_inst_MROW_C_0_tr0 = ~ MROW_stage_0;
  EdgeDetect_MagAng_run_dx_in_rsci EdgeDetect_MagAng_run_dx_in_rsci_inst (
      .dx_in_rsc_dat(dx_in_rsc_dat),
      .dx_in_rsc_vld(dx_in_rsc_vld),
      .dx_in_rsc_rdy(dx_in_rsc_rdy),
      .run_wen(run_wen),
      .dx_in_rsci_oswt(reg_pix_in_rsci_oswt_cse),
      .dx_in_rsci_wen_comp(dx_in_rsci_wen_comp),
      .dx_in_rsci_idat_mxwt(dx_in_rsci_idat_mxwt)
    );
  EdgeDetect_MagAng_run_dy_in_rsci EdgeDetect_MagAng_run_dy_in_rsci_inst (
      .dy_in_rsc_dat(dy_in_rsc_dat),
      .dy_in_rsc_vld(dy_in_rsc_vld),
      .dy_in_rsc_rdy(dy_in_rsc_rdy),
      .run_wen(run_wen),
      .dy_in_rsci_oswt(reg_pix_in_rsci_oswt_cse),
      .dy_in_rsci_wen_comp(dy_in_rsci_wen_comp),
      .dy_in_rsci_idat_mxwt(dy_in_rsci_idat_mxwt)
    );
  EdgeDetect_MagAng_run_pix_in_rsci EdgeDetect_MagAng_run_pix_in_rsci_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .pix_in_rsc_dat(pix_in_rsc_dat),
      .pix_in_rsc_vld(pix_in_rsc_vld),
      .pix_in_rsc_rdy(pix_in_rsc_rdy),
      .run_wen(run_wen),
      .pix_in_rsci_oswt(reg_pix_in_rsci_oswt_cse),
      .pix_in_rsci_wen_comp(pix_in_rsci_wen_comp),
      .pix_in_rsci_idat_mxwt(pix_in_rsci_idat_mxwt)
    );
  EdgeDetect_MagAng_run_dat_out_rsci EdgeDetect_MagAng_run_dat_out_rsci_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .dat_out_rsc_dat(dat_out_rsc_dat),
      .dat_out_rsc_vld(dat_out_rsc_vld),
      .dat_out_rsc_rdy(dat_out_rsc_rdy),
      .run_wen(run_wen),
      .dat_out_rsci_oswt(reg_dat_out_rsci_iswt0_cse),
      .dat_out_rsci_wen_comp(dat_out_rsci_wen_comp),
      .dat_out_rsci_idat(nl_EdgeDetect_MagAng_run_dat_out_rsci_inst_dat_out_rsci_idat[33:0])
    );
  EdgeDetect_MagAng_run_crc32_pix_in_triosy_obj EdgeDetect_MagAng_run_crc32_pix_in_triosy_obj_inst
      (
      .crc32_pix_in_triosy_lz(crc32_pix_in_triosy_lz),
      .run_wten(run_wten),
      .crc32_pix_in_triosy_obj_iswt0(reg_crc32_dat_out_triosy_obj_iswt0_cse)
    );
  EdgeDetect_MagAng_run_crc32_dat_out_triosy_obj EdgeDetect_MagAng_run_crc32_dat_out_triosy_obj_inst
      (
      .crc32_dat_out_triosy_lz(crc32_dat_out_triosy_lz),
      .run_wten(run_wten),
      .crc32_dat_out_triosy_obj_iswt0(reg_crc32_dat_out_triosy_obj_iswt0_cse)
    );
  EdgeDetect_MagAng_run_staller EdgeDetect_MagAng_run_staller_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .dx_in_rsci_wen_comp(dx_in_rsci_wen_comp),
      .dy_in_rsci_wen_comp(dy_in_rsci_wen_comp),
      .pix_in_rsci_wen_comp(pix_in_rsci_wen_comp),
      .dat_out_rsci_wen_comp(dat_out_rsci_wen_comp)
    );
  EdgeDetect_MagAng_run_run_fsm EdgeDetect_MagAng_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .MROW_C_0_tr0(nl_EdgeDetect_MagAng_run_run_fsm_inst_MROW_C_0_tr0)
    );
  assign crc32_dat_out_rsci_idat = {not_64 , not_65 , not_66 , not_67 , not_68 ,
      not_69 , not_70 , not_71 , not_72 , not_73 , not_74 , not_75 , not_76 , not_77
      , not_78 , not_79 , not_80 , not_81 , not_82 , not_83 , not_84 , not_85 , not_86
      , not_87 , not_88 , not_89 , not_90 , not_91 , not_92 , not_93 , not_94 , not_95};
  assign crc32_pix_in_rsci_idat = {not_96 , not_97 , not_98 , not_99 , not_100 ,
      not_101 , not_102 , not_103 , not_104 , not_105 , not_106 , not_107 , not_108
      , not_109 , not_110 , not_111 , not_112 , not_113 , not_114 , not_115 , not_116
      , not_117 , not_118 , not_119 , not_120 , not_121 , not_122 , not_123 , not_124
      , not_125 , not_126 , not_127};
  assign nand_6_cse = ~(nor_cse & MROW_equal_tmp);
  assign nand_5_cse = ~(nand_6_cse & MROW_stage_0);
  assign MCOL_and_cse = run_wen & ((MROW_stage_0 & (~ sw_in) & (fsm_output[1])) |
      or_tmp_2);
  assign MCOL_and_4_cse = run_wen & MROW_stage_0 & (fsm_output[1]);
  assign nor_cse = ~(MCOL_unequal_itm | (operator_11_true_acc_psp_sva_1[8]));
  assign and_307_cse = run_wen & (~(MROW_stage_0 | (~ (fsm_output[1]))));
  assign magn_out_7_0_lpi_2_dfm_mx0w1 = MUX_v_8_2_2((MCOL_for_abs_sum_clip_asn_sat_1_sva_1[7:0]),
      8'b11111111, (MCOL_for_abs_sum_clip_asn_sat_1_sva_1[8]));
  assign magn_out_15_8_lpi_2_dfm_mx0w1 = MUX_v_8_2_2((MCOL_for_abs_sum_clip_asn_sat_2_sva_1[7:0]),
      8'b11111111, (MCOL_for_abs_sum_clip_asn_sat_2_sva_1[8]));
  assign magn_out_23_16_lpi_2_dfm_mx0w1 = MUX_v_8_2_2((MCOL_for_abs_sum_clip_asn_sat_3_sva_1[7:0]),
      8'b11111111, (MCOL_for_abs_sum_clip_asn_sat_3_sva_1[8]));
  assign magn_out_31_24_lpi_2_dfm_mx0w1 = MUX_v_8_2_2((MCOL_for_abs_sum_clip_asn_sat_sva_1[7:0]),
      8'b11111111, (MCOL_for_abs_sum_clip_asn_sat_sva_1[8]));
  assign MCOL_unequal_itm = MCOL_x_9_2_sva != (operator_11_true_acc_psp_sva_1[7:0]);
  assign magn_out_7_0_lpi_2_dfm_mx0 = MUX_v_8_2_2((pix_in_rsci_idat_mxwt[7:0]), magn_out_7_0_lpi_2_dfm_mx0w1,
      sw_in);
  assign magn_out_15_8_lpi_2_dfm_mx0 = MUX_v_8_2_2((pix_in_rsci_idat_mxwt[15:8]),
      magn_out_15_8_lpi_2_dfm_mx0w1, sw_in);
  assign magn_out_23_16_lpi_2_dfm_mx0 = MUX_v_8_2_2((pix_in_rsci_idat_mxwt[23:16]),
      magn_out_23_16_lpi_2_dfm_mx0w1, sw_in);
  assign magn_out_31_24_lpi_2_dfm_mx0 = MUX_v_8_2_2((pix_in_rsci_idat_mxwt[31:24]),
      magn_out_31_24_lpi_2_dfm_mx0w1, sw_in);
  assign MCOL_for_1_ac_math_ac_abs_9_8_xabs_xor_nl = (signext_8_1(dx_in_rsci_idat_mxwt[8]))
      ^ (dx_in_rsci_idat_mxwt[7:0]);
  assign nl_MCOL_for_1_ac_math_ac_abs_9_8_xabs_acc_nl = MCOL_for_1_ac_math_ac_abs_9_8_xabs_xor_nl
      + conv_u2u_1_8(dx_in_rsci_idat_mxwt[8]);
  assign MCOL_for_1_ac_math_ac_abs_9_8_xabs_acc_nl = nl_MCOL_for_1_ac_math_ac_abs_9_8_xabs_acc_nl[7:0];
  assign MCOL_for_1_ac_math_ac_abs_9_8_1_xabs_xor_nl = (signext_8_1(dy_in_rsci_idat_mxwt[8]))
      ^ (dy_in_rsci_idat_mxwt[7:0]);
  assign nl_MCOL_for_1_ac_math_ac_abs_9_8_1_xabs_acc_nl = MCOL_for_1_ac_math_ac_abs_9_8_1_xabs_xor_nl
      + conv_u2u_1_8(dy_in_rsci_idat_mxwt[8]);
  assign MCOL_for_1_ac_math_ac_abs_9_8_1_xabs_acc_nl = nl_MCOL_for_1_ac_math_ac_abs_9_8_1_xabs_acc_nl[7:0];
  assign nl_MCOL_for_abs_sum_clip_asn_sat_1_sva_1 = conv_u2u_8_9(MCOL_for_1_ac_math_ac_abs_9_8_xabs_acc_nl)
      + conv_u2u_8_9(MCOL_for_1_ac_math_ac_abs_9_8_1_xabs_acc_nl);
  assign MCOL_for_abs_sum_clip_asn_sat_1_sva_1 = nl_MCOL_for_abs_sum_clip_asn_sat_1_sva_1[8:0];
  assign MCOL_for_2_ac_math_ac_abs_9_8_xabs_xor_nl = (signext_8_1(dx_in_rsci_idat_mxwt[17]))
      ^ (dx_in_rsci_idat_mxwt[16:9]);
  assign nl_MCOL_for_2_ac_math_ac_abs_9_8_xabs_acc_nl = MCOL_for_2_ac_math_ac_abs_9_8_xabs_xor_nl
      + conv_u2u_1_8(dx_in_rsci_idat_mxwt[17]);
  assign MCOL_for_2_ac_math_ac_abs_9_8_xabs_acc_nl = nl_MCOL_for_2_ac_math_ac_abs_9_8_xabs_acc_nl[7:0];
  assign MCOL_for_2_ac_math_ac_abs_9_8_1_xabs_xor_nl = (signext_8_1(dy_in_rsci_idat_mxwt[17]))
      ^ (dy_in_rsci_idat_mxwt[16:9]);
  assign nl_MCOL_for_2_ac_math_ac_abs_9_8_1_xabs_acc_nl = MCOL_for_2_ac_math_ac_abs_9_8_1_xabs_xor_nl
      + conv_u2u_1_8(dy_in_rsci_idat_mxwt[17]);
  assign MCOL_for_2_ac_math_ac_abs_9_8_1_xabs_acc_nl = nl_MCOL_for_2_ac_math_ac_abs_9_8_1_xabs_acc_nl[7:0];
  assign nl_MCOL_for_abs_sum_clip_asn_sat_2_sva_1 = conv_u2u_8_9(MCOL_for_2_ac_math_ac_abs_9_8_xabs_acc_nl)
      + conv_u2u_8_9(MCOL_for_2_ac_math_ac_abs_9_8_1_xabs_acc_nl);
  assign MCOL_for_abs_sum_clip_asn_sat_2_sva_1 = nl_MCOL_for_abs_sum_clip_asn_sat_2_sva_1[8:0];
  assign MCOL_for_3_ac_math_ac_abs_9_8_xabs_xor_nl = (signext_8_1(dx_in_rsci_idat_mxwt[26]))
      ^ (dx_in_rsci_idat_mxwt[25:18]);
  assign nl_MCOL_for_3_ac_math_ac_abs_9_8_xabs_acc_nl = MCOL_for_3_ac_math_ac_abs_9_8_xabs_xor_nl
      + conv_u2u_1_8(dx_in_rsci_idat_mxwt[26]);
  assign MCOL_for_3_ac_math_ac_abs_9_8_xabs_acc_nl = nl_MCOL_for_3_ac_math_ac_abs_9_8_xabs_acc_nl[7:0];
  assign MCOL_for_3_ac_math_ac_abs_9_8_1_xabs_xor_nl = (signext_8_1(dy_in_rsci_idat_mxwt[26]))
      ^ (dy_in_rsci_idat_mxwt[25:18]);
  assign nl_MCOL_for_3_ac_math_ac_abs_9_8_1_xabs_acc_nl = MCOL_for_3_ac_math_ac_abs_9_8_1_xabs_xor_nl
      + conv_u2u_1_8(dy_in_rsci_idat_mxwt[26]);
  assign MCOL_for_3_ac_math_ac_abs_9_8_1_xabs_acc_nl = nl_MCOL_for_3_ac_math_ac_abs_9_8_1_xabs_acc_nl[7:0];
  assign nl_MCOL_for_abs_sum_clip_asn_sat_3_sva_1 = conv_u2u_8_9(MCOL_for_3_ac_math_ac_abs_9_8_xabs_acc_nl)
      + conv_u2u_8_9(MCOL_for_3_ac_math_ac_abs_9_8_1_xabs_acc_nl);
  assign MCOL_for_abs_sum_clip_asn_sat_3_sva_1 = nl_MCOL_for_abs_sum_clip_asn_sat_3_sva_1[8:0];
  assign MCOL_for_4_ac_math_ac_abs_9_8_xabs_xor_nl = (signext_8_1(dx_in_rsci_idat_mxwt[35]))
      ^ (dx_in_rsci_idat_mxwt[34:27]);
  assign nl_MCOL_for_4_ac_math_ac_abs_9_8_xabs_acc_nl = MCOL_for_4_ac_math_ac_abs_9_8_xabs_xor_nl
      + conv_u2u_1_8(dx_in_rsci_idat_mxwt[35]);
  assign MCOL_for_4_ac_math_ac_abs_9_8_xabs_acc_nl = nl_MCOL_for_4_ac_math_ac_abs_9_8_xabs_acc_nl[7:0];
  assign MCOL_for_4_ac_math_ac_abs_9_8_1_xabs_xor_nl = (signext_8_1(dy_in_rsci_idat_mxwt[35]))
      ^ (dy_in_rsci_idat_mxwt[34:27]);
  assign nl_MCOL_for_4_ac_math_ac_abs_9_8_1_xabs_acc_nl = MCOL_for_4_ac_math_ac_abs_9_8_1_xabs_xor_nl
      + conv_u2u_1_8(dy_in_rsci_idat_mxwt[35]);
  assign MCOL_for_4_ac_math_ac_abs_9_8_1_xabs_acc_nl = nl_MCOL_for_4_ac_math_ac_abs_9_8_1_xabs_acc_nl[7:0];
  assign nl_MCOL_for_abs_sum_clip_asn_sat_sva_1 = conv_u2u_8_9(MCOL_for_4_ac_math_ac_abs_9_8_xabs_acc_nl)
      + conv_u2u_8_9(MCOL_for_4_ac_math_ac_abs_9_8_1_xabs_acc_nl);
  assign MCOL_for_abs_sum_clip_asn_sat_sva_1 = nl_MCOL_for_abs_sum_clip_asn_sat_sva_1[8:0];
  assign nl_operator_9_false_acc_nl = heightIn + 9'b111111111;
  assign operator_9_false_acc_nl = nl_operator_9_false_acc_nl[8:0];
  assign MROW_equal_tmp = MROW_y_sva == operator_9_false_acc_nl;
  assign nl_operator_11_true_acc_psp_sva_1 = conv_u2s_8_9(widthIn[9:2]) + 9'b111111111;
  assign operator_11_true_acc_psp_sva_1 = nl_operator_11_true_acc_psp_sva_1[8:0];
  assign and_dcpl_7 = (~ nand_6_cse) & MROW_stage_0;
  assign and_dcpl_9 = nand_6_cse & MROW_stage_0;
  assign or_tmp_2 = MROW_stage_0 & sw_in & (fsm_output[1]);
  assign xor_cse = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[7])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_31_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[7]);
  assign xor_cse_3 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[0])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_25_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[6]);
  assign xor_cse_6 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[3])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[6]);
  assign xor_cse_9 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[7])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[1]);
  assign xor_cse_12 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[1])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[2]);
  assign xor_cse_15 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[5])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_21_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[3]);
  assign xor_cse_18 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_24_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[5]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva_1 = xor_cse ^ xor_cse_3
      ^ xor_cse_6 ^ xor_cse_9 ^ xor_cse_12 ^ xor_cse_15 ^ xor_cse_18;
  assign xor_cse_20 = xor_cse ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva
      ^ (magn_out_15_8_lpi_2_dfm_mx0[7]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_21_sva;
  assign xor_cse_22 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[5])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_9_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[0]);
  assign xor_cse_24 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[5])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[1]);
  assign xor_cse_28 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[4])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[4]);
  assign xor_cse_31 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_31_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[4])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[2]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_9_sva_mx1w1 = xor_cse_20 ^ (magn_out_23_16_lpi_2_dfm_mx0[3])
      ^ xor_cse_3 ^ xor_cse_22 ^ xor_cse_24 ^ xor_cse_28 ^ xor_cse_31;
  assign xor_cse_35 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[6])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[1]);
  assign xor_cse_37 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[6])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[2]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_30_sva_mx1w0 = xor_cse_20 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_25_sva
      ^ (magn_out_23_16_lpi_2_dfm_mx0[6]) ^ (magn_out_23_16_lpi_2_dfm_mx0[3]) ^ xor_cse_35
      ^ xor_cse_37 ^ xor_cse_28 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_27_sva
      ^ (magn_out_31_24_lpi_2_dfm_mx0[0]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[3]);
  assign xor_cse_43 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_28_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[4])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_31_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[4]);
  assign xor_cse_45 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[2])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[7]);
  assign xor_cse_42 = xor_cse_43 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva
      ^ (magn_out_31_24_lpi_2_dfm_mx0[1]) ^ xor_cse_45;
  assign xor_cse_48 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_30_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[3])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_21_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[3]);
  assign xor_cse_50 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[0])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[4]);
  assign xor_cse_52 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[5])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[0]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_27_sva_mx1w1 = xor_cse_42 ^ xor_cse
      ^ xor_cse_48 ^ xor_cse_50 ^ xor_cse_52 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_sva
      ^ (magn_out_15_8_lpi_2_dfm_mx0[3]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[1]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva
      ^ (magn_out_31_24_lpi_2_dfm_mx0[5]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[6]);
  assign xor_cse_58 = xor_cse ^ xor_cse_37 ^ xor_cse_35 ^ xor_cse_3;
  assign xor_cse_60 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_27_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[0])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[5]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_sva_mx1w0 = xor_cse_58 ^ xor_cse_60
      ^ xor_cse_24 ^ xor_cse_9 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva
      ^ (magn_out_23_16_lpi_2_dfm_mx0[7]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[5]);
  assign xor_cse_62 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[2])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[2]);
  assign xor_cse_65 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_30_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[3])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[3]);
  assign xor_cse_66 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[2])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_27_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[0]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva_mx1w1 = xor_cse ^ xor_cse_35
      ^ xor_cse_62 ^ xor_cse_43 ^ xor_cse_65 ^ xor_cse_66 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[2]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[3]) ^ xor_cse_18;
  assign xor_cse_69 = xor_cse_3 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[4]);
  assign xor_cse_71 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[0])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva;
  assign xor_cse_73 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[6])
      ^ (magn_out_31_24_lpi_2_dfm_mx0[6]);
  assign xor_cse_74 = (magn_out_15_8_lpi_2_dfm_mx0[6]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva
      ^ (magn_out_23_16_lpi_2_dfm_mx0[7]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva_mx1w0 = xor_cse_69 ^
      xor_cse_60 ^ xor_cse_43 ^ xor_cse_24 ^ xor_cse_71 ^ xor_cse_73 ^ xor_cse_74
      ^ xor_cse_18;
  assign xor_cse_76 = xor_cse_62 ^ xor_cse_45 ^ xor_cse_60;
  assign xor_cse_79 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[1])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[1]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_25_sva_mx1w1 = xor_cse_76 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva
      ^ (magn_out_23_16_lpi_2_dfm_mx0[4]) ^ xor_cse_35 ^ xor_cse_79 ^ xor_cse_65
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[1])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[6]);
  assign xor_cse_84 = EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[1])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_24_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[5]);
  assign xor_cse_85 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[7])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_28_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[4]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_24_sva_mx1w1 = xor_cse_76 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_9_sva
      ^ (magn_out_15_8_lpi_2_dfm_mx0[0]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva
      ^ (magn_out_23_16_lpi_2_dfm_mx0[0]) ^ xor_cse ^ xor_cse_6 ^ xor_cse_84 ^ xor_cse_85;
  assign xor_cse_86 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[3])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[6]);
  assign xor_cse_87 = (magn_out_31_24_lpi_2_dfm_mx0[6]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_9_sva;
  assign xor_cse_88 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_28_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[4])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[7]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva_mx1w1 = xor_cse_48 ^ xor_cse_84
      ^ xor_cse_86 ^ xor_cse_87 ^ xor_cse_88 ^ (magn_out_15_8_lpi_2_dfm_mx0[0]) ^
      (magn_out_23_16_lpi_2_dfm_mx0[4]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_31_sva
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[0])
      ^ (magn_out_31_24_lpi_2_dfm_mx0[7]);
  assign xor_cse_91 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[2])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[2]);
  assign xor_cse_92 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[7])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[5]);
  assign xor_cse_93 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[5])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_25_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[6]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva_mx1w1 = xor_cse_48 ^
      xor_cse_91 ^ xor_cse_87 ^ xor_cse_92 ^ xor_cse_93 ^ (magn_out_15_8_lpi_2_dfm_mx0[0])
      ^ (magn_out_23_16_lpi_2_dfm_mx0[4]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva
      ^ (magn_out_23_16_lpi_2_dfm_mx0[2]);
  assign xor_cse_95 = xor_cse_43 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva
      ^ (magn_out_23_16_lpi_2_dfm_mx0[2]);
  assign xor_cse_98 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[7])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[5]);
  assign xor_cse_99 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[3])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[1]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_21_sva_mx1w1 = xor_cse_95 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva
      ^ (magn_out_31_24_lpi_2_dfm_mx0[5]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_31_sva
      ^ (magn_out_31_24_lpi_2_dfm_mx0[7]) ^ xor_cse_3 ^ xor_cse_91 ^ xor_cse_98 ^
      xor_cse_99;
  assign xor_cse_100 = xor_cse_3 ^ xor_cse_6 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_28_sva
      ^ (magn_out_31_24_lpi_2_dfm_mx0[4]);
  assign xor_cse_102 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[4])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[3]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva_mx1w1 = xor_cse_100 ^ xor_cse
      ^ xor_cse_102 ^ xor_cse_48 ^ xor_cse_98 ^ xor_cse_71 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva
      ^ (magn_out_23_16_lpi_2_dfm_mx0[1]) ^ (magn_out_15_8_lpi_2_dfm_mx0[6]) ^ (magn_out_31_24_lpi_2_dfm_mx0[6]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva_mx1w1 = xor_cse_100 ^
      EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[1])
      ^ xor_cse_22 ^ xor_cse_12 ^ xor_cse_66 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[4]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva
      ^ (magn_out_15_8_lpi_2_dfm_mx0[2]);
  assign xor_cse_110 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[4])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[1]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva_mx1w1 = xor_cse_58 ^ (magn_out_15_8_lpi_2_dfm_mx0[5])
      ^ (magn_out_31_24_lpi_2_dfm_mx0[5]) ^ xor_cse_62 ^ xor_cse_48 ^ xor_cse_110
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[0])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva;
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva_mx1w1 = xor_cse_95 ^
      xor_cse_6 ^ xor_cse_60 ^ xor_cse_35 ^ xor_cse_24 ^ xor_cse_84 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_sva
      ^ (magn_out_31_24_lpi_2_dfm_mx0[2]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva
      ^ (magn_out_15_8_lpi_2_dfm_mx0[7]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[0]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva_mx1w1 = xor_cse_42 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva
      ^ (magn_out_15_8_lpi_2_dfm_mx0[6]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva
      ^ (magn_out_23_16_lpi_2_dfm_mx0[1]) ^ xor_cse_60 ^ xor_cse_22 ^ xor_cse_50
      ^ xor_cse_65;
  assign xor_cse_119 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_27_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[0])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[7]);
  assign xor_cse_118 = xor_cse_102 ^ xor_cse_62 ^ xor_cse_119;
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva_mx1w1 = xor_cse_118
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[0])
      ^ xor_cse_48 ^ xor_cse_9 ^ xor_cse_88 ^ xor_cse_93;
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva_mx1w1 = xor_cse ^ xor_cse_45
      ^ xor_cse_62 ^ xor_cse_48 ^ xor_cse_37 ^ xor_cse_79 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_31_sva
      ^ (magn_out_15_8_lpi_2_dfm_mx0[4]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[5]);
  assign xor_cse_123 = (magn_out_15_8_lpi_2_dfm_mx0[0]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_9_sva
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[2]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_31_sva_mx1w1 = xor_cse_3 ^
      xor_cse_35 ^ xor_cse_102 ^ xor_cse_24 ^ xor_cse_79 ^ xor_cse_123 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[6]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva
      ^ (magn_out_23_16_lpi_2_dfm_mx0[2]);
  assign xor_cse_125 = xor_cse_22 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva
      ^ (magn_out_31_24_lpi_2_dfm_mx0[1]);
  assign xor_cse_128 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[2])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_24_sva ^ (magn_out_23_16_lpi_2_dfm_mx0[5]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_sva_mx1w1 = xor_cse_125 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva
      ^ (magn_out_23_16_lpi_2_dfm_mx0[0]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[0]) ^ xor_cse_60 ^ xor_cse_99 ^ xor_cse_128 ^
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva ^ (magn_out_7_0_lpi_2_dfm_mx0[7])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_31_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[4]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva_mx1w1 = xor_cse_45 ^
      xor_cse_102 ^ xor_cse_50 ^ xor_cse_119 ^ xor_cse_85 ^ EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva
      ^ (magn_out_15_8_lpi_2_dfm_mx0[1]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[6]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_sva_mx1w1 = EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva
      ^ xor_cse_6 ^ xor_cse_22 ^ xor_cse_48 ^ xor_cse_9 ^ xor_cse_74 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_25_sva
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[2])
      ^ (magn_out_23_16_lpi_2_dfm_mx0[6]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva_mx1w1 = xor_cse_69 ^
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva ^ (magn_out_15_8_lpi_2_dfm_mx0[5])
      ^ xor_cse_37 ^ xor_cse_84 ^ xor_cse_91 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[7]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[5]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva_mx1w1 = xor_cse_45 ^
      xor_cse_22 ^ xor_cse_84 ^ xor_cse_119 ^ xor_cse_99 ^ xor_cse_110 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_30_sva
      ^ (magn_out_31_24_lpi_2_dfm_mx0[3]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_28_sva_mx1w1 = xor_cse_3 ^ xor_cse_45
      ^ xor_cse_6 ^ xor_cse_50 ^ xor_cse_110 ^ xor_cse_123 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva
      ^ (magn_out_7_0_lpi_2_dfm_mx0[7]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva_mx1w1 = xor_cse_3 ^ xor_cse_35
      ^ xor_cse_102 ^ xor_cse_37 ^ xor_cse_98 ^ xor_cse_31 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva
      ^ (magn_out_23_16_lpi_2_dfm_mx0[0]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_31_sva
      ^ (magn_out_31_24_lpi_2_dfm_mx0[7]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva_mx1w1 = xor_cse_60 ^
      xor_cse_102 ^ xor_cse_24 ^ xor_cse_9 ^ xor_cse_86 ^ xor_cse_128 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva
      ^ (magn_out_31_24_lpi_2_dfm_mx0[6]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva_mx1w1 = xor_cse_45 ^
      xor_cse_43 ^ xor_cse_50 ^ xor_cse_86 ^ xor_cse_52 ^ EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva
      ^ (magn_out_15_8_lpi_2_dfm_mx0[1]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva
      ^ (magn_out_15_8_lpi_2_dfm_mx0[2]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva
      ^ (magn_out_31_24_lpi_2_dfm_mx0[5]);
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva_mx1w1 = xor_cse_125 ^ xor_cse
      ^ xor_cse_6 ^ xor_cse_43 ^ xor_cse_84 ^ xor_cse_52 ^ xor_cse_65;
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_31_sva_mx1w1 = xor_cse_118 ^
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_30_sva ^ (magn_out_31_24_lpi_2_dfm_mx0[3])
      ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva
      ^ (magn_out_23_16_lpi_2_dfm_mx0[4]) ^ xor_cse_22 ^ xor_cse_31 ^ xor_cse_73;
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva_mx1w0 = xor_cse_6 ^ xor_cse_102
      ^ xor_cse_62 ^ xor_cse_79 ^ xor_cse_92 ^ xor_cse_15 ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva
      ^ (magn_out_31_24_lpi_2_dfm_mx0[1]) ^ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva
      ^ (magn_out_23_16_lpi_2_dfm_mx0[7]);
  assign xor_cse_146 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva ^ (pix_in_rsci_idat_mxwt[7])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_31_sva ^ (pix_in_rsci_idat_mxwt[31]);
  assign xor_cse_149 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva ^ (pix_in_rsci_idat_mxwt[0])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_25_sva ^ (pix_in_rsci_idat_mxwt[22]);
  assign xor_cse_152 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva ^ (pix_in_rsci_idat_mxwt[3])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva ^ (pix_in_rsci_idat_mxwt[6]);
  assign xor_cse_155 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva ^ (pix_in_rsci_idat_mxwt[15])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_sva ^ (pix_in_rsci_idat_mxwt[1]);
  assign xor_cse_158 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva ^ (pix_in_rsci_idat_mxwt[25])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva ^ (pix_in_rsci_idat_mxwt[2]);
  assign xor_cse_161 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva ^ (pix_in_rsci_idat_mxwt[5])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_21_sva ^ (pix_in_rsci_idat_mxwt[19]);
  assign xor_cse_164 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_24_sva ^ (pix_in_rsci_idat_mxwt[21]);
  assign EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva_1 = xor_cse_146 ^ xor_cse_149
      ^ xor_cse_152 ^ xor_cse_155 ^ xor_cse_158 ^ xor_cse_161 ^ xor_cse_164;
  assign xor_cse_166 = xor_cse_146 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva
      ^ (pix_in_rsci_idat_mxwt[15]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_21_sva;
  assign xor_cse_168 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva ^ (pix_in_rsci_idat_mxwt[5])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_9_sva ^ (pix_in_rsci_idat_mxwt[8]);
  assign xor_cse_170 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva ^ (pix_in_rsci_idat_mxwt[13])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva ^ (pix_in_rsci_idat_mxwt[17]);
  assign xor_cse_174 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva ^ (pix_in_rsci_idat_mxwt[4])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva ^ (pix_in_rsci_idat_mxwt[20]);
  assign xor_cse_177 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_31_sva ^ (pix_in_rsci_idat_mxwt[12])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva ^ (pix_in_rsci_idat_mxwt[2]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_9_sva_mx1w1 = xor_cse_166 ^ (pix_in_rsci_idat_mxwt[19])
      ^ xor_cse_149 ^ xor_cse_168 ^ xor_cse_170 ^ xor_cse_174 ^ xor_cse_177;
  assign xor_cse_181 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva ^ (pix_in_rsci_idat_mxwt[30])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva ^ (pix_in_rsci_idat_mxwt[25]);
  assign xor_cse_183 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva ^ (pix_in_rsci_idat_mxwt[14])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva ^ (pix_in_rsci_idat_mxwt[18]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_30_sva_mx1w0 = xor_cse_166 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_25_sva
      ^ (pix_in_rsci_idat_mxwt[22]) ^ (pix_in_rsci_idat_mxwt[19]) ^ xor_cse_181 ^
      xor_cse_183 ^ xor_cse_174 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_27_sva
      ^ (pix_in_rsci_idat_mxwt[24]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva
      ^ (pix_in_rsci_idat_mxwt[3]);
  assign xor_cse_189 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_28_sva ^ (pix_in_rsci_idat_mxwt[28])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_31_sva ^ (pix_in_rsci_idat_mxwt[12]);
  assign xor_cse_191 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva ^ (pix_in_rsci_idat_mxwt[2])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva ^ (pix_in_rsci_idat_mxwt[23]);
  assign xor_cse_188 = xor_cse_189 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva
      ^ (pix_in_rsci_idat_mxwt[25]) ^ xor_cse_191;
  assign xor_cse_194 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_30_sva ^ (pix_in_rsci_idat_mxwt[27])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_21_sva ^ (pix_in_rsci_idat_mxwt[19]);
  assign xor_cse_196 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva ^ (pix_in_rsci_idat_mxwt[16])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva ^ (pix_in_rsci_idat_mxwt[20]);
  assign xor_cse_198 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva ^ (pix_in_rsci_idat_mxwt[13])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva ^ (pix_in_rsci_idat_mxwt[0]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_27_sva_mx1w1 = xor_cse_188 ^ xor_cse_146
      ^ xor_cse_194 ^ xor_cse_196 ^ xor_cse_198 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_sva
      ^ (pix_in_rsci_idat_mxwt[11]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_sva
      ^ (pix_in_rsci_idat_mxwt[1]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva
      ^ (pix_in_rsci_idat_mxwt[29]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva
      ^ (pix_in_rsci_idat_mxwt[6]);
  assign xor_cse_204 = xor_cse_146 ^ xor_cse_183 ^ xor_cse_181 ^ xor_cse_149;
  assign xor_cse_206 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_27_sva ^ (pix_in_rsci_idat_mxwt[24])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva ^ (pix_in_rsci_idat_mxwt[29]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_sva_mx1w0 = xor_cse_204 ^ xor_cse_206
      ^ xor_cse_170 ^ xor_cse_155 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva
      ^ (pix_in_rsci_idat_mxwt[23]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva
      ^ (pix_in_rsci_idat_mxwt[5]);
  assign xor_cse_208 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_sva ^ (pix_in_rsci_idat_mxwt[26])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva ^ (pix_in_rsci_idat_mxwt[10]);
  assign xor_cse_211 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_30_sva ^ (pix_in_rsci_idat_mxwt[27])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_sva ^ (pix_in_rsci_idat_mxwt[11]);
  assign xor_cse_212 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva ^ (pix_in_rsci_idat_mxwt[18])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_27_sva ^ (pix_in_rsci_idat_mxwt[24]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva_mx1w1 = xor_cse_146 ^ xor_cse_181
      ^ xor_cse_208 ^ xor_cse_189 ^ xor_cse_211 ^ xor_cse_212 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva
      ^ (pix_in_rsci_idat_mxwt[2]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva
      ^ (pix_in_rsci_idat_mxwt[3]) ^ xor_cse_164;
  assign xor_cse_215 = xor_cse_149 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva
      ^ (pix_in_rsci_idat_mxwt[4]);
  assign xor_cse_217 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva ^ (pix_in_rsci_idat_mxwt[16])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva;
  assign xor_cse_219 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva ^ (pix_in_rsci_idat_mxwt[6])
      ^ (pix_in_rsci_idat_mxwt[30]);
  assign xor_cse_220 = (pix_in_rsci_idat_mxwt[14]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva
      ^ (pix_in_rsci_idat_mxwt[23]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva_mx1w0 = xor_cse_215 ^
      xor_cse_206 ^ xor_cse_189 ^ xor_cse_170 ^ xor_cse_217 ^ xor_cse_219 ^ xor_cse_220
      ^ xor_cse_164;
  assign xor_cse_222 = xor_cse_208 ^ xor_cse_191 ^ xor_cse_206;
  assign xor_cse_225 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_sva ^ (pix_in_rsci_idat_mxwt[1])
      ^ EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva ^ (pix_in_rsci_idat_mxwt[9]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_25_sva_mx1w1 = xor_cse_222 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva
      ^ (pix_in_rsci_idat_mxwt[20]) ^ xor_cse_181 ^ xor_cse_225 ^ xor_cse_211 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva
      ^ (pix_in_rsci_idat_mxwt[17]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva
      ^ (pix_in_rsci_idat_mxwt[6]);
  assign xor_cse_230 = EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva ^ (pix_in_rsci_idat_mxwt[9])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_24_sva ^ (pix_in_rsci_idat_mxwt[21]);
  assign xor_cse_231 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva ^ (pix_in_rsci_idat_mxwt[15])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_28_sva ^ (pix_in_rsci_idat_mxwt[28]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_24_sva_mx1w1 = xor_cse_222 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_9_sva
      ^ (pix_in_rsci_idat_mxwt[8]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva
      ^ (pix_in_rsci_idat_mxwt[16]) ^ xor_cse_146 ^ xor_cse_152 ^ xor_cse_230 ^ xor_cse_231;
  assign xor_cse_232 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva ^ (pix_in_rsci_idat_mxwt[3])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva ^ (pix_in_rsci_idat_mxwt[14]);
  assign xor_cse_233 = (pix_in_rsci_idat_mxwt[30]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_9_sva;
  assign xor_cse_234 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_28_sva ^ (pix_in_rsci_idat_mxwt[28])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva ^ (pix_in_rsci_idat_mxwt[23]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva_mx1w1 = xor_cse_194 ^ xor_cse_230
      ^ xor_cse_232 ^ xor_cse_233 ^ xor_cse_234 ^ (pix_in_rsci_idat_mxwt[8]) ^ (pix_in_rsci_idat_mxwt[20])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_31_sva ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva
      ^ (pix_in_rsci_idat_mxwt[0]) ^ (pix_in_rsci_idat_mxwt[31]);
  assign xor_cse_237 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva ^ (pix_in_rsci_idat_mxwt[2])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_sva ^ (pix_in_rsci_idat_mxwt[26]);
  assign xor_cse_238 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva ^ (pix_in_rsci_idat_mxwt[7])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva ^ (pix_in_rsci_idat_mxwt[29]);
  assign xor_cse_239 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva ^ (pix_in_rsci_idat_mxwt[13])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_25_sva ^ (pix_in_rsci_idat_mxwt[22]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva_mx1w1 = xor_cse_194 ^
      xor_cse_237 ^ xor_cse_233 ^ xor_cse_238 ^ xor_cse_239 ^ (pix_in_rsci_idat_mxwt[8])
      ^ (pix_in_rsci_idat_mxwt[20]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva
      ^ (pix_in_rsci_idat_mxwt[18]);
  assign xor_cse_241 = xor_cse_189 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva
      ^ (pix_in_rsci_idat_mxwt[18]);
  assign xor_cse_244 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva ^ (pix_in_rsci_idat_mxwt[15])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva ^ (pix_in_rsci_idat_mxwt[5]);
  assign xor_cse_245 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva ^ (pix_in_rsci_idat_mxwt[3])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva ^ (pix_in_rsci_idat_mxwt[17]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_21_sva_mx1w1 = xor_cse_241 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva
      ^ (pix_in_rsci_idat_mxwt[29]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_31_sva
      ^ (pix_in_rsci_idat_mxwt[31]) ^ xor_cse_149 ^ xor_cse_237 ^ xor_cse_244 ^ xor_cse_245;
  assign xor_cse_246 = xor_cse_149 ^ xor_cse_152 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_28_sva
      ^ (pix_in_rsci_idat_mxwt[28]);
  assign xor_cse_248 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva ^ (pix_in_rsci_idat_mxwt[4])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_sva ^ (pix_in_rsci_idat_mxwt[11]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva_mx1w1 = xor_cse_246 ^ xor_cse_146
      ^ xor_cse_248 ^ xor_cse_194 ^ xor_cse_244 ^ xor_cse_217 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva
      ^ (pix_in_rsci_idat_mxwt[17]) ^ (pix_in_rsci_idat_mxwt[14]) ^ (pix_in_rsci_idat_mxwt[30]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva_mx1w1 = xor_cse_246 ^ EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva
      ^ (pix_in_rsci_idat_mxwt[9]) ^ xor_cse_168 ^ xor_cse_158 ^ xor_cse_212 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva
      ^ (pix_in_rsci_idat_mxwt[4]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva
      ^ (pix_in_rsci_idat_mxwt[10]);
  assign xor_cse_256 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva ^ (pix_in_rsci_idat_mxwt[4])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_sva ^ (pix_in_rsci_idat_mxwt[1]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva_mx1w1 = xor_cse_204 ^ (pix_in_rsci_idat_mxwt[13])
      ^ (pix_in_rsci_idat_mxwt[29]) ^ xor_cse_208 ^ xor_cse_194 ^ xor_cse_256 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva
      ^ (pix_in_rsci_idat_mxwt[16]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva;
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva_mx1w1 = xor_cse_241 ^
      xor_cse_152 ^ xor_cse_206 ^ xor_cse_181 ^ xor_cse_170 ^ xor_cse_230 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_sva
      ^ (pix_in_rsci_idat_mxwt[26]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva
      ^ (pix_in_rsci_idat_mxwt[15]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva
      ^ (pix_in_rsci_idat_mxwt[0]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva_mx1w1 = xor_cse_188 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva
      ^ (pix_in_rsci_idat_mxwt[14]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva
      ^ (pix_in_rsci_idat_mxwt[17]) ^ xor_cse_206 ^ xor_cse_168 ^ xor_cse_196 ^ xor_cse_211;
  assign xor_cse_265 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_27_sva ^ (pix_in_rsci_idat_mxwt[24])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva ^ (pix_in_rsci_idat_mxwt[7]);
  assign xor_cse_264 = xor_cse_248 ^ xor_cse_208 ^ xor_cse_265;
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva_mx1w1 = xor_cse_264 ^
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva ^ (pix_in_rsci_idat_mxwt[16])
      ^ xor_cse_194 ^ xor_cse_155 ^ xor_cse_234 ^ xor_cse_239;
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva_mx1w1 = xor_cse_146 ^ xor_cse_191
      ^ xor_cse_208 ^ xor_cse_194 ^ xor_cse_183 ^ xor_cse_225 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_31_sva
      ^ (pix_in_rsci_idat_mxwt[12]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva
      ^ (pix_in_rsci_idat_mxwt[5]);
  assign xor_cse_269 = (pix_in_rsci_idat_mxwt[8]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_9_sva
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_sva ^ (pix_in_rsci_idat_mxwt[26]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_31_sva_mx1w1 = xor_cse_149 ^
      xor_cse_181 ^ xor_cse_248 ^ xor_cse_170 ^ xor_cse_225 ^ xor_cse_269 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva
      ^ (pix_in_rsci_idat_mxwt[6]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva
      ^ (pix_in_rsci_idat_mxwt[18]);
  assign xor_cse_271 = xor_cse_168 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva
      ^ (pix_in_rsci_idat_mxwt[25]);
  assign xor_cse_274 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva ^ (pix_in_rsci_idat_mxwt[10])
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_24_sva ^ (pix_in_rsci_idat_mxwt[21]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_sva_mx1w1 = xor_cse_271 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva
      ^ (pix_in_rsci_idat_mxwt[16]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva
      ^ (pix_in_rsci_idat_mxwt[0]) ^ xor_cse_206 ^ xor_cse_245 ^ xor_cse_274 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva
      ^ (pix_in_rsci_idat_mxwt[7]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_31_sva
      ^ (pix_in_rsci_idat_mxwt[12]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva_mx1w1 = xor_cse_191 ^
      xor_cse_248 ^ xor_cse_196 ^ xor_cse_265 ^ xor_cse_231 ^ EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva
      ^ (pix_in_rsci_idat_mxwt[9]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva
      ^ (pix_in_rsci_idat_mxwt[6]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_sva_mx1w1 = EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva
      ^ xor_cse_152 ^ xor_cse_168 ^ xor_cse_194 ^ xor_cse_155 ^ xor_cse_220 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_25_sva
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva ^ (pix_in_rsci_idat_mxwt[10])
      ^ (pix_in_rsci_idat_mxwt[22]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva_mx1w1 = xor_cse_215 ^
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva ^ (pix_in_rsci_idat_mxwt[13])
      ^ xor_cse_183 ^ xor_cse_230 ^ xor_cse_237 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva
      ^ (pix_in_rsci_idat_mxwt[7]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva
      ^ (pix_in_rsci_idat_mxwt[5]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva_mx1w1 = xor_cse_191 ^ xor_cse_168
      ^ xor_cse_230 ^ xor_cse_265 ^ xor_cse_245 ^ xor_cse_256 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_30_sva
      ^ (pix_in_rsci_idat_mxwt[27]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_28_sva_mx1w1 = xor_cse_149 ^ xor_cse_191
      ^ xor_cse_152 ^ xor_cse_196 ^ xor_cse_256 ^ xor_cse_269 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva
      ^ (pix_in_rsci_idat_mxwt[7]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva_mx1w1 = xor_cse_149 ^ xor_cse_181
      ^ xor_cse_248 ^ xor_cse_183 ^ xor_cse_244 ^ xor_cse_177 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva
      ^ (pix_in_rsci_idat_mxwt[16]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_31_sva
      ^ (pix_in_rsci_idat_mxwt[31]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva_mx1w1 = xor_cse_206 ^ xor_cse_248
      ^ xor_cse_170 ^ xor_cse_155 ^ xor_cse_232 ^ xor_cse_274 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva
      ^ (pix_in_rsci_idat_mxwt[30]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva_mx1w1 = xor_cse_191 ^ xor_cse_189
      ^ xor_cse_196 ^ xor_cse_232 ^ xor_cse_198 ^ EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva
      ^ (pix_in_rsci_idat_mxwt[9]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva
      ^ (pix_in_rsci_idat_mxwt[10]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva
      ^ (pix_in_rsci_idat_mxwt[29]);
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva_mx1w1 = xor_cse_271 ^ xor_cse_146
      ^ xor_cse_152 ^ xor_cse_189 ^ xor_cse_230 ^ xor_cse_198 ^ xor_cse_211;
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_31_sva_mx1w1 = xor_cse_264 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_30_sva
      ^ (pix_in_rsci_idat_mxwt[27]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva
      ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva ^ (pix_in_rsci_idat_mxwt[20])
      ^ xor_cse_168 ^ xor_cse_177 ^ xor_cse_219;
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva_mx1w0 = xor_cse_152 ^ xor_cse_248
      ^ xor_cse_208 ^ xor_cse_225 ^ xor_cse_238 ^ xor_cse_161 ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva
      ^ (pix_in_rsci_idat_mxwt[25]) ^ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva
      ^ (pix_in_rsci_idat_mxwt[23]);
  assign and_373_itm = ((operator_11_true_acc_psp_sva_1[8]) | MCOL_unequal_itm) &
      (fsm_output[1]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_pix_in_rsci_oswt_cse <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_27_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_25_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_24_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_21_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_9_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_28_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_27_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_25_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_24_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_21_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_9_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_28_sva <= 1'b0;
      MROW_stage_0 <= 1'b0;
      reg_crc32_dat_out_triosy_obj_iswt0_cse <= 1'b0;
      reg_dat_out_rsci_iswt0_cse <= 1'b0;
    end
    else if ( rst ) begin
      reg_pix_in_rsci_oswt_cse <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_27_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_25_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_24_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_21_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_9_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_28_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_27_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_25_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_24_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_21_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_9_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_31_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva <= 1'b0;
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_28_sva <= 1'b0;
      MROW_stage_0 <= 1'b0;
      reg_crc32_dat_out_triosy_obj_iswt0_cse <= 1'b0;
      reg_dat_out_rsci_iswt0_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_pix_in_rsci_oswt_cse <= ~((nand_5_cse & (fsm_output[1])) | (fsm_output[2]));
      EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva <= EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_mux1h_1_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_30_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_1_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_3_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_5_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_27_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_7_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_9_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_25_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_11_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_24_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_13_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_15_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_17_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_21_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_19_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_21_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_23_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_25_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_27_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_29_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_31_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_31_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_33_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_35_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_37_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_39_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_41_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_9_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_43_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_45_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_47_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_49_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_51_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_31_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_53_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_55_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_57_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_59_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_28_sva <= EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_61_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva <= EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_mux1h_1_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_30_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_1_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_3_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_5_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_27_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_7_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_9_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_25_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_11_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_24_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_13_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_15_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_17_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_21_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_19_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_21_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_23_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_25_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_27_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_29_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_31_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_31_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_33_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_35_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_37_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_39_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_41_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_9_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_43_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_45_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_47_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_49_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_51_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_31_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_53_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_55_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_57_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_59_nl
          | (~ (fsm_output[1]));
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_28_sva <= EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_61_nl
          | (~ (fsm_output[1]));
      MROW_stage_0 <= ~(nand_5_cse & (fsm_output[1]));
      reg_crc32_dat_out_triosy_obj_iswt0_cse <= (~ MROW_stage_0) & (fsm_output[1]);
      reg_dat_out_rsci_iswt0_cse <= MROW_stage_0 & (fsm_output[1]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dat_out_rsci_idat_7_0 <= 8'b00000000;
      dat_out_rsci_idat_15_8 <= 8'b00000000;
      dat_out_rsci_idat_23_16 <= 8'b00000000;
      dat_out_rsci_idat_31_24 <= 8'b00000000;
    end
    else if ( rst ) begin
      dat_out_rsci_idat_7_0 <= 8'b00000000;
      dat_out_rsci_idat_15_8 <= 8'b00000000;
      dat_out_rsci_idat_23_16 <= 8'b00000000;
      dat_out_rsci_idat_31_24 <= 8'b00000000;
    end
    else if ( MCOL_and_cse ) begin
      dat_out_rsci_idat_7_0 <= MUX_v_8_2_2((pix_in_rsci_idat_mxwt[7:0]), magn_out_7_0_lpi_2_dfm_mx0w1,
          or_tmp_2);
      dat_out_rsci_idat_15_8 <= MUX_v_8_2_2((pix_in_rsci_idat_mxwt[15:8]), magn_out_15_8_lpi_2_dfm_mx0w1,
          or_tmp_2);
      dat_out_rsci_idat_23_16 <= MUX_v_8_2_2((pix_in_rsci_idat_mxwt[23:16]), magn_out_23_16_lpi_2_dfm_mx0w1,
          or_tmp_2);
      dat_out_rsci_idat_31_24 <= MUX_v_8_2_2((pix_in_rsci_idat_mxwt[31:24]), magn_out_31_24_lpi_2_dfm_mx0w1,
          or_tmp_2);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dat_out_rsci_idat_32 <= 1'b0;
      dat_out_rsci_idat_33 <= 1'b0;
    end
    else if ( rst ) begin
      dat_out_rsci_idat_32 <= 1'b0;
      dat_out_rsci_idat_33 <= 1'b0;
    end
    else if ( MCOL_and_4_cse ) begin
      dat_out_rsci_idat_32 <= ~((MROW_y_sva!=9'b000000000) | (MCOL_x_9_2_sva!=8'b00000000));
      dat_out_rsci_idat_33 <= nor_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      MROW_y_sva <= 9'b000000000;
    end
    else if ( rst ) begin
      MROW_y_sva <= 9'b000000000;
    end
    else if ( (~((~(nor_cse & MROW_stage_0)) & (fsm_output[1]))) & run_wen ) begin
      MROW_y_sva <= MUX_v_9_2_2(9'b000000000, z_out, (fsm_output[1]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      MCOL_x_9_2_sva <= 8'b00000000;
    end
    else if ( rst ) begin
      MCOL_x_9_2_sva <= 8'b00000000;
    end
    else if ( (MROW_stage_0 | (~ (fsm_output[1]))) & run_wen ) begin
      MCOL_x_9_2_sva <= (z_out[7:0]) & (signext_8_1(MCOL_if_1_MCOL_if_1_or_nl)) &
          (signext_8_1(fsm_output[1]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      not_95 <= 1'b0;
      not_94 <= 1'b0;
      not_93 <= 1'b0;
      not_92 <= 1'b0;
      not_91 <= 1'b0;
      not_90 <= 1'b0;
      not_89 <= 1'b0;
      not_88 <= 1'b0;
      not_87 <= 1'b0;
      not_86 <= 1'b0;
      not_85 <= 1'b0;
      not_84 <= 1'b0;
      not_83 <= 1'b0;
      not_82 <= 1'b0;
      not_81 <= 1'b0;
      not_80 <= 1'b0;
      not_79 <= 1'b0;
      not_78 <= 1'b0;
      not_77 <= 1'b0;
      not_76 <= 1'b0;
      not_75 <= 1'b0;
      not_74 <= 1'b0;
      not_73 <= 1'b0;
      not_72 <= 1'b0;
      not_71 <= 1'b0;
      not_70 <= 1'b0;
      not_69 <= 1'b0;
      not_68 <= 1'b0;
      not_67 <= 1'b0;
      not_66 <= 1'b0;
      not_65 <= 1'b0;
      not_64 <= 1'b0;
      not_127 <= 1'b0;
      not_126 <= 1'b0;
      not_125 <= 1'b0;
      not_124 <= 1'b0;
      not_123 <= 1'b0;
      not_122 <= 1'b0;
      not_121 <= 1'b0;
      not_120 <= 1'b0;
      not_119 <= 1'b0;
      not_118 <= 1'b0;
      not_117 <= 1'b0;
      not_116 <= 1'b0;
      not_115 <= 1'b0;
      not_114 <= 1'b0;
      not_113 <= 1'b0;
      not_112 <= 1'b0;
      not_111 <= 1'b0;
      not_110 <= 1'b0;
      not_109 <= 1'b0;
      not_108 <= 1'b0;
      not_107 <= 1'b0;
      not_106 <= 1'b0;
      not_105 <= 1'b0;
      not_104 <= 1'b0;
      not_103 <= 1'b0;
      not_102 <= 1'b0;
      not_101 <= 1'b0;
      not_100 <= 1'b0;
      not_99 <= 1'b0;
      not_98 <= 1'b0;
      not_97 <= 1'b0;
      not_96 <= 1'b0;
    end
    else if ( rst ) begin
      not_95 <= 1'b0;
      not_94 <= 1'b0;
      not_93 <= 1'b0;
      not_92 <= 1'b0;
      not_91 <= 1'b0;
      not_90 <= 1'b0;
      not_89 <= 1'b0;
      not_88 <= 1'b0;
      not_87 <= 1'b0;
      not_86 <= 1'b0;
      not_85 <= 1'b0;
      not_84 <= 1'b0;
      not_83 <= 1'b0;
      not_82 <= 1'b0;
      not_81 <= 1'b0;
      not_80 <= 1'b0;
      not_79 <= 1'b0;
      not_78 <= 1'b0;
      not_77 <= 1'b0;
      not_76 <= 1'b0;
      not_75 <= 1'b0;
      not_74 <= 1'b0;
      not_73 <= 1'b0;
      not_72 <= 1'b0;
      not_71 <= 1'b0;
      not_70 <= 1'b0;
      not_69 <= 1'b0;
      not_68 <= 1'b0;
      not_67 <= 1'b0;
      not_66 <= 1'b0;
      not_65 <= 1'b0;
      not_64 <= 1'b0;
      not_127 <= 1'b0;
      not_126 <= 1'b0;
      not_125 <= 1'b0;
      not_124 <= 1'b0;
      not_123 <= 1'b0;
      not_122 <= 1'b0;
      not_121 <= 1'b0;
      not_120 <= 1'b0;
      not_119 <= 1'b0;
      not_118 <= 1'b0;
      not_117 <= 1'b0;
      not_116 <= 1'b0;
      not_115 <= 1'b0;
      not_114 <= 1'b0;
      not_113 <= 1'b0;
      not_112 <= 1'b0;
      not_111 <= 1'b0;
      not_110 <= 1'b0;
      not_109 <= 1'b0;
      not_108 <= 1'b0;
      not_107 <= 1'b0;
      not_106 <= 1'b0;
      not_105 <= 1'b0;
      not_104 <= 1'b0;
      not_103 <= 1'b0;
      not_102 <= 1'b0;
      not_101 <= 1'b0;
      not_100 <= 1'b0;
      not_99 <= 1'b0;
      not_98 <= 1'b0;
      not_97 <= 1'b0;
      not_96 <= 1'b0;
    end
    else if ( and_307_cse ) begin
      not_95 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_28_sva;
      not_94 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva;
      not_93 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva;
      not_92 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva;
      not_91 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_31_sva;
      not_90 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva;
      not_89 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva;
      not_88 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva;
      not_87 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva;
      not_86 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_9_sva;
      not_85 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva;
      not_84 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_sva;
      not_83 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva;
      not_82 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_sva;
      not_81 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_31_sva;
      not_80 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva;
      not_79 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva;
      not_78 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva;
      not_77 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva;
      not_76 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva;
      not_75 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva;
      not_74 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_21_sva;
      not_73 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva;
      not_72 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva;
      not_71 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_24_sva;
      not_70 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_25_sva;
      not_69 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva;
      not_68 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_27_sva;
      not_67 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva;
      not_66 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_sva;
      not_65 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_30_sva;
      not_64 <= ~ EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva;
      not_127 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_28_sva;
      not_126 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva;
      not_125 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva;
      not_124 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva;
      not_123 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_31_sva;
      not_122 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva;
      not_121 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva;
      not_120 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva;
      not_119 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva;
      not_118 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_9_sva;
      not_117 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva;
      not_116 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_sva;
      not_115 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva;
      not_114 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_sva;
      not_113 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_31_sva;
      not_112 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva;
      not_111 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva;
      not_110 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva;
      not_109 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva;
      not_108 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva;
      not_107 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva;
      not_106 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_21_sva;
      not_105 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva;
      not_104 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva;
      not_103 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_24_sva;
      not_102 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_25_sva;
      not_101 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva;
      not_100 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_27_sva;
      not_99 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva;
      not_98 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_sva;
      not_97 <= ~ EdgeDetect_MagAng_calc_crc32_32_crc_tmp_30_sva;
      not_96 <= ~ EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva;
    end
  end
  assign EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_mux1h_1_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva_1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_9_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_1_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_30_sva_mx1w0,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_27_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_30_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_3_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_sva_mx1w0,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_5_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva_mx1w0,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_25_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_7_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_27_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_24_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_27_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_9_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_26_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_11_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_25_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_25_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_13_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_24_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_21_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_24_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_15_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_17_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_23_31_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_19_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_21_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_21_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_21_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_20_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_23_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_25_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_19_31_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_27_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_29_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_31_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_17_31_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_31_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_33_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_31_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_15_31_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_35_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_37_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_14_30_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_39_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_41_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_28_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_12_30_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_43_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_9_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_9_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_45_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_47_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_31_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_49_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_8_30_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_51_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_31_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_53_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_31_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_for_tmp_bit_sva_1, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_5_31_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_55_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva_mx1w0,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_30_sva_mx1w0, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_57_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_sva_mx1w0, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_30_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_59_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_sva_mx1w0, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_29_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_mux1h_61_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_28_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_29_31_sva_mx1w0, EdgeDetect_MagAng_calc_crc32_32_1_crc_tmp_4_28_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_mux1h_1_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva_1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_9_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_1_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_30_sva_mx1w0,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_27_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_30_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_3_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_sva_mx1w0,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_5_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva_mx1w0,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_25_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_7_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_27_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_24_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_27_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_9_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_26_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_11_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_25_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_25_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_13_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_24_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_21_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_24_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_15_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_17_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_23_31_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_19_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_21_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_21_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_21_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_20_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_23_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_25_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_19_31_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_27_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_29_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_31_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_17_31_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_31_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_33_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_31_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_15_31_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_35_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_37_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_14_30_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_39_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_41_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_28_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_12_30_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_43_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_9_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_9_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_45_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_47_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_31_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_49_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_8_30_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_51_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_31_sva_mx1w1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_53_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_31_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_for_tmp_bit_sva_1, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_5_31_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_55_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva_mx1w0,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_30_sva_mx1w0, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_57_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_sva_mx1w0, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_30_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_59_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_sva_mx1w0, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_29_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign EdgeDetect_MagAng_calc_crc32_32_crc_tmp_mux1h_61_nl = MUX1HOT_s_1_3_2(EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_28_sva_mx1w1,
      EdgeDetect_MagAng_calc_crc32_32_crc_tmp_29_31_sva_mx1w0, EdgeDetect_MagAng_calc_crc32_32_crc_tmp_4_28_sva,
      {and_dcpl_7 , and_dcpl_9 , (~ MROW_stage_0)});
  assign MCOL_if_1_MCOL_if_1_or_nl = MROW_equal_tmp | (~ nor_cse);
  assign MROW_MROW_and_1_nl = (MROW_y_sva[8]) & (~ and_373_itm);
  assign MROW_mux_2_nl = MUX_v_8_2_2((MROW_y_sva[7:0]), MCOL_x_9_2_sva, and_373_itm);
  assign nl_z_out = ({MROW_MROW_and_1_nl , MROW_mux_2_nl}) + 9'b000000001;
  assign z_out = nl_z_out[8:0];

  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [7:0] signext_8_1;
    input  vector;
  begin
    signext_8_1= {{7{vector}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_1_8 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_8 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_VerDer
// ------------------------------------------------------------------


module EdgeDetect_VerDer (
  clk, rst, arst_n, dat_in_rsc_dat, dat_in_rsc_vld, dat_in_rsc_rdy, widthIn, heightIn,
      pix_out_rsc_dat, pix_out_rsc_vld, pix_out_rsc_rdy, dy_rsc_dat, dy_rsc_vld,
      dy_rsc_rdy, line_buf0_rsc_en, line_buf0_rsc_q, line_buf0_rsc_we, line_buf0_rsc_d,
      line_buf0_rsc_adr, line_buf1_rsc_en, line_buf1_rsc_q, line_buf1_rsc_we, line_buf1_rsc_d,
      line_buf1_rsc_adr
);
  input clk;
  input rst;
  input arst_n;
  input [33:0] dat_in_rsc_dat;
  input dat_in_rsc_vld;
  output dat_in_rsc_rdy;
  input [9:0] widthIn;
  input [8:0] heightIn;
  output [31:0] pix_out_rsc_dat;
  output pix_out_rsc_vld;
  input pix_out_rsc_rdy;
  output [35:0] dy_rsc_dat;
  output dy_rsc_vld;
  input dy_rsc_rdy;
  output line_buf0_rsc_en;
  input [63:0] line_buf0_rsc_q;
  output line_buf0_rsc_we;
  output [63:0] line_buf0_rsc_d;
  output [6:0] line_buf0_rsc_adr;
  output line_buf1_rsc_en;
  input [63:0] line_buf1_rsc_q;
  output line_buf1_rsc_we;
  output [63:0] line_buf1_rsc_d;
  output [6:0] line_buf1_rsc_adr;


  // Interconnect Declarations
  wire [63:0] line_buf0_rsci_d_d;
  wire line_buf0_rsci_en_d;
  wire [63:0] line_buf0_rsci_q_d;
  wire [63:0] line_buf1_rsci_d_d;
  wire [63:0] line_buf1_rsci_q_d;
  wire [6:0] line_buf0_rsci_adr_d_iff;
  wire line_buf0_rsci_we_d_iff;
  wire line_buf0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_iff;


  // Interconnect Declarations for Component Instantiations 
  EdgeDetect_VerDer_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_6_64_7_80_80_64_5_gen
      line_buf0_rsci (
      .en(line_buf0_rsc_en),
      .q(line_buf0_rsc_q),
      .we(line_buf0_rsc_we),
      .d(line_buf0_rsc_d),
      .adr(line_buf0_rsc_adr),
      .adr_d(line_buf0_rsci_adr_d_iff),
      .d_d(line_buf0_rsci_d_d),
      .en_d(line_buf0_rsci_en_d),
      .we_d(line_buf0_rsci_we_d_iff),
      .q_d(line_buf0_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(line_buf0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_iff),
      .port_0_rw_ram_ir_internal_WMASK_B_d(line_buf0_rsci_we_d_iff)
    );
  EdgeDetect_VerDer_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_7_64_7_80_80_64_5_gen
      line_buf1_rsci (
      .en(line_buf1_rsc_en),
      .q(line_buf1_rsc_q),
      .we(line_buf1_rsc_we),
      .d(line_buf1_rsc_d),
      .adr(line_buf1_rsc_adr),
      .adr_d(line_buf0_rsci_adr_d_iff),
      .d_d(line_buf1_rsci_d_d),
      .en_d(line_buf0_rsci_en_d),
      .we_d(line_buf0_rsci_we_d_iff),
      .q_d(line_buf1_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(line_buf0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_iff),
      .port_0_rw_ram_ir_internal_WMASK_B_d(line_buf0_rsci_we_d_iff)
    );
  EdgeDetect_VerDer_run EdgeDetect_VerDer_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .dat_in_rsc_dat(dat_in_rsc_dat),
      .dat_in_rsc_vld(dat_in_rsc_vld),
      .dat_in_rsc_rdy(dat_in_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .pix_out_rsc_dat(pix_out_rsc_dat),
      .pix_out_rsc_vld(pix_out_rsc_vld),
      .pix_out_rsc_rdy(pix_out_rsc_rdy),
      .dy_rsc_dat(dy_rsc_dat),
      .dy_rsc_vld(dy_rsc_vld),
      .dy_rsc_rdy(dy_rsc_rdy),
      .line_buf0_rsci_d_d(line_buf0_rsci_d_d),
      .line_buf0_rsci_en_d(line_buf0_rsci_en_d),
      .line_buf0_rsci_q_d(line_buf0_rsci_q_d),
      .line_buf1_rsci_d_d(line_buf1_rsci_d_d),
      .line_buf1_rsci_q_d(line_buf1_rsci_q_d),
      .line_buf0_rsci_adr_d_pff(line_buf0_rsci_adr_d_iff),
      .line_buf0_rsci_we_d_pff(line_buf0_rsci_we_d_iff),
      .line_buf0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_pff(line_buf0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_HorDer
// ------------------------------------------------------------------


module EdgeDetect_HorDer (
  clk, rst, arst_n, pix_in_rsc_dat, pix_in_rsc_vld, pix_in_rsc_rdy, widthIn, heightIn,
      pix_out_rsc_dat, pix_out_rsc_vld, pix_out_rsc_rdy, dx_rsc_dat, dx_rsc_vld,
      dx_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] pix_in_rsc_dat;
  input pix_in_rsc_vld;
  output pix_in_rsc_rdy;
  input [9:0] widthIn;
  input [8:0] heightIn;
  output [31:0] pix_out_rsc_dat;
  output pix_out_rsc_vld;
  input pix_out_rsc_rdy;
  output [35:0] dx_rsc_dat;
  output dx_rsc_vld;
  input dx_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  EdgeDetect_HorDer_run EdgeDetect_HorDer_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .pix_in_rsc_dat(pix_in_rsc_dat),
      .pix_in_rsc_vld(pix_in_rsc_vld),
      .pix_in_rsc_rdy(pix_in_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .pix_out_rsc_dat(pix_out_rsc_dat),
      .pix_out_rsc_vld(pix_out_rsc_vld),
      .pix_out_rsc_rdy(pix_out_rsc_rdy),
      .dx_rsc_dat(dx_rsc_dat),
      .dx_rsc_vld(dx_rsc_vld),
      .dx_rsc_rdy(dx_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_MagAng
// ------------------------------------------------------------------


module EdgeDetect_MagAng (
  clk, rst, arst_n, dx_in_rsc_dat, dx_in_rsc_vld, dx_in_rsc_rdy, dy_in_rsc_dat, dy_in_rsc_vld,
      dy_in_rsc_rdy, pix_in_rsc_dat, pix_in_rsc_vld, pix_in_rsc_rdy, widthIn, heightIn,
      sw_in, crc32_pix_in_rsc_dat, crc32_pix_in_triosy_lz, crc32_dat_out_rsc_dat,
      crc32_dat_out_triosy_lz, dat_out_rsc_dat, dat_out_rsc_vld, dat_out_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input [35:0] dx_in_rsc_dat;
  input dx_in_rsc_vld;
  output dx_in_rsc_rdy;
  input [35:0] dy_in_rsc_dat;
  input dy_in_rsc_vld;
  output dy_in_rsc_rdy;
  input [31:0] pix_in_rsc_dat;
  input pix_in_rsc_vld;
  output pix_in_rsc_rdy;
  input [9:0] widthIn;
  input [8:0] heightIn;
  input sw_in;
  output [31:0] crc32_pix_in_rsc_dat;
  output crc32_pix_in_triosy_lz;
  output [31:0] crc32_dat_out_rsc_dat;
  output crc32_dat_out_triosy_lz;
  output [33:0] dat_out_rsc_dat;
  output dat_out_rsc_vld;
  input dat_out_rsc_rdy;


  // Interconnect Declarations
  wire [31:0] crc32_pix_in_rsci_idat;
  wire [31:0] crc32_dat_out_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_v1 #(.rscid(32'sd20),
  .width(32'sd32)) crc32_pix_in_rsci (
      .idat(crc32_pix_in_rsci_idat),
      .dat(crc32_pix_in_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd21),
  .width(32'sd32)) crc32_dat_out_rsci (
      .idat(crc32_dat_out_rsci_idat),
      .dat(crc32_dat_out_rsc_dat)
    );
  EdgeDetect_MagAng_run EdgeDetect_MagAng_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .dx_in_rsc_dat(dx_in_rsc_dat),
      .dx_in_rsc_vld(dx_in_rsc_vld),
      .dx_in_rsc_rdy(dx_in_rsc_rdy),
      .dy_in_rsc_dat(dy_in_rsc_dat),
      .dy_in_rsc_vld(dy_in_rsc_vld),
      .dy_in_rsc_rdy(dy_in_rsc_rdy),
      .pix_in_rsc_dat(pix_in_rsc_dat),
      .pix_in_rsc_vld(pix_in_rsc_vld),
      .pix_in_rsc_rdy(pix_in_rsc_rdy),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .sw_in(sw_in),
      .crc32_pix_in_triosy_lz(crc32_pix_in_triosy_lz),
      .crc32_dat_out_triosy_lz(crc32_dat_out_triosy_lz),
      .dat_out_rsc_dat(dat_out_rsc_dat),
      .dat_out_rsc_vld(dat_out_rsc_vld),
      .dat_out_rsc_rdy(dat_out_rsc_rdy),
      .crc32_pix_in_rsci_idat(crc32_pix_in_rsci_idat),
      .crc32_dat_out_rsci_idat(crc32_dat_out_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_Top_struct
// ------------------------------------------------------------------


module EdgeDetect_Top_struct (
  clk, rst, arst_n, widthIn, heightIn, sw_in, crc32_pix_in_rsc_dat, crc32_pix_in_triosy_lz,
      crc32_dat_out_rsc_dat, crc32_dat_out_triosy_lz, dat_in_rsc_dat_eol, dat_in_rsc_dat_sof,
      dat_in_rsc_dat_pix, dat_in_rsc_vld, dat_in_rsc_rdy, dat_out_rsc_dat_eol, dat_out_rsc_dat_sof,
      dat_out_rsc_dat_pix, dat_out_rsc_vld, dat_out_rsc_rdy, line_buf0_rsc_en, line_buf0_rsc_q,
      line_buf0_rsc_we, line_buf0_rsc_d, line_buf0_rsc_adr, line_buf1_rsc_en, line_buf1_rsc_q,
      line_buf1_rsc_we, line_buf1_rsc_d, line_buf1_rsc_adr
);
  input clk;
  input rst;
  input arst_n;
  input [9:0] widthIn;
  input [8:0] heightIn;
  input sw_in;
  output [31:0] crc32_pix_in_rsc_dat;
  output crc32_pix_in_triosy_lz;
  output [31:0] crc32_dat_out_rsc_dat;
  output crc32_dat_out_triosy_lz;
  input dat_in_rsc_dat_eol;
  input dat_in_rsc_dat_sof;
  input [31:0] dat_in_rsc_dat_pix;
  input dat_in_rsc_vld;
  output dat_in_rsc_rdy;
  output dat_out_rsc_dat_eol;
  output dat_out_rsc_dat_sof;
  output [31:0] dat_out_rsc_dat_pix;
  output dat_out_rsc_vld;
  input dat_out_rsc_rdy;
  output line_buf0_rsc_en;
  input [63:0] line_buf0_rsc_q;
  output line_buf0_rsc_we;
  output [63:0] line_buf0_rsc_d;
  output [6:0] line_buf0_rsc_adr;
  output line_buf1_rsc_en;
  input [63:0] line_buf1_rsc_q;
  output line_buf1_rsc_we;
  output [63:0] line_buf1_rsc_d;
  output [6:0] line_buf1_rsc_adr;


  // Interconnect Declarations
  wire [31:0] pix_out_rsc_dat_n_VerDer_inst;
  wire [35:0] dy_rsc_dat_n_VerDer_inst;
  wire dy_rsc_rdy_n_VerDer_inst;
  wire line_buf0_rsc_en_n_VerDer_inst;
  wire [63:0] line_buf0_rsc_d_n_VerDer_inst;
  wire [6:0] line_buf0_rsc_adr_n_VerDer_inst;
  wire line_buf1_rsc_en_n_VerDer_inst;
  wire [63:0] line_buf1_rsc_d_n_VerDer_inst;
  wire [6:0] line_buf1_rsc_adr_n_VerDer_inst;
  wire [31:0] pix_out_rsc_dat_n_HorDer_inst;
  wire [35:0] dx_rsc_dat_n_HorDer_inst;
  wire [35:0] dy_in_rsc_dat_n_MagAng_inst;
  wire dy_in_rsc_vld_n_MagAng_inst;
  wire [31:0] crc32_pix_in_rsc_dat_n_MagAng_inst;
  wire [31:0] crc32_dat_out_rsc_dat_n_MagAng_inst;
  wire [33:0] dat_out_rsc_dat_n_MagAng_inst;
  wire dat_in_rsc_rdy_n_VerDer_inst_bud;
  wire pix_out_rsc_vld_n_VerDer_inst_bud;
  wire pix_in_rsc_rdy_n_HorDer_inst_bud;
  wire dy_rsc_vld_n_VerDer_inst_bud;
  wire dy_in_rsc_rdy_n_MagAng_inst_bud;
  wire line_buf0_rsc_we_n_VerDer_inst_bud;
  wire line_buf1_rsc_we_n_VerDer_inst_bud;
  wire pix_out_rsc_vld_n_HorDer_inst_bud;
  wire pix_in_rsc_rdy_n_MagAng_inst_bud;
  wire dx_rsc_vld_n_HorDer_inst_bud;
  wire dx_in_rsc_rdy_n_MagAng_inst_bud;
  wire crc32_pix_in_triosy_lz_n_MagAng_inst_bud;
  wire crc32_dat_out_triosy_lz_n_MagAng_inst_bud;
  wire dat_out_rsc_vld_n_MagAng_inst_bud;
  wire dy_chan_unc_1;
  wire dy_chan_idle;


  // Interconnect Declarations for Component Instantiations 
  wire [33:0] nl_VerDer_inst_dat_in_rsc_dat;
  assign nl_VerDer_inst_dat_in_rsc_dat = {dat_in_rsc_dat_eol , dat_in_rsc_dat_sof
      , dat_in_rsc_dat_pix};
  ccs_pipe_v6 #(.rscid(32'sd35),
  .width(32'sd36),
  .sz_width(32'sd1),
  .fifo_sz(32'sd2),
  .log2_sz(32'sd1),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd1)) dy_chan_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(rst),
      .din_rdy(dy_rsc_rdy_n_VerDer_inst),
      .din_vld(dy_rsc_vld_n_VerDer_inst_bud),
      .din(dy_rsc_dat_n_VerDer_inst),
      .dout_rdy(dy_in_rsc_rdy_n_MagAng_inst_bud),
      .dout_vld(dy_in_rsc_vld_n_MagAng_inst),
      .dout(dy_in_rsc_dat_n_MagAng_inst),
      .sz(dy_chan_unc_1),
      .sz_req(1'b0),
      .is_idle(dy_chan_idle)
    );
  EdgeDetect_VerDer VerDer_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .dat_in_rsc_dat(nl_VerDer_inst_dat_in_rsc_dat[33:0]),
      .dat_in_rsc_vld(dat_in_rsc_vld),
      .dat_in_rsc_rdy(dat_in_rsc_rdy_n_VerDer_inst_bud),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .pix_out_rsc_dat(pix_out_rsc_dat_n_VerDer_inst),
      .pix_out_rsc_vld(pix_out_rsc_vld_n_VerDer_inst_bud),
      .pix_out_rsc_rdy(pix_in_rsc_rdy_n_HorDer_inst_bud),
      .dy_rsc_dat(dy_rsc_dat_n_VerDer_inst),
      .dy_rsc_vld(dy_rsc_vld_n_VerDer_inst_bud),
      .dy_rsc_rdy(dy_rsc_rdy_n_VerDer_inst),
      .line_buf0_rsc_en(line_buf0_rsc_en_n_VerDer_inst),
      .line_buf0_rsc_q(line_buf0_rsc_q),
      .line_buf0_rsc_we(line_buf0_rsc_we_n_VerDer_inst_bud),
      .line_buf0_rsc_d(line_buf0_rsc_d_n_VerDer_inst),
      .line_buf0_rsc_adr(line_buf0_rsc_adr_n_VerDer_inst),
      .line_buf1_rsc_en(line_buf1_rsc_en_n_VerDer_inst),
      .line_buf1_rsc_q(line_buf1_rsc_q),
      .line_buf1_rsc_we(line_buf1_rsc_we_n_VerDer_inst_bud),
      .line_buf1_rsc_d(line_buf1_rsc_d_n_VerDer_inst),
      .line_buf1_rsc_adr(line_buf1_rsc_adr_n_VerDer_inst)
    );
  EdgeDetect_HorDer HorDer_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .pix_in_rsc_dat(pix_out_rsc_dat_n_VerDer_inst),
      .pix_in_rsc_vld(pix_out_rsc_vld_n_VerDer_inst_bud),
      .pix_in_rsc_rdy(pix_in_rsc_rdy_n_HorDer_inst_bud),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .pix_out_rsc_dat(pix_out_rsc_dat_n_HorDer_inst),
      .pix_out_rsc_vld(pix_out_rsc_vld_n_HorDer_inst_bud),
      .pix_out_rsc_rdy(pix_in_rsc_rdy_n_MagAng_inst_bud),
      .dx_rsc_dat(dx_rsc_dat_n_HorDer_inst),
      .dx_rsc_vld(dx_rsc_vld_n_HorDer_inst_bud),
      .dx_rsc_rdy(dx_in_rsc_rdy_n_MagAng_inst_bud)
    );
  EdgeDetect_MagAng MagAng_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .dx_in_rsc_dat(dx_rsc_dat_n_HorDer_inst),
      .dx_in_rsc_vld(dx_rsc_vld_n_HorDer_inst_bud),
      .dx_in_rsc_rdy(dx_in_rsc_rdy_n_MagAng_inst_bud),
      .dy_in_rsc_dat(dy_in_rsc_dat_n_MagAng_inst),
      .dy_in_rsc_vld(dy_in_rsc_vld_n_MagAng_inst),
      .dy_in_rsc_rdy(dy_in_rsc_rdy_n_MagAng_inst_bud),
      .pix_in_rsc_dat(pix_out_rsc_dat_n_HorDer_inst),
      .pix_in_rsc_vld(pix_out_rsc_vld_n_HorDer_inst_bud),
      .pix_in_rsc_rdy(pix_in_rsc_rdy_n_MagAng_inst_bud),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .sw_in(sw_in),
      .crc32_pix_in_rsc_dat(crc32_pix_in_rsc_dat_n_MagAng_inst),
      .crc32_pix_in_triosy_lz(crc32_pix_in_triosy_lz_n_MagAng_inst_bud),
      .crc32_dat_out_rsc_dat(crc32_dat_out_rsc_dat_n_MagAng_inst),
      .crc32_dat_out_triosy_lz(crc32_dat_out_triosy_lz_n_MagAng_inst_bud),
      .dat_out_rsc_dat(dat_out_rsc_dat_n_MagAng_inst),
      .dat_out_rsc_vld(dat_out_rsc_vld_n_MagAng_inst_bud),
      .dat_out_rsc_rdy(dat_out_rsc_rdy)
    );
  assign dat_out_rsc_dat_pix = dat_out_rsc_dat_n_MagAng_inst[31:0];
  assign dat_out_rsc_dat_sof = dat_out_rsc_dat_n_MagAng_inst[32];
  assign dat_out_rsc_dat_eol = dat_out_rsc_dat_n_MagAng_inst[33];
  assign dat_in_rsc_rdy = dat_in_rsc_rdy_n_VerDer_inst_bud;
  assign line_buf0_rsc_en = line_buf0_rsc_en_n_VerDer_inst;
  assign line_buf0_rsc_we = line_buf0_rsc_we_n_VerDer_inst_bud;
  assign line_buf0_rsc_d = line_buf0_rsc_d_n_VerDer_inst;
  assign line_buf0_rsc_adr = line_buf0_rsc_adr_n_VerDer_inst;
  assign line_buf1_rsc_en = line_buf1_rsc_en_n_VerDer_inst;
  assign line_buf1_rsc_we = line_buf1_rsc_we_n_VerDer_inst_bud;
  assign line_buf1_rsc_d = line_buf1_rsc_d_n_VerDer_inst;
  assign line_buf1_rsc_adr = line_buf1_rsc_adr_n_VerDer_inst;
  assign crc32_pix_in_rsc_dat = crc32_pix_in_rsc_dat_n_MagAng_inst;
  assign crc32_pix_in_triosy_lz = crc32_pix_in_triosy_lz_n_MagAng_inst_bud;
  assign crc32_dat_out_rsc_dat = crc32_dat_out_rsc_dat_n_MagAng_inst;
  assign crc32_dat_out_triosy_lz = crc32_dat_out_triosy_lz_n_MagAng_inst_bud;
  assign dat_out_rsc_vld = dat_out_rsc_vld_n_MagAng_inst_bud;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    EdgeDetect_Top
// ------------------------------------------------------------------


module EdgeDetect_Top (
  clk, rst, arst_n, widthIn, heightIn, sw_in, crc32_pix_in_rsc_dat, crc32_pix_in_triosy_lz,
      crc32_dat_out_rsc_dat, crc32_dat_out_triosy_lz, dat_in_rsc_dat, dat_in_rsc_vld,
      dat_in_rsc_rdy, dat_out_rsc_dat, dat_out_rsc_vld, dat_out_rsc_rdy, line_buf0_rsc_en,
      line_buf0_rsc_q, line_buf0_rsc_we, line_buf0_rsc_d, line_buf0_rsc_adr, line_buf1_rsc_en,
      line_buf1_rsc_q, line_buf1_rsc_we, line_buf1_rsc_d, line_buf1_rsc_adr
);
  input clk;
  input rst;
  input arst_n;
  input [9:0] widthIn;
  input [8:0] heightIn;
  input sw_in;
  output [31:0] crc32_pix_in_rsc_dat;
  output crc32_pix_in_triosy_lz;
  output [31:0] crc32_dat_out_rsc_dat;
  output crc32_dat_out_triosy_lz;
  input [33:0] dat_in_rsc_dat;
  input dat_in_rsc_vld;
  output dat_in_rsc_rdy;
  output [33:0] dat_out_rsc_dat;
  output dat_out_rsc_vld;
  input dat_out_rsc_rdy;
  output line_buf0_rsc_en;
  input [63:0] line_buf0_rsc_q;
  output line_buf0_rsc_we;
  output [63:0] line_buf0_rsc_d;
  output [6:0] line_buf0_rsc_adr;
  output line_buf1_rsc_en;
  input [63:0] line_buf1_rsc_q;
  output line_buf1_rsc_we;
  output [63:0] line_buf1_rsc_d;
  output [6:0] line_buf1_rsc_adr;


  // Interconnect Declarations
  wire dat_out_rsc_dat_eol;
  wire dat_out_rsc_dat_sof;
  wire [31:0] dat_out_rsc_dat_pix;


  // Interconnect Declarations for Component Instantiations 
  wire  nl_EdgeDetect_Top_struct_inst_dat_in_rsc_dat_eol;
  assign nl_EdgeDetect_Top_struct_inst_dat_in_rsc_dat_eol = dat_in_rsc_dat[33];
  wire  nl_EdgeDetect_Top_struct_inst_dat_in_rsc_dat_sof;
  assign nl_EdgeDetect_Top_struct_inst_dat_in_rsc_dat_sof = dat_in_rsc_dat[32];
  wire [31:0] nl_EdgeDetect_Top_struct_inst_dat_in_rsc_dat_pix;
  assign nl_EdgeDetect_Top_struct_inst_dat_in_rsc_dat_pix = dat_in_rsc_dat[31:0];
  EdgeDetect_Top_struct EdgeDetect_Top_struct_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .widthIn(widthIn),
      .heightIn(heightIn),
      .sw_in(sw_in),
      .crc32_pix_in_rsc_dat(crc32_pix_in_rsc_dat),
      .crc32_pix_in_triosy_lz(crc32_pix_in_triosy_lz),
      .crc32_dat_out_rsc_dat(crc32_dat_out_rsc_dat),
      .crc32_dat_out_triosy_lz(crc32_dat_out_triosy_lz),
      .dat_in_rsc_dat_eol(nl_EdgeDetect_Top_struct_inst_dat_in_rsc_dat_eol),
      .dat_in_rsc_dat_sof(nl_EdgeDetect_Top_struct_inst_dat_in_rsc_dat_sof),
      .dat_in_rsc_dat_pix(nl_EdgeDetect_Top_struct_inst_dat_in_rsc_dat_pix[31:0]),
      .dat_in_rsc_vld(dat_in_rsc_vld),
      .dat_in_rsc_rdy(dat_in_rsc_rdy),
      .dat_out_rsc_dat_eol(dat_out_rsc_dat_eol),
      .dat_out_rsc_dat_sof(dat_out_rsc_dat_sof),
      .dat_out_rsc_dat_pix(dat_out_rsc_dat_pix),
      .dat_out_rsc_vld(dat_out_rsc_vld),
      .dat_out_rsc_rdy(dat_out_rsc_rdy),
      .line_buf0_rsc_en(line_buf0_rsc_en),
      .line_buf0_rsc_q(line_buf0_rsc_q),
      .line_buf0_rsc_we(line_buf0_rsc_we),
      .line_buf0_rsc_d(line_buf0_rsc_d),
      .line_buf0_rsc_adr(line_buf0_rsc_adr),
      .line_buf1_rsc_en(line_buf1_rsc_en),
      .line_buf1_rsc_q(line_buf1_rsc_q),
      .line_buf1_rsc_we(line_buf1_rsc_we),
      .line_buf1_rsc_d(line_buf1_rsc_d),
      .line_buf1_rsc_adr(line_buf1_rsc_adr)
    );
  assign dat_out_rsc_dat = {dat_out_rsc_dat_eol , dat_out_rsc_dat_sof , dat_out_rsc_dat_pix};
endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Wed May 22 01:04:35 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    In_copy_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_2_64_10_1024_1024_64_5_gen
// ------------------------------------------------------------------


module In_copy_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_2_64_10_1024_1024_64_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [9:0] adr;
  input [9:0] adr_d;
  input [63:0] d_d;
  input en_d;
  input we_d;
  output [63:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module In_copy_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output, for_C_3_tr0
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [6:0] fsm_output;
  reg [6:0] fsm_output;
  input for_C_3_tr0;


  // FSM State Type Declaration for In_copy_run_run_fsm_1
  parameter
    run_rlp_C_0 = 3'd0,
    main_C_0 = 3'd1,
    for_C_0 = 3'd2,
    for_C_1 = 3'd3,
    for_C_2 = 3'd4,
    for_C_3 = 3'd5,
    main_C_1 = 3'd6;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : In_copy_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 7'b0000010;
        state_var_NS = for_C_0;
      end
      for_C_0 : begin
        fsm_output = 7'b0000100;
        state_var_NS = for_C_1;
      end
      for_C_1 : begin
        fsm_output = 7'b0001000;
        state_var_NS = for_C_2;
      end
      for_C_2 : begin
        fsm_output = 7'b0010000;
        state_var_NS = for_C_3;
      end
      for_C_3 : begin
        fsm_output = 7'b0100000;
        if ( for_C_3_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 7'b1000000;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 7'b0000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy_run_staller
// ------------------------------------------------------------------


module In_copy_run_staller (
  clk, rst, arst_n, run_wen, run_wten, in_data_rsci_wen_comp, ap_done_rsci_wen_comp,
      ap_start_rsci_wen_comp
);
  input clk;
  input rst;
  input arst_n;
  output run_wen;
  output run_wten;
  reg run_wten;
  input in_data_rsci_wen_comp;
  input ap_done_rsci_wen_comp;
  input ap_start_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = in_data_rsci_wen_comp & ap_done_rsci_wen_comp & ap_start_rsci_wen_comp;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten <= 1'b0;
    end
    else if ( rst ) begin
      run_wten <= 1'b0;
    end
    else begin
      run_wten <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy_run_mode_triosy_obj_mode_triosy_wait_ctrl
// ------------------------------------------------------------------


module In_copy_run_mode_triosy_obj_mode_triosy_wait_ctrl (
  run_wten, mode_triosy_obj_iswt0, mode_triosy_obj_biwt
);
  input run_wten;
  input mode_triosy_obj_iswt0;
  output mode_triosy_obj_biwt;



  // Interconnect Declarations for Component Instantiations 
  assign mode_triosy_obj_biwt = (~ run_wten) & mode_triosy_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy_run_qin_triosy_obj_qin_triosy_wait_ctrl
// ------------------------------------------------------------------


module In_copy_run_qin_triosy_obj_qin_triosy_wait_ctrl (
  run_wten, qin_triosy_obj_iswt0, qin_triosy_obj_biwt
);
  input run_wten;
  input qin_triosy_obj_iswt0;
  output qin_triosy_obj_biwt;



  // Interconnect Declarations for Component Instantiations 
  assign qin_triosy_obj_biwt = (~ run_wten) & qin_triosy_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy_run_ap_start_rsci_ap_start_wait_ctrl
// ------------------------------------------------------------------


module In_copy_run_ap_start_rsci_ap_start_wait_ctrl (
  ap_start_rsci_iswt0, ap_start_rsci_biwt, ap_start_rsci_ivld
);
  input ap_start_rsci_iswt0;
  output ap_start_rsci_biwt;
  input ap_start_rsci_ivld;



  // Interconnect Declarations for Component Instantiations 
  assign ap_start_rsci_biwt = ap_start_rsci_iswt0 & ap_start_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy_run_ap_done_rsci_ap_done_wait_ctrl
// ------------------------------------------------------------------


module In_copy_run_ap_done_rsci_ap_done_wait_ctrl (
  ap_done_rsci_iswt0, ap_done_rsci_biwt, ap_done_rsci_irdy
);
  input ap_done_rsci_iswt0;
  output ap_done_rsci_biwt;
  input ap_done_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign ap_done_rsci_biwt = ap_done_rsci_iswt0 & ap_done_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy_run_wait_dp
// ------------------------------------------------------------------


module In_copy_run_wait_dp (
  qin_rsci_en_d, run_wen, qin_rsci_cgo, qin_rsci_cgo_ir_unreg
);
  output qin_rsci_en_d;
  input run_wen;
  input qin_rsci_cgo;
  input qin_rsci_cgo_ir_unreg;



  // Interconnect Declarations for Component Instantiations 
  assign qin_rsci_en_d = run_wen & (qin_rsci_cgo | qin_rsci_cgo_ir_unreg);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy_run_in_data_rsci_in_data_wait_ctrl
// ------------------------------------------------------------------


module In_copy_run_in_data_rsci_in_data_wait_ctrl (
  in_data_rsci_iswt0, in_data_rsci_biwt, in_data_rsci_ivld
);
  input in_data_rsci_iswt0;
  output in_data_rsci_biwt;
  input in_data_rsci_ivld;



  // Interconnect Declarations for Component Instantiations 
  assign in_data_rsci_biwt = in_data_rsci_iswt0 & in_data_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy_run_mode_triosy_obj
// ------------------------------------------------------------------


module In_copy_run_mode_triosy_obj (
  mode_triosy_lz, run_wten, mode_triosy_obj_iswt0
);
  output mode_triosy_lz;
  input run_wten;
  input mode_triosy_obj_iswt0;


  // Interconnect Declarations
  wire mode_triosy_obj_biwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) mode_triosy_obj (
      .ld(mode_triosy_obj_biwt),
      .lz(mode_triosy_lz)
    );
  In_copy_run_mode_triosy_obj_mode_triosy_wait_ctrl In_copy_run_mode_triosy_obj_mode_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .mode_triosy_obj_iswt0(mode_triosy_obj_iswt0),
      .mode_triosy_obj_biwt(mode_triosy_obj_biwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy_run_qin_triosy_obj
// ------------------------------------------------------------------


module In_copy_run_qin_triosy_obj (
  qin_triosy_lz, run_wten, qin_triosy_obj_iswt0
);
  output qin_triosy_lz;
  input run_wten;
  input qin_triosy_obj_iswt0;


  // Interconnect Declarations
  wire qin_triosy_obj_biwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) qin_triosy_obj (
      .ld(qin_triosy_obj_biwt),
      .lz(qin_triosy_lz)
    );
  In_copy_run_qin_triosy_obj_qin_triosy_wait_ctrl In_copy_run_qin_triosy_obj_qin_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .qin_triosy_obj_iswt0(qin_triosy_obj_iswt0),
      .qin_triosy_obj_biwt(qin_triosy_obj_biwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy_run_ap_start_rsci
// ------------------------------------------------------------------


module In_copy_run_ap_start_rsci (
  ap_start_rsc_dat, ap_start_rsc_vld, ap_start_rsc_rdy, ap_start_rsci_oswt, ap_start_rsci_wen_comp
);
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  input ap_start_rsci_oswt;
  output ap_start_rsci_wen_comp;


  // Interconnect Declarations
  wire ap_start_rsci_biwt;
  wire ap_start_rsci_ivld;
  wire ap_start_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd4),
  .width(32'sd1)) ap_start_rsci (
      .rdy(ap_start_rsc_rdy),
      .vld(ap_start_rsc_vld),
      .dat(ap_start_rsc_dat),
      .irdy(ap_start_rsci_oswt),
      .ivld(ap_start_rsci_ivld),
      .idat(ap_start_rsci_idat)
    );
  In_copy_run_ap_start_rsci_ap_start_wait_ctrl In_copy_run_ap_start_rsci_ap_start_wait_ctrl_inst
      (
      .ap_start_rsci_iswt0(ap_start_rsci_oswt),
      .ap_start_rsci_biwt(ap_start_rsci_biwt),
      .ap_start_rsci_ivld(ap_start_rsci_ivld)
    );
  assign ap_start_rsci_wen_comp = (~ ap_start_rsci_oswt) | ap_start_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy_run_ap_done_rsci
// ------------------------------------------------------------------


module In_copy_run_ap_done_rsci (
  ap_done_rsc_dat, ap_done_rsc_vld, ap_done_rsc_rdy, ap_done_rsci_oswt, ap_done_rsci_wen_comp
);
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input ap_done_rsci_oswt;
  output ap_done_rsci_wen_comp;


  // Interconnect Declarations
  wire ap_done_rsci_biwt;
  wire ap_done_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd1)) ap_done_rsci (
      .irdy(ap_done_rsci_irdy),
      .ivld(ap_done_rsci_oswt),
      .idat(1'b1),
      .rdy(ap_done_rsc_rdy),
      .vld(ap_done_rsc_vld),
      .dat(ap_done_rsc_dat)
    );
  In_copy_run_ap_done_rsci_ap_done_wait_ctrl In_copy_run_ap_done_rsci_ap_done_wait_ctrl_inst
      (
      .ap_done_rsci_iswt0(ap_done_rsci_oswt),
      .ap_done_rsci_biwt(ap_done_rsci_biwt),
      .ap_done_rsci_irdy(ap_done_rsci_irdy)
    );
  assign ap_done_rsci_wen_comp = (~ ap_done_rsci_oswt) | ap_done_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy_run_in_data_rsci
// ------------------------------------------------------------------


module In_copy_run_in_data_rsci (
  in_data_rsc_dat, in_data_rsc_vld, in_data_rsc_rdy, in_data_rsci_oswt, in_data_rsci_wen_comp,
      in_data_rsci_idat_mxwt
);
  input [31:0] in_data_rsc_dat;
  input in_data_rsc_vld;
  output in_data_rsc_rdy;
  input in_data_rsci_oswt;
  output in_data_rsci_wen_comp;
  output [31:0] in_data_rsci_idat_mxwt;


  // Interconnect Declarations
  wire in_data_rsci_biwt;
  wire in_data_rsci_ivld;
  wire [31:0] in_data_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd32)) in_data_rsci (
      .rdy(in_data_rsc_rdy),
      .vld(in_data_rsc_vld),
      .dat(in_data_rsc_dat),
      .irdy(in_data_rsci_oswt),
      .ivld(in_data_rsci_ivld),
      .idat(in_data_rsci_idat)
    );
  In_copy_run_in_data_rsci_in_data_wait_ctrl In_copy_run_in_data_rsci_in_data_wait_ctrl_inst
      (
      .in_data_rsci_iswt0(in_data_rsci_oswt),
      .in_data_rsci_biwt(in_data_rsci_biwt),
      .in_data_rsci_ivld(in_data_rsci_ivld)
    );
  assign in_data_rsci_idat_mxwt = in_data_rsci_idat;
  assign in_data_rsci_wen_comp = (~ in_data_rsci_oswt) | in_data_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy_run
// ------------------------------------------------------------------


module In_copy_run (
  clk, rst, arst_n, in_data_rsc_dat, in_data_rsc_vld, in_data_rsc_rdy, qin_triosy_lz,
      ap_done_rsc_dat, ap_done_rsc_vld, ap_done_rsc_rdy, ap_start_rsc_dat, ap_start_rsc_vld,
      ap_start_rsc_rdy, mode_rsc_dat, mode_triosy_lz, qin_rsci_adr_d, qin_rsci_d_d,
      qin_rsci_en_d, qin_rsci_we_d_pff
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] in_data_rsc_dat;
  input in_data_rsc_vld;
  output in_data_rsc_rdy;
  output qin_triosy_lz;
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  input mode_rsc_dat;
  output mode_triosy_lz;
  output [9:0] qin_rsci_adr_d;
  output [63:0] qin_rsci_d_d;
  output qin_rsci_en_d;
  output qin_rsci_we_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire in_data_rsci_wen_comp;
  wire [31:0] in_data_rsci_idat_mxwt;
  wire ap_done_rsci_wen_comp;
  wire ap_start_rsci_wen_comp;
  wire mode_rsci_idat;
  wire [6:0] fsm_output;
  wire [10:0] for_x_10_0_sva_2;
  wire [11:0] nl_for_x_10_0_sva_2;
  reg for_io_read_mode_rsc_svs_st;
  reg reg_mode_triosy_obj_iswt0_cse;
  reg reg_ap_start_rsci_iswt0_cse;
  reg reg_qin_rsci_cgo_ir_cse;
  reg reg_in_data_rsci_iswt0_cse;
  wire or_5_rmff;
  reg [31:0] tmp1_63_32_sva_dfm_1;
  reg [31:0] for_mux_1_itm_1;
  reg [9:0] for_x_10_0_sva_9_0;

  wire[31:0] for_if_mux_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_In_copy_run_run_fsm_inst_for_C_3_tr0;
  assign nl_In_copy_run_run_fsm_inst_for_C_3_tr0 = for_x_10_0_sva_2[10];
  ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd1)) mode_rsci (
      .dat(mode_rsc_dat),
      .idat(mode_rsci_idat)
    );
  In_copy_run_in_data_rsci In_copy_run_in_data_rsci_inst (
      .in_data_rsc_dat(in_data_rsc_dat),
      .in_data_rsc_vld(in_data_rsc_vld),
      .in_data_rsc_rdy(in_data_rsc_rdy),
      .in_data_rsci_oswt(reg_in_data_rsci_iswt0_cse),
      .in_data_rsci_wen_comp(in_data_rsci_wen_comp),
      .in_data_rsci_idat_mxwt(in_data_rsci_idat_mxwt)
    );
  In_copy_run_wait_dp In_copy_run_wait_dp_inst (
      .qin_rsci_en_d(qin_rsci_en_d),
      .run_wen(run_wen),
      .qin_rsci_cgo(reg_qin_rsci_cgo_ir_cse),
      .qin_rsci_cgo_ir_unreg(or_5_rmff)
    );
  In_copy_run_ap_done_rsci In_copy_run_ap_done_rsci_inst (
      .ap_done_rsc_dat(ap_done_rsc_dat),
      .ap_done_rsc_vld(ap_done_rsc_vld),
      .ap_done_rsc_rdy(ap_done_rsc_rdy),
      .ap_done_rsci_oswt(reg_mode_triosy_obj_iswt0_cse),
      .ap_done_rsci_wen_comp(ap_done_rsci_wen_comp)
    );
  In_copy_run_ap_start_rsci In_copy_run_ap_start_rsci_inst (
      .ap_start_rsc_dat(ap_start_rsc_dat),
      .ap_start_rsc_vld(ap_start_rsc_vld),
      .ap_start_rsc_rdy(ap_start_rsc_rdy),
      .ap_start_rsci_oswt(reg_ap_start_rsci_iswt0_cse),
      .ap_start_rsci_wen_comp(ap_start_rsci_wen_comp)
    );
  In_copy_run_qin_triosy_obj In_copy_run_qin_triosy_obj_inst (
      .qin_triosy_lz(qin_triosy_lz),
      .run_wten(run_wten),
      .qin_triosy_obj_iswt0(reg_mode_triosy_obj_iswt0_cse)
    );
  In_copy_run_mode_triosy_obj In_copy_run_mode_triosy_obj_inst (
      .mode_triosy_lz(mode_triosy_lz),
      .run_wten(run_wten),
      .mode_triosy_obj_iswt0(reg_mode_triosy_obj_iswt0_cse)
    );
  In_copy_run_staller In_copy_run_staller_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .in_data_rsci_wen_comp(in_data_rsci_wen_comp),
      .ap_done_rsci_wen_comp(ap_done_rsci_wen_comp),
      .ap_start_rsci_wen_comp(ap_start_rsci_wen_comp)
    );
  In_copy_run_run_fsm In_copy_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .for_C_3_tr0(nl_In_copy_run_run_fsm_inst_for_C_3_tr0)
    );
  assign or_5_rmff = (fsm_output[5:4]!=2'b00);
  assign nl_for_x_10_0_sva_2 = conv_u2s_10_11(for_x_10_0_sva_9_0) + 11'b00000000001;
  assign for_x_10_0_sva_2 = nl_for_x_10_0_sva_2[10:0];
  assign qin_rsci_adr_d = for_x_10_0_sva_9_0;
  assign for_if_mux_nl = MUX_v_32_2_2(in_data_rsci_idat_mxwt, tmp1_63_32_sva_dfm_1,
      for_io_read_mode_rsc_svs_st);
  assign qin_rsci_d_d = {for_if_mux_nl , for_mux_1_itm_1};
  assign qin_rsci_we_d_pff = fsm_output[4];
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_mode_triosy_obj_iswt0_cse <= 1'b0;
      reg_ap_start_rsci_iswt0_cse <= 1'b0;
      reg_qin_rsci_cgo_ir_cse <= 1'b0;
      reg_in_data_rsci_iswt0_cse <= 1'b0;
      for_mux_1_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      reg_mode_triosy_obj_iswt0_cse <= 1'b0;
      reg_ap_start_rsci_iswt0_cse <= 1'b0;
      reg_qin_rsci_cgo_ir_cse <= 1'b0;
      reg_in_data_rsci_iswt0_cse <= 1'b0;
      for_mux_1_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen ) begin
      reg_mode_triosy_obj_iswt0_cse <= (for_x_10_0_sva_2[10]) & (fsm_output[5]);
      reg_ap_start_rsci_iswt0_cse <= (fsm_output[6]) | (fsm_output[0]);
      reg_qin_rsci_cgo_ir_cse <= or_5_rmff;
      reg_in_data_rsci_iswt0_cse <= ((~ for_io_read_mode_rsc_svs_st) & (fsm_output[3]))
          | (fsm_output[2]);
      for_mux_1_itm_1 <= in_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      tmp1_63_32_sva_dfm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      tmp1_63_32_sva_dfm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & (~ for_io_read_mode_rsc_svs_st) & (fsm_output[4]) ) begin
      tmp1_63_32_sva_dfm_1 <= in_data_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_x_10_0_sva_9_0 <= 10'b0000000000;
    end
    else if ( rst ) begin
      for_x_10_0_sva_9_0 <= 10'b0000000000;
    end
    else if ( run_wen & ((fsm_output[1]) | (fsm_output[5])) ) begin
      for_x_10_0_sva_9_0 <= MUX_v_10_2_2(10'b0000000000, (for_x_10_0_sva_2[9:0]),
          (fsm_output[5]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_io_read_mode_rsc_svs_st <= 1'b0;
    end
    else if ( rst ) begin
      for_io_read_mode_rsc_svs_st <= 1'b0;
    end
    else if ( run_wen & (fsm_output[2]) ) begin
      for_io_read_mode_rsc_svs_st <= mode_rsci_idat;
    end
  end

  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input  sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    In_copy
// ------------------------------------------------------------------


module In_copy (
  clk, rst, arst_n, in_data_rsc_dat, in_data_rsc_vld, in_data_rsc_rdy, qin_rsc_adr,
      qin_rsc_d, qin_rsc_we, qin_rsc_q, qin_rsc_en, qin_triosy_lz, ap_done_rsc_dat,
      ap_done_rsc_vld, ap_done_rsc_rdy, ap_start_rsc_dat, ap_start_rsc_vld, ap_start_rsc_rdy,
      mode_rsc_dat, mode_triosy_lz
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] in_data_rsc_dat;
  input in_data_rsc_vld;
  output in_data_rsc_rdy;
  output [9:0] qin_rsc_adr;
  output [63:0] qin_rsc_d;
  output qin_rsc_we;
  input [63:0] qin_rsc_q;
  output qin_rsc_en;
  output qin_triosy_lz;
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  input mode_rsc_dat;
  output mode_triosy_lz;


  // Interconnect Declarations
  wire [9:0] qin_rsci_adr_d;
  wire [63:0] qin_rsci_d_d;
  wire qin_rsci_en_d;
  wire [63:0] qin_rsci_q_d;
  wire qin_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  In_copy_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_2_64_10_1024_1024_64_5_gen
      qin_rsci (
      .en(qin_rsc_en),
      .q(qin_rsc_q),
      .we(qin_rsc_we),
      .d(qin_rsc_d),
      .adr(qin_rsc_adr),
      .adr_d(qin_rsci_adr_d),
      .d_d(qin_rsci_d_d),
      .en_d(qin_rsci_en_d),
      .we_d(qin_rsci_we_d_iff),
      .q_d(qin_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(qin_rsci_we_d_iff)
    );
  In_copy_run In_copy_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .in_data_rsc_dat(in_data_rsc_dat),
      .in_data_rsc_vld(in_data_rsc_vld),
      .in_data_rsc_rdy(in_data_rsc_rdy),
      .qin_triosy_lz(qin_triosy_lz),
      .ap_done_rsc_dat(ap_done_rsc_dat),
      .ap_done_rsc_vld(ap_done_rsc_vld),
      .ap_done_rsc_rdy(ap_done_rsc_rdy),
      .ap_start_rsc_dat(ap_start_rsc_dat),
      .ap_start_rsc_vld(ap_start_rsc_vld),
      .ap_start_rsc_rdy(ap_start_rsc_rdy),
      .mode_rsc_dat(mode_rsc_dat),
      .mode_triosy_lz(mode_triosy_lz),
      .qin_rsci_adr_d(qin_rsci_adr_d),
      .qin_rsci_d_d(qin_rsci_d_d),
      .qin_rsci_en_d(qin_rsci_en_d),
      .qin_rsci_we_d_pff(qin_rsci_we_d_iff)
    );
endmodule



module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);
  parameter integer rscid = 1;
  parameter integer width = 8;
  output [width-1:0] idat;
  output rdy;
  output ivld;
  input [width-1:0] dat;
  input irdy;
  input vld;
  wire [width-1:0] idat;
  wire rdy;
  wire ivld;
  localparam stallOff = 0;
  wire stall_ctrl;
  assign stall_ctrl = stallOff;
  assign idat = dat;
  assign rdy = irdy && !stall_ctrl;
  assign ivld = vld && !stall_ctrl;
endmodule
module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);
  parameter integer rscid = 1;
  parameter integer width = 8;
  output [width-1:0] dat;
  output irdy;
  output vld;
  input [width-1:0] idat;
  input rdy;
  input ivld;
  wire [width-1:0] dat;
  wire irdy;
  wire vld;
  localparam stallOff = 0;
  wire stall_ctrl;
  assign stall_ctrl = stallOff;
  assign dat = idat;
  assign irdy = rdy && !stall_ctrl;
  assign vld = ivld && !stall_ctrl;
endmodule
module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;
    input ld;
    output lz;
    wire lz;
    assign lz = ld;
endmodule
module ccs_in_v1 (idat, dat);
  parameter integer rscid = 1;
  parameter integer width = 8;
  output [width-1:0] idat;
  input [width-1:0] dat;
  wire [width-1:0] idat;
  assign idat = dat;
endmodule
module leading_sign_57_0_1_0 (
  mantissa, all_same, rtn
);
  input [56:0] mantissa;
  output all_same;
  output [5:0] rtn;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_18_3_sdt_3;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_42_4_sdt_4;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_62_3_sdt_3;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_90_5_sdt_5;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_110_3_sdt_3;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_134_4_sdt_4;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_154_3_sdt_3;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_168_6_sdt_6;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_14_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_34_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_58_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_78_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_106_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_126_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_150_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_24;
  wire c_h_1_25;
  wire c_h_1_26;
  wire c_h_1_27;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_and_221_nl;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_and_219_nl;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_nl;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_or_4_nl;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_2 = ~((mantissa[54:53]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_1 = ~((mantissa[56:55]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_14_2_sdt_1 = ~((mantissa[52:51]!=2'b00));
  assign c_h_1_2 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_2;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_18_3_sdt_3 = (mantissa[50:49]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_14_2_sdt_1;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_2 = ~((mantissa[46:45]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_1 = ~((mantissa[48:47]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_34_2_sdt_1 = ~((mantissa[44:43]!=2'b00));
  assign c_h_1_5 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_18_3_sdt_3;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_42_4_sdt_4 = (mantissa[42:41]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_34_2_sdt_1 & c_h_1_5;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_2 = ~((mantissa[38:37]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_1 = ~((mantissa[40:39]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_58_2_sdt_1 = ~((mantissa[36:35]!=2'b00));
  assign c_h_1_9 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_2;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_62_3_sdt_3 = (mantissa[34:33]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_58_2_sdt_1;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_2 = ~((mantissa[30:29]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_1 = ~((mantissa[32:31]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_78_2_sdt_1 = ~((mantissa[28:27]!=2'b00));
  assign c_h_1_12 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_42_4_sdt_4;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_90_5_sdt_5 = (mantissa[26:25]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_78_2_sdt_1 & c_h_1_12
      & c_h_1_13;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_2 = ~((mantissa[22:21]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_1 = ~((mantissa[24:23]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_106_2_sdt_1 = ~((mantissa[20:19]!=2'b00));
  assign c_h_1_17 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_2;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_110_3_sdt_3 = (mantissa[18:17]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_106_2_sdt_1;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_2 = ~((mantissa[14:13]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_1 = ~((mantissa[16:15]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_126_2_sdt_1 = ~((mantissa[12:11]!=2'b00));
  assign c_h_1_20 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_110_3_sdt_3;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_134_4_sdt_4 = (mantissa[10:9]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_126_2_sdt_1 & c_h_1_20;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_2 = ~((mantissa[6:5]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_1 = ~((mantissa[8:7]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_150_2_sdt_1 = ~((mantissa[4:3]!=2'b00));
  assign c_h_1_24 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_2;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_154_3_sdt_3 = (mantissa[2:1]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_150_2_sdt_1;
  assign c_h_1_25 = c_h_1_24 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_154_3_sdt_3;
  assign c_h_1_26 = c_h_1_21 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_134_4_sdt_4;
  assign c_h_1_27 = c_h_1_14 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_90_5_sdt_5;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_168_6_sdt_6 = (~
      (mantissa[0])) & c_h_1_25 & c_h_1_26 & c_h_1_27;
  assign all_same = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_168_6_sdt_6;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_and_221_nl = c_h_1_14 &
      (c_h_1_26 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_90_5_sdt_5));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_and_219_nl = c_h_1_6 &
      (c_h_1_13 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_42_4_sdt_4))
      & (~((~(c_h_1_21 & (c_h_1_25 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_134_4_sdt_4))))
      & c_h_1_27));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_nl
      = c_h_1_2 & (c_h_1_5 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_18_3_sdt_3))
      & (~((~(c_h_1_9 & (c_h_1_12 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~((~(c_h_1_17 & (c_h_1_20 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_110_3_sdt_3))
      & (~((~(c_h_1_24 & (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_154_3_sdt_3)))
      & c_h_1_26)))) & c_h_1_27));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_1_nl
      = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_1 & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_14_2_sdt_1
      | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_2)) & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_34_2_sdt_1 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_58_2_sdt_1 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_2))
      & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_1 &
      (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_78_2_sdt_1 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_106_2_sdt_1 | (~
      return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_2)) & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_126_2_sdt_1 | (~
      return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_2)))) & c_h_1_21))
      & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_150_2_sdt_1 | (~
      return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_2)) & (~ c_h_1_25)))
      & c_h_1_26)))) & c_h_1_27));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_or_4_nl
      = ((~((mantissa[56]) | (~((mantissa[55:54]!=2'b01))))) & (~(((mantissa[52])
      | (~((mantissa[51:50]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[48]) | (~((mantissa[47:46]!=2'b01)))))
      & (~(((mantissa[44]) | (~((mantissa[43:42]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[40]) | (~((mantissa[39:38]!=2'b01))))) & (~(((mantissa[36])
      | (~((mantissa[35:34]!=2'b01)))) & c_h_1_9)) & (~((~((~((mantissa[32]) | (~((mantissa[31:30]!=2'b01)))))
      & (~(((mantissa[28]) | (~((mantissa[27:26]!=2'b01)))) & c_h_1_12)))) & c_h_1_13))))
      & c_h_1_14)) & (~((~((~((mantissa[24]) | (~((mantissa[23:22]!=2'b01))))) &
      (~(((mantissa[20]) | (~((mantissa[19:18]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[16])
      | (~((mantissa[15:14]!=2'b01))))) & (~(((mantissa[12]) | (~((mantissa[11:10]!=2'b01))))
      & c_h_1_20)))) & c_h_1_21)) & (~(((mantissa[8]) | (~((mantissa[7:6]!=2'b01)))
      | (((mantissa[4]) | (~((mantissa[3:2]!=2'b01)))) & c_h_1_24) | c_h_1_25) &
      c_h_1_26)))) & c_h_1_27))) | return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_168_6_sdt_6;
  assign rtn = {c_h_1_27 , return_add_generic_AC_RND_CONV_false_ls_all_sign_and_221_nl
      , return_add_generic_AC_RND_CONV_false_ls_all_sign_and_219_nl , return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_nl
      , return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_1_nl
      , return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_or_4_nl};
endmodule
module mgc_shift_r_v5(a,s,z);
   parameter width_a = 4;
   parameter signd_a = 1;
   parameter width_s = 2;
   parameter width_z = 8;
   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;
   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u = result[olen-1:0];
      end
   endfunction
endmodule
module leading_sign_53_0 (
  mantissa, rtn
);
  input [52:0] mantissa;
  output [5:0] rtn;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_18_3_sdt_3;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_42_4_sdt_4;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_62_3_sdt_3;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_90_5_sdt_5;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_110_3_sdt_3;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_134_4_sdt_4;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_14_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_34_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_58_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_78_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_106_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_126_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_23;
  wire c_h_1_24;
  wire c_h_1_25;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_205_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_216_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_3_nl;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_2
      = ~((mantissa[50:49]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_1
      = ~((mantissa[52:51]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_14_2_sdt_1
      = ~((mantissa[48:47]!=2'b00));
  assign c_h_1_2 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_2;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_18_3_sdt_3
      = (mantissa[46:45]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_14_2_sdt_1;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_2
      = ~((mantissa[42:41]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_1
      = ~((mantissa[44:43]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_34_2_sdt_1
      = ~((mantissa[40:39]!=2'b00));
  assign c_h_1_5 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_18_3_sdt_3;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_42_4_sdt_4
      = (mantissa[38:37]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_34_2_sdt_1
      & c_h_1_5;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_2
      = ~((mantissa[34:33]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_1
      = ~((mantissa[36:35]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_58_2_sdt_1
      = ~((mantissa[32:31]!=2'b00));
  assign c_h_1_9 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_2;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_62_3_sdt_3
      = (mantissa[30:29]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_58_2_sdt_1;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_2
      = ~((mantissa[26:25]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_1
      = ~((mantissa[28:27]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_78_2_sdt_1
      = ~((mantissa[24:23]!=2'b00));
  assign c_h_1_12 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_42_4_sdt_4;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_90_5_sdt_5
      = (mantissa[22:21]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_78_2_sdt_1
      & c_h_1_12 & c_h_1_13;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_2
      = ~((mantissa[18:17]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_1
      = ~((mantissa[20:19]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_106_2_sdt_1
      = ~((mantissa[16:15]!=2'b00));
  assign c_h_1_17 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_2;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_110_3_sdt_3
      = (mantissa[14:13]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_106_2_sdt_1;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_2
      = ~((mantissa[10:9]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_1
      = ~((mantissa[12:11]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_126_2_sdt_1
      = ~((mantissa[8:7]!=2'b00));
  assign c_h_1_20 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_110_3_sdt_3;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_134_4_sdt_4
      = (mantissa[6:5]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_126_2_sdt_1
      & c_h_1_20;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_2
      = ~((mantissa[2:1]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_1
      = ~((mantissa[4:3]!=2'b00));
  assign c_h_1_23 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_2;
  assign c_h_1_24 = c_h_1_21 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_25 = c_h_1_14 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_90_5_sdt_5;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_205_nl
      = c_h_1_14 & (c_h_1_24 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_90_5_sdt_5));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_nl
      = c_h_1_6 & (c_h_1_13 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_42_4_sdt_4))
      & (~((~(c_h_1_21 & (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_134_4_sdt_4)))
      & c_h_1_25));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_216_nl
      = c_h_1_2 & (c_h_1_5 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_18_3_sdt_3))
      & (~((~(c_h_1_9 & (c_h_1_12 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~((~(c_h_1_17 & (c_h_1_20 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_110_3_sdt_3))
      & (c_h_1_23 | (~ c_h_1_24)))) & c_h_1_25));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_1_nl
      = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_14_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_34_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_58_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_2))
      & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_78_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_106_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_2))
      & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_126_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_2))))
      & c_h_1_21)) & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_1
      & (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_2)))
      & c_h_1_24)))) & c_h_1_25));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_3_nl
      = ((~((mantissa[52]) | (~((mantissa[51:50]!=2'b01))))) & (~(((mantissa[48])
      | (~((mantissa[47:46]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[44]) | (~((mantissa[43:42]!=2'b01)))))
      & (~(((mantissa[40]) | (~((mantissa[39:38]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[36]) | (~((mantissa[35:34]!=2'b01))))) & (~(((mantissa[32])
      | (~((mantissa[31:30]!=2'b01)))) & c_h_1_9)) & (~((~((~((mantissa[28]) | (~((mantissa[27:26]!=2'b01)))))
      & (~(((mantissa[24]) | (~((mantissa[23:22]!=2'b01)))) & c_h_1_12)))) & c_h_1_13))))
      & c_h_1_14)) & (~((~((~((mantissa[20]) | (~((mantissa[19:18]!=2'b01))))) &
      (~(((mantissa[16]) | (~((mantissa[15:14]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[12])
      | (~((mantissa[11:10]!=2'b01))))) & (~(((mantissa[8]) | (~((mantissa[7:6]!=2'b01))))
      & c_h_1_20)))) & c_h_1_21)) & (~(((mantissa[4]) | (~((mantissa[3:2]!=2'b01)))
      | c_h_1_23) & c_h_1_24)))) & c_h_1_25))) | ((~ (mantissa[0])) & c_h_1_23 &
      c_h_1_24 & c_h_1_25);
  assign rtn = {c_h_1_25 , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_205_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_216_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_1_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_3_nl};
endmodule
module mgc_shift_l_v5(a,s,z);
   parameter width_a = 4;
   parameter signd_a = 1;
   parameter width_s = 2;
   parameter width_z = 8;
   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;
   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate
   function [width_z-1:0] fshl_u_1;
      input [width_a :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 = result[olen-1:0];
      end
   endfunction
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction
endmodule
module mgc_generic_reg (d, clk, en, a_rst, s_rst, q);
   parameter width = 8;
   parameter ph_clk = 1;
   parameter ph_en = 1;
   parameter ph_a_rst = 1;
   parameter ph_s_rst = 1;
   parameter a_rst_used = 1;
   parameter s_rst_used = 0;
   parameter en_used = 0;
   input [width-1:0] d;
   input clk;
   input en;
   input a_rst;
   input s_rst;
   output reg [width-1:0] q;
   generate
      if (ph_clk==1 && ph_a_rst==1)
      begin: GEN_CLK1_ARST1
         always@(posedge a_rst or posedge clk)
           if (a_rst == 1'b1)
             q <= {width{1'b0}};
           else if (s_rst == $unsigned(ph_s_rst))
             q <= {width{1'b0}};
           else if (en == $unsigned(ph_en))
             q <= d;
      end
      else if (ph_clk==1 && ph_a_rst==0)
      begin: GEN_CLK1_ARST0
         always@(negedge a_rst or posedge clk)
           if (a_rst == 1'b0)
             q <= {width{1'b0}};
           else if (s_rst == $unsigned(ph_s_rst))
             q <= {width{1'b0}};
           else if (en == $unsigned(ph_en))
             q <= d;
      end
      else if (ph_clk==0 && ph_a_rst==1)
      begin: GEN_CLK0_ARST1
         always@(posedge a_rst or negedge clk)
           if (a_rst == 1'b1)
             q <= {width{1'b0}};
           else if (s_rst == $unsigned(ph_s_rst))
             q <= {width{1'b0}};
           else if (en == $unsigned(ph_en))
             q <= d;
      end
      else if (ph_clk==0 && ph_a_rst==0)
      begin: GEN_CLK0_ARST0
         always@(negedge a_rst or negedge clk)
           if (a_rst == 1'b0)
             q <= {width{1'b0}};
           else if (s_rst == $unsigned(ph_s_rst))
             q <= {width{1'b0}};
           else if (en == $unsigned(ph_en))
             q <= d;
      end
   endgenerate
endmodule
module stagemgc_rom_sync_regout_14_1024_14_1_0_0_1_0_1_0_0_0_1_60 (addr, data_out,
    clk, s_rst, a_rst, en
);
  input [9:0]addr ;
  output [13:0]data_out ;
  input clk ;
  input s_rst ;
  input a_rst ;
  input en ;
  parameter n_width = 14;
  parameter n_size = 1024;
  parameter n_numports = 1;
  parameter n_addr_w = 10;
  parameter n_inreg = 0;
  parameter n_outreg = 1;
  wire [9:0] addr_f;
  wire [9:0] addr_reg [n_inreg:0];
  genvar i;
  generate if (n_inreg > 0)
  begin
    for( i=n_inreg-1; i >= 1; i=i-1)
    begin: addr_reg_stage
      mgc_generic_reg #(
        .width(10),
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_addr_reg (
        .d(addr_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(addr_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(10),
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_addr_reg_init (
      .d(addr),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(addr_reg[0])
    );
    assign addr_f = addr_reg[n_inreg-1];
  end
  else
  begin
    assign addr_f = addr;
  end
  endgenerate
  wire [13:0] mem [1023:0];
  reg [13:0] data_out_t;
  assign mem[0] = 14'b00111111111011;
  assign mem[1] = 14'b01111011010000;
  assign mem[2] = 14'b10101100110100;
  assign mem[3] = 14'b10101111001000;
  assign mem[4] = 14'b01101100110000;
  assign mem[5] = 14'b01000011110110;
  assign mem[6] = 14'b01100010000011;
  assign mem[7] = 14'b10011000011111;
  assign mem[8] = 14'b00011000110111;
  assign mem[9] = 14'b01100011111111;
  assign mem[10] = 14'b10010100000101;
  assign mem[11] = 14'b01010010010010;
  assign mem[12] = 14'b00001001001010;
  assign mem[13] = 14'b01011011000001;
  assign mem[14] = 14'b01110101110010;
  assign mem[15] = 14'b10010111101110;
  assign mem[16] = 14'b00010001101110;
  assign mem[17] = 14'b01100100000111;
  assign mem[18] = 14'b00011010101111;
  assign mem[19] = 14'b00001111000101;
  assign mem[20] = 14'b01101110111011;
  assign mem[21] = 14'b01110111111010;
  assign mem[22] = 14'b00111010011111;
  assign mem[23] = 14'b01100100101010;
  assign mem[24] = 14'b10100010101110;
  assign mem[25] = 14'b01111110100100;
  assign mem[26] = 14'b00011101011101;
  assign mem[27] = 14'b00011010011000;
  assign mem[28] = 14'b00010101010100;
  assign mem[29] = 14'b10100001011001;
  assign mem[30] = 14'b10011110110100;
  assign mem[31] = 14'b10001111011100;
  assign mem[32] = 14'b10111110110010;
  assign mem[33] = 14'b01100001100000;
  assign mem[34] = 14'b00001111100101;
  assign mem[35] = 14'b00000001110101;
  assign mem[36] = 14'b01001010101111;
  assign mem[37] = 14'b01000100110111;
  assign mem[38] = 14'b00011000001101;
  assign mem[39] = 14'b01101110100000;
  assign mem[40] = 14'b00101100001101;
  assign mem[41] = 14'b01100100111010;
  assign mem[42] = 14'b01000101001111;
  assign mem[43] = 14'b10001010101101;
  assign mem[44] = 14'b01101111101000;
  assign mem[45] = 14'b00101000000100;
  assign mem[46] = 14'b01011000100000;
  assign mem[47] = 14'b00111111001010;
  assign mem[48] = 14'b10111110011101;
  assign mem[49] = 14'b00000110110000;
  assign mem[50] = 14'b10100111111111;
  assign mem[51] = 14'b00010011010101;
  assign mem[52] = 14'b01110110111010;
  assign mem[53] = 14'b00010111111110;
  assign mem[54] = 14'b00111110001111;
  assign mem[55] = 14'b01111010110111;
  assign mem[56] = 14'b00100010000101;
  assign mem[57] = 14'b01100010100100;
  assign mem[58] = 14'b10001000010000;
  assign mem[59] = 14'b01100110101010;
  assign mem[60] = 14'b01001011101011;
  assign mem[61] = 14'b00011010011010;
  assign mem[62] = 14'b00000000001110;
  assign mem[63] = 14'b00111100100000;
  assign mem[64] = 14'b01010111000001;
  assign mem[65] = 14'b10010010011000;
  assign mem[66] = 14'b10111110000011;
  assign mem[67] = 14'b00011111100011;
  assign mem[68] = 14'b01110101110111;
  assign mem[69] = 14'b00100100001011;
  assign mem[70] = 14'b01001001000001;
  assign mem[71] = 14'b01110010101100;
  assign mem[72] = 14'b00011000010001;
  assign mem[73] = 14'b00010010000100;
  assign mem[74] = 14'b10000011010001;
  assign mem[75] = 14'b10110001111101;
  assign mem[76] = 14'b00001111111100;
  assign mem[77] = 14'b00101110010111;
  assign mem[78] = 14'b10101000010100;
  assign mem[79] = 14'b01101110000101;
  assign mem[80] = 14'b00110011110100;
  assign mem[81] = 14'b10101111100100;
  assign mem[82] = 14'b01010010100101;
  assign mem[83] = 14'b10110100111010;
  assign mem[84] = 14'b10100110001101;
  assign mem[85] = 14'b10011101100110;
  assign mem[86] = 14'b10010100010101;
  assign mem[87] = 14'b01100000100100;
  assign mem[88] = 14'b10010000111101;
  assign mem[89] = 14'b01011111110010;
  assign mem[90] = 14'b00110011111011;
  assign mem[91] = 14'b00001101110011;
  assign mem[92] = 14'b10100011100101;
  assign mem[93] = 14'b00000111101001;
  assign mem[94] = 14'b00010111011110;
  assign mem[95] = 14'b00101100100011;
  assign mem[96] = 14'b10101100110101;
  assign mem[97] = 14'b10011000000001;
  assign mem[98] = 14'b00101010110110;
  assign mem[99] = 14'b10111111010001;
  assign mem[100] = 14'b01001101101010;
  assign mem[101] = 14'b10100011110001;
  assign mem[102] = 14'b10011101011110;
  assign mem[103] = 14'b00010010101011;
  assign mem[104] = 14'b00001011011010;
  assign mem[105] = 14'b00011011100010;
  assign mem[106] = 14'b00111100001110;
  assign mem[107] = 14'b00011111101110;
  assign mem[108] = 14'b01011100000100;
  assign mem[109] = 14'b10101010101010;
  assign mem[110] = 14'b10001100111100;
  assign mem[111] = 14'b01010010011010;
  assign mem[112] = 14'b10001111011011;
  assign mem[113] = 14'b00111000010100;
  assign mem[114] = 14'b00111011000110;
  assign mem[115] = 14'b10011111011110;
  assign mem[116] = 14'b00110001101100;
  assign mem[117] = 14'b00110110001011;
  assign mem[118] = 14'b01001000111100;
  assign mem[119] = 14'b00100110001110;
  assign mem[120] = 14'b01110110111101;
  assign mem[121] = 14'b10010010101010;
  assign mem[122] = 14'b00001101000010;
  assign mem[123] = 14'b01111000010111;
  assign mem[124] = 14'b01101010110100;
  assign mem[125] = 14'b00110101001011;
  assign mem[126] = 14'b01010011100111;
  assign mem[127] = 14'b10111111110100;
  assign mem[128] = 14'b00110111111100;
  assign mem[129] = 14'b00011011001011;
  assign mem[130] = 14'b10101001000100;
  assign mem[131] = 14'b10011000111011;
  assign mem[132] = 14'b10011111100001;
  assign mem[133] = 14'b00111111100110;
  assign mem[134] = 14'b10111111011010;
  assign mem[135] = 14'b10000101001101;
  assign mem[136] = 14'b10100010100001;
  assign mem[137] = 14'b00101010111101;
  assign mem[138] = 14'b01110010101010;
  assign mem[139] = 14'b10100101001110;
  assign mem[140] = 14'b01011110011000;
  assign mem[141] = 14'b00001110101111;
  assign mem[142] = 14'b10010001110010;
  assign mem[143] = 14'b00010111000101;
  assign mem[144] = 14'b01101011010001;
  assign mem[145] = 14'b10010111000100;
  assign mem[146] = 14'b00111000000001;
  assign mem[147] = 14'b01100111101001;
  assign mem[148] = 14'b10111101110001;
  assign mem[149] = 14'b00111111011111;
  assign mem[150] = 14'b00111001100100;
  assign mem[151] = 14'b01111000000000;
  assign mem[152] = 14'b01111111111100;
  assign mem[153] = 14'b01101011110110;
  assign mem[154] = 14'b00110111001101;
  assign mem[155] = 14'b10011001001111;
  assign mem[156] = 14'b01011111001010;
  assign mem[157] = 14'b00001011010111;
  assign mem[158] = 14'b10011101110011;
  assign mem[159] = 14'b01101101011011;
  assign mem[160] = 14'b01101100100001;
  assign mem[161] = 14'b00011110011101;
  assign mem[162] = 14'b10011000000011;
  assign mem[163] = 14'b10100100111111;
  assign mem[164] = 14'b01011110101001;
  assign mem[165] = 14'b00000101111010;
  assign mem[166] = 14'b01111010111111;
  assign mem[167] = 14'b10001000111011;
  assign mem[168] = 14'b10001011000101;
  assign mem[169] = 14'b10010000001101;
  assign mem[170] = 14'b10001010001110;
  assign mem[171] = 14'b01000111000111;
  assign mem[172] = 14'b10010101110101;
  assign mem[173] = 14'b10110110010000;
  assign mem[174] = 14'b01110111001110;
  assign mem[175] = 14'b10001001110101;
  assign mem[176] = 14'b01011000110000;
  assign mem[177] = 14'b01001101011100;
  assign mem[178] = 14'b01100001101011;
  assign mem[179] = 14'b10000011000100;
  assign mem[180] = 14'b10011110101100;
  assign mem[181] = 14'b10001000010011;
  assign mem[182] = 14'b00100100100101;
  assign mem[183] = 14'b00110001010111;
  assign mem[184] = 14'b00010110111011;
  assign mem[185] = 14'b01010101010100;
  assign mem[186] = 14'b10000101101001;
  assign mem[187] = 14'b01111001100111;
  assign mem[188] = 14'b00101001011001;
  assign mem[189] = 14'b00100100010000;
  assign mem[190] = 14'b10001101001100;
  assign mem[191] = 14'b01100000101100;
  assign mem[192] = 14'b00001011100001;
  assign mem[193] = 14'b00111001110010;
  assign mem[194] = 14'b01001001011011;
  assign mem[195] = 14'b01011001111001;
  assign mem[196] = 14'b10001101010110;
  assign mem[197] = 14'b00111001100111;
  assign mem[198] = 14'b00000000010000;
  assign mem[199] = 14'b00001110010010;
  assign mem[200] = 14'b01010001000010;
  assign mem[201] = 14'b10100100100011;
  assign mem[202] = 14'b01000111001000;
  assign mem[203] = 14'b00011110101100;
  assign mem[204] = 14'b00110110110101;
  assign mem[205] = 14'b10000011110100;
  assign mem[206] = 14'b01110101011100;
  assign mem[207] = 14'b01010100000101;
  assign mem[208] = 14'b10100111101101;
  assign mem[209] = 14'b00110011010001;
  assign mem[210] = 14'b01101101111101;
  assign mem[211] = 14'b00010000100100;
  assign mem[212] = 14'b00101101001111;
  assign mem[213] = 14'b01101111110100;
  assign mem[214] = 14'b10001010110111;
  assign mem[215] = 14'b01010011101101;
  assign mem[216] = 14'b01100100001001;
  assign mem[217] = 14'b10000000000101;
  assign mem[218] = 14'b00101110010010;
  assign mem[219] = 14'b01100011100111;
  assign mem[220] = 14'b01001111001000;
  assign mem[221] = 14'b01100111101010;
  assign mem[222] = 14'b01010111111001;
  assign mem[223] = 14'b00000100010110;
  assign mem[224] = 14'b00001110100100;
  assign mem[225] = 14'b10011111110101;
  assign mem[226] = 14'b10001011011111;
  assign mem[227] = 14'b01110111011010;
  assign mem[228] = 14'b00000101011111;
  assign mem[229] = 14'b10010001010010;
  assign mem[230] = 14'b00000011101101;
  assign mem[231] = 14'b01011011100010;
  assign mem[232] = 14'b01111000001100;
  assign mem[233] = 14'b00110001001010;
  assign mem[234] = 14'b10111101011110;
  assign mem[235] = 14'b01110110100010;
  assign mem[236] = 14'b00100000000101;
  assign mem[237] = 14'b10110000010101;
  assign mem[238] = 14'b00111011011010;
  assign mem[239] = 14'b01010001010100;
  assign mem[240] = 14'b01000111111010;
  assign mem[241] = 14'b00011011010100;
  assign mem[242] = 14'b10110000100100;
  assign mem[243] = 14'b00000101010100;
  assign mem[244] = 14'b00111001111111;
  assign mem[245] = 14'b01001000000110;
  assign mem[246] = 14'b00000100101100;
  assign mem[247] = 14'b10101011110001;
  assign mem[248] = 14'b01001111001110;
  assign mem[249] = 14'b10011101000001;
  assign mem[250] = 14'b10110101100000;
  assign mem[251] = 14'b10111111010111;
  assign mem[252] = 14'b01110011111101;
  assign mem[253] = 14'b10100111010011;
  assign mem[254] = 14'b01011001110010;
  assign mem[255] = 14'b01011000010110;
  assign mem[256] = 14'b00111011111011;
  assign mem[257] = 14'b01010110110001;
  assign mem[258] = 14'b00010011001000;
  assign mem[259] = 14'b10000100011100;
  assign mem[260] = 14'b10010000010101;
  assign mem[261] = 14'b00111100000101;
  assign mem[262] = 14'b00000011111010;
  assign mem[263] = 14'b10101111001001;
  assign mem[264] = 14'b01000010000001;
  assign mem[265] = 14'b01100010110110;
  assign mem[266] = 14'b10010111010000;
  assign mem[267] = 14'b10111111011110;
  assign mem[268] = 14'b01000000101000;
  assign mem[269] = 14'b00101011011010;
  assign mem[270] = 14'b00001010110100;
  assign mem[271] = 14'b10001001101000;
  assign mem[272] = 14'b01100100001010;
  assign mem[273] = 14'b01101000111110;
  assign mem[274] = 14'b10011101111001;
  assign mem[275] = 14'b10100010110010;
  assign mem[276] = 14'b00111010101111;
  assign mem[277] = 14'b01110010111100;
  assign mem[278] = 14'b10110001100001;
  assign mem[279] = 14'b10000011110001;
  assign mem[280] = 14'b01100100100101;
  assign mem[281] = 14'b00111001000100;
  assign mem[282] = 14'b01100011000110;
  assign mem[283] = 14'b10001100010010;
  assign mem[284] = 14'b01010100001111;
  assign mem[285] = 14'b00100011100000;
  assign mem[286] = 14'b01100101001100;
  assign mem[287] = 14'b01110011111000;
  assign mem[288] = 14'b10000011100010;
  assign mem[289] = 14'b10101001001000;
  assign mem[290] = 14'b10111011010010;
  assign mem[291] = 14'b01011001100101;
  assign mem[292] = 14'b00001101101100;
  assign mem[293] = 14'b01101101110110;
  assign mem[294] = 14'b00100001110111;
  assign mem[295] = 14'b00100110000100;
  assign mem[296] = 14'b00110101110010;
  assign mem[297] = 14'b10010000000001;
  assign mem[298] = 14'b10000000001110;
  assign mem[299] = 14'b01001011111010;
  assign mem[300] = 14'b01011101001100;
  assign mem[301] = 14'b00101010111010;
  assign mem[302] = 14'b01110000001010;
  assign mem[303] = 14'b00010110011010;
  assign mem[304] = 14'b01110011011101;
  assign mem[305] = 14'b10001010101111;
  assign mem[306] = 14'b10100110100101;
  assign mem[307] = 14'b10110011000001;
  assign mem[308] = 14'b01000001111100;
  assign mem[309] = 14'b00010110011000;
  assign mem[310] = 14'b10101001010000;
  assign mem[311] = 14'b01000011101000;
  assign mem[312] = 14'b10000101101101;
  assign mem[313] = 14'b00011101001011;
  assign mem[314] = 14'b10010011101110;
  assign mem[315] = 14'b00100101110000;
  assign mem[316] = 14'b00111011101000;
  assign mem[317] = 14'b10001101110100;
  assign mem[318] = 14'b00001010101110;
  assign mem[319] = 14'b01010100010001;
  assign mem[320] = 14'b00100111011011;
  assign mem[321] = 14'b01000011110011;
  assign mem[322] = 14'b01011111100011;
  assign mem[323] = 14'b00001001101011;
  assign mem[324] = 14'b00001110101001;
  assign mem[325] = 14'b00101100010010;
  assign mem[326] = 14'b01111001011111;
  assign mem[327] = 14'b00110011001111;
  assign mem[328] = 14'b00100100111011;
  assign mem[329] = 14'b01110101000000;
  assign mem[330] = 14'b01011111100000;
  assign mem[331] = 14'b01001111000000;
  assign mem[332] = 14'b00001100111000;
  assign mem[333] = 14'b10011111011100;
  assign mem[334] = 14'b10110110101010;
  assign mem[335] = 14'b00010001011001;
  assign mem[336] = 14'b00101010100111;
  assign mem[337] = 14'b10011001111000;
  assign mem[338] = 14'b00001110000000;
  assign mem[339] = 14'b00011111101100;
  assign mem[340] = 14'b01001111010011;
  assign mem[341] = 14'b00101001011110;
  assign mem[342] = 14'b10100011100000;
  assign mem[343] = 14'b01111011001100;
  assign mem[344] = 14'b10111110001001;
  assign mem[345] = 14'b01010100111010;
  assign mem[346] = 14'b00101111111110;
  assign mem[347] = 14'b01100100000000;
  assign mem[348] = 14'b10001110101100;
  assign mem[349] = 14'b10110110011000;
  assign mem[350] = 14'b10111101111001;
  assign mem[351] = 14'b01000110101000;
  assign mem[352] = 14'b00010011111001;
  assign mem[353] = 14'b10011000001011;
  assign mem[354] = 14'b10110011001100;
  assign mem[355] = 14'b10011011010001;
  assign mem[356] = 14'b10011100110111;
  assign mem[357] = 14'b10010111111000;
  assign mem[358] = 14'b00100011010110;
  assign mem[359] = 14'b10010010110111;
  assign mem[360] = 14'b10101110111000;
  assign mem[361] = 14'b00000100111011;
  assign mem[362] = 14'b01000110011111;
  assign mem[363] = 14'b00010010000110;
  assign mem[364] = 14'b01011110101101;
  assign mem[365] = 14'b01101001011111;
  assign mem[366] = 14'b10111001011001;
  assign mem[367] = 14'b00000101100101;
  assign mem[368] = 14'b01110011000111;
  assign mem[369] = 14'b01000111000110;
  assign mem[370] = 14'b00001111010111;
  assign mem[371] = 14'b10000101010110;
  assign mem[372] = 14'b10000010100000;
  assign mem[373] = 14'b10011110001110;
  assign mem[374] = 14'b01110101101010;
  assign mem[375] = 14'b10010000100101;
  assign mem[376] = 14'b01000100001111;
  assign mem[377] = 14'b01010001100101;
  assign mem[378] = 14'b00111110011111;
  assign mem[379] = 14'b10001001001001;
  assign mem[380] = 14'b00110001011001;
  assign mem[381] = 14'b01101101001110;
  assign mem[382] = 14'b01000000100010;
  assign mem[383] = 14'b10110110000100;
  assign mem[384] = 14'b00110100101110;
  assign mem[385] = 14'b10110011010101;
  assign mem[386] = 14'b00011011011001;
  assign mem[387] = 14'b00000100100100;
  assign mem[388] = 14'b10000111101001;
  assign mem[389] = 14'b00101011110110;
  assign mem[390] = 14'b10100010001010;
  assign mem[391] = 14'b10111110011100;
  assign mem[392] = 14'b01011010101000;
  assign mem[393] = 14'b10111000100011;
  assign mem[394] = 14'b00110001101101;
  assign mem[395] = 14'b00011111000100;
  assign mem[396] = 14'b00010000000000;
  assign mem[397] = 14'b10010001111100;
  assign mem[398] = 14'b00100110101101;
  assign mem[399] = 14'b10101010110000;
  assign mem[400] = 14'b01000111100110;
  assign mem[401] = 14'b01101001011110;
  assign mem[402] = 14'b00111000100011;
  assign mem[403] = 14'b01010101111111;
  assign mem[404] = 14'b01010001110001;
  assign mem[405] = 14'b00100110011111;
  assign mem[406] = 14'b10000100010110;
  assign mem[407] = 14'b01110111100010;
  assign mem[408] = 14'b01111100011100;
  assign mem[409] = 14'b01100011111011;
  assign mem[410] = 14'b00010000101111;
  assign mem[411] = 14'b00010011111000;
  assign mem[412] = 14'b00110110010010;
  assign mem[413] = 14'b10101100100101;
  assign mem[414] = 14'b00110011011011;
  assign mem[415] = 14'b10110001010000;
  assign mem[416] = 14'b10000100110110;
  assign mem[417] = 14'b10010100000110;
  assign mem[418] = 14'b10011001101101;
  assign mem[419] = 14'b00010011100101;
  assign mem[420] = 14'b00011101000001;
  assign mem[421] = 14'b01100001011001;
  assign mem[422] = 14'b01001001110000;
  assign mem[423] = 14'b10110100101001;
  assign mem[424] = 14'b01011110010010;
  assign mem[425] = 14'b10011001011001;
  assign mem[426] = 14'b00110100001011;
  assign mem[427] = 14'b00011100000101;
  assign mem[428] = 14'b00101100111111;
  assign mem[429] = 14'b01100001100010;
  assign mem[430] = 14'b01010001010000;
  assign mem[431] = 14'b00100001000010;
  assign mem[432] = 14'b01111100011010;
  assign mem[433] = 14'b10010010001001;
  assign mem[434] = 14'b10110001100011;
  assign mem[435] = 14'b01010101100011;
  assign mem[436] = 14'b01011111000100;
  assign mem[437] = 14'b10010110000001;
  assign mem[438] = 14'b01000000001100;
  assign mem[439] = 14'b01110010011011;
  assign mem[440] = 14'b10100011000110;
  assign mem[441] = 14'b10010011111111;
  assign mem[442] = 14'b00010011110111;
  assign mem[443] = 14'b00000110011000;
  assign mem[444] = 14'b01101011111111;
  assign mem[445] = 14'b00110000000111;
  assign mem[446] = 14'b00000101101000;
  assign mem[447] = 14'b10000001010100;
  assign mem[448] = 14'b10110100001111;
  assign mem[449] = 14'b10001111000100;
  assign mem[450] = 14'b10001101011001;
  assign mem[451] = 14'b10110100010011;
  assign mem[452] = 14'b00001101010010;
  assign mem[453] = 14'b10000110101001;
  assign mem[454] = 14'b00001100010000;
  assign mem[455] = 14'b01111011101111;
  assign mem[456] = 14'b10000010001110;
  assign mem[457] = 14'b10111110001010;
  assign mem[458] = 14'b00011100110110;
  assign mem[459] = 14'b10011111100101;
  assign mem[460] = 14'b10111110011000;
  assign mem[461] = 14'b01111010010011;
  assign mem[462] = 14'b10111001111111;
  assign mem[463] = 14'b01010111100000;
  assign mem[464] = 14'b10011000110011;
  assign mem[465] = 14'b00001111110100;
  assign mem[466] = 14'b00001011010001;
  assign mem[467] = 14'b00101011100000;
  assign mem[468] = 14'b01101000010100;
  assign mem[469] = 14'b01100110011000;
  assign mem[470] = 14'b01010011100100;
  assign mem[471] = 14'b01000101001000;
  assign mem[472] = 14'b01101010100000;
  assign mem[473] = 14'b10000011010101;
  assign mem[474] = 14'b10011011100111;
  assign mem[475] = 14'b01010000011110;
  assign mem[476] = 14'b00100100110100;
  assign mem[477] = 14'b01010110110000;
  assign mem[478] = 14'b01010010010011;
  assign mem[479] = 14'b00010100110101;
  assign mem[480] = 14'b10001001100001;
  assign mem[481] = 14'b10010110111101;
  assign mem[482] = 14'b01110010001100;
  assign mem[483] = 14'b01011010011100;
  assign mem[484] = 14'b01001100101110;
  assign mem[485] = 14'b00001110001101;
  assign mem[486] = 14'b10110101011101;
  assign mem[487] = 14'b01000100101011;
  assign mem[488] = 14'b10000000101110;
  assign mem[489] = 14'b01101000011110;
  assign mem[490] = 14'b01000011001110;
  assign mem[491] = 14'b00101111100100;
  assign mem[492] = 14'b00100011101101;
  assign mem[493] = 14'b10111111011001;
  assign mem[494] = 14'b00011110101011;
  assign mem[495] = 14'b10010000000000;
  assign mem[496] = 14'b01000011001000;
  assign mem[497] = 14'b10111010001110;
  assign mem[498] = 14'b00001010110111;
  assign mem[499] = 14'b01000100010011;
  assign mem[500] = 14'b10011001000001;
  assign mem[501] = 14'b01001100010100;
  assign mem[502] = 14'b00100101101011;
  assign mem[503] = 14'b10011111110110;
  assign mem[504] = 14'b00101001011010;
  assign mem[505] = 14'b00001101001001;
  assign mem[506] = 14'b00111100110010;
  assign mem[507] = 14'b10011111110111;
  assign mem[508] = 14'b01110001010000;
  assign mem[509] = 14'b10000100111001;
  assign mem[510] = 14'b10101110111100;
  assign mem[511] = 14'b01101000100000;
  assign mem[512] = 14'b00111111011011;
  assign mem[513] = 14'b01011110101100;
  assign mem[514] = 14'b00111001100110;
  assign mem[515] = 14'b01001001110010;
  assign mem[516] = 14'b10111001001101;
  assign mem[517] = 14'b01011010111000;
  assign mem[518] = 14'b01101110010010;
  assign mem[519] = 14'b01101011010100;
  assign mem[520] = 14'b10101110000001;
  assign mem[521] = 14'b01111011110110;
  assign mem[522] = 14'b01001100011110;
  assign mem[523] = 14'b10111111111100;
  assign mem[524] = 14'b01000000000110;
  assign mem[525] = 14'b00111101000100;
  assign mem[526] = 14'b00111000011010;
  assign mem[527] = 14'b01100101111101;
  assign mem[528] = 14'b01111100000010;
  assign mem[529] = 14'b01111100101110;
  assign mem[530] = 14'b10111011001001;
  assign mem[531] = 14'b01101001100011;
  assign mem[532] = 14'b00001000011001;
  assign mem[533] = 14'b01000111010010;
  assign mem[534] = 14'b00011001010111;
  assign mem[535] = 14'b10000000100011;
  assign mem[536] = 14'b10110010111101;
  assign mem[537] = 14'b01110101111000;
  assign mem[538] = 14'b00001110001010;
  assign mem[539] = 14'b10111000101000;
  assign mem[540] = 14'b10010101001100;
  assign mem[541] = 14'b10101001101010;
  assign mem[542] = 14'b10010111100111;
  assign mem[543] = 14'b00101011111111;
  assign mem[544] = 14'b10110111011000;
  assign mem[545] = 14'b01101010011101;
  assign mem[546] = 14'b01101101000011;
  assign mem[547] = 14'b00001100110011;
  assign mem[548] = 14'b10001011000111;
  assign mem[549] = 14'b01100001111111;
  assign mem[550] = 14'b10101001011011;
  assign mem[551] = 14'b00000101011100;
  assign mem[552] = 14'b01110101011010;
  assign mem[553] = 14'b10000010010011;
  assign mem[554] = 14'b01100100100111;
  assign mem[555] = 14'b00001010110110;
  assign mem[556] = 14'b00001101010100;
  assign mem[557] = 14'b01011000011011;
  assign mem[558] = 14'b00101011011101;
  assign mem[559] = 14'b00111010000100;
  assign mem[560] = 14'b10110101000101;
  assign mem[561] = 14'b00101111010000;
  assign mem[562] = 14'b00010111110011;
  assign mem[563] = 14'b10000111010011;
  assign mem[564] = 14'b01000000010010;
  assign mem[565] = 14'b10100111110010;
  assign mem[566] = 14'b00110011100111;
  assign mem[567] = 14'b01011011111101;
  assign mem[568] = 14'b00101110100010;
  assign mem[569] = 14'b01110001111001;
  assign mem[570] = 14'b10111001101100;
  assign mem[571] = 14'b10001110100011;
  assign mem[572] = 14'b10010001101011;
  assign mem[573] = 14'b10111000110110;
  assign mem[574] = 14'b00000001100010;
  assign mem[575] = 14'b00100111011110;
  assign mem[576] = 14'b00100001000100;
  assign mem[577] = 14'b01000000100011;
  assign mem[578] = 14'b10110010001111;
  assign mem[579] = 14'b00011100110100;
  assign mem[580] = 14'b00111000111101;
  assign mem[581] = 14'b00111101001100;
  assign mem[582] = 14'b01111111000101;
  assign mem[583] = 14'b00100010110000;
  assign mem[584] = 14'b10101001110111;
  assign mem[585] = 14'b01111110011100;
  assign mem[586] = 14'b10010110110011;
  assign mem[587] = 14'b01011101100101;
  assign mem[588] = 14'b01101111100100;
  assign mem[589] = 14'b10000100100000;
  assign mem[590] = 14'b00011010000110;
  assign mem[591] = 14'b00000010011111;
  assign mem[592] = 14'b10101010101011;
  assign mem[593] = 14'b01001100110110;
  assign mem[594] = 14'b00000010000000;
  assign mem[595] = 14'b01110010010000;
  assign mem[596] = 14'b00001011010101;
  assign mem[597] = 14'b10001111000101;
  assign mem[598] = 14'b01001110001110;
  assign mem[599] = 14'b01100011111001;
  assign mem[600] = 14'b00110110100110;
  assign mem[601] = 14'b01011110011011;
  assign mem[602] = 14'b10101011011100;
  assign mem[603] = 14'b01100000100101;
  assign mem[604] = 14'b10111000111110;
  assign mem[605] = 14'b00110101011111;
  assign mem[606] = 14'b10100100010010;
  assign mem[607] = 14'b01110111110100;
  assign mem[608] = 14'b00111001101101;
  assign mem[609] = 14'b01101000000010;
  assign mem[610] = 14'b01101011111001;
  assign mem[611] = 14'b10111010110001;
  assign mem[612] = 14'b10011111100100;
  assign mem[613] = 14'b10111010010010;
  assign mem[614] = 14'b10001110001101;
  assign mem[615] = 14'b10000010101101;
  assign mem[616] = 14'b01001111110110;
  assign mem[617] = 14'b00000000101101;
  assign mem[618] = 14'b00100101100000;
  assign mem[619] = 14'b00011110000001;
  assign mem[620] = 14'b01000100011001;
  assign mem[621] = 14'b00101010100000;
  assign mem[622] = 14'b00011010011111;
  assign mem[623] = 14'b00000000110011;
  assign mem[624] = 14'b00101011111000;
  assign mem[625] = 14'b00001010001010;
  assign mem[626] = 14'b00011101101000;
  assign mem[627] = 14'b10011100001101;
  assign mem[628] = 14'b10011011110011;
  assign mem[629] = 14'b10111011001100;
  assign mem[630] = 14'b01111110100010;
  assign mem[631] = 14'b01001011100001;
  assign mem[632] = 14'b01000000100111;
  assign mem[633] = 14'b01000010100001;
  assign mem[634] = 14'b01011011001110;
  assign mem[635] = 14'b01001010011101;
  assign mem[636] = 14'b10101011101001;
  assign mem[637] = 14'b10110100001100;
  assign mem[638] = 14'b00001001001110;
  assign mem[639] = 14'b10111110100110;
  assign mem[640] = 14'b00000111100010;
  assign mem[641] = 14'b10111110001101;
  assign mem[642] = 14'b00011111010110;
  assign mem[643] = 14'b01101110011000;
  assign mem[644] = 14'b10011100100010;
  assign mem[645] = 14'b00111101001000;
  assign mem[646] = 14'b10111011110000;
  assign mem[647] = 14'b10100100010111;
  assign mem[648] = 14'b10110001100010;
  assign mem[649] = 14'b01101100101010;
  assign mem[650] = 14'b00100010100010;
  assign mem[651] = 14'b00000100011100;
  assign mem[652] = 14'b01010100100101;
  assign mem[653] = 14'b01100111001001;
  assign mem[654] = 14'b00111100011001;
  assign mem[655] = 14'b10100001100011;
  assign mem[656] = 14'b10101110110100;
  assign mem[657] = 14'b01100001010111;
  assign mem[658] = 14'b00001000000101;
  assign mem[659] = 14'b10010101011100;
  assign mem[660] = 14'b10110000010001;
  assign mem[661] = 14'b00111100010111;
  assign mem[662] = 14'b00010010111010;
  assign mem[663] = 14'b01000111111100;
  assign mem[664] = 14'b01111111100000;
  assign mem[665] = 14'b10110010110111;
  assign mem[666] = 14'b00000010011001;
  assign mem[667] = 14'b01110000100100;
  assign mem[668] = 14'b01011010000011;
  assign mem[669] = 14'b01001111100001;
  assign mem[670] = 14'b10010000100000;
  assign mem[671] = 14'b10111101111010;
  assign mem[672] = 14'b10110111100100;
  assign mem[673] = 14'b00010101001010;
  assign mem[674] = 14'b01101000010000;
  assign mem[675] = 14'b00000010110011;
  assign mem[676] = 14'b01010110011100;
  assign mem[677] = 14'b00101001010110;
  assign mem[678] = 14'b01011100110101;
  assign mem[679] = 14'b10111110011001;
  assign mem[680] = 14'b00001101011110;
  assign mem[681] = 14'b00110001010110;
  assign mem[682] = 14'b00000111011101;
  assign mem[683] = 14'b01110001101111;
  assign mem[684] = 14'b01011000101110;
  assign mem[685] = 14'b01111011101010;
  assign mem[686] = 14'b01000010011110;
  assign mem[687] = 14'b00000100101110;
  assign mem[688] = 14'b00101101001101;
  assign mem[689] = 14'b10011110000010;
  assign mem[690] = 14'b01101011101010;
  assign mem[691] = 14'b10010101011000;
  assign mem[692] = 14'b10010110101111;
  assign mem[693] = 14'b10111010000001;
  assign mem[694] = 14'b01000000000010;
  assign mem[695] = 14'b10011001100000;
  assign mem[696] = 14'b10100000011101;
  assign mem[697] = 14'b00010101001001;
  assign mem[698] = 14'b10100111011011;
  assign mem[699] = 14'b01010011001101;
  assign mem[700] = 14'b01100001101110;
  assign mem[701] = 14'b00111101101111;
  assign mem[702] = 14'b00011100001111;
  assign mem[703] = 14'b01100100110001;
  assign mem[704] = 14'b01010000100111;
  assign mem[705] = 14'b00010100011100;
  assign mem[706] = 14'b10000001111011;
  assign mem[707] = 14'b00110101001100;
  assign mem[708] = 14'b00011101010101;
  assign mem[709] = 14'b00010011001111;
  assign mem[710] = 14'b00000001110000;
  assign mem[711] = 14'b01100011111110;
  assign mem[712] = 14'b10110111001100;
  assign mem[713] = 14'b10111111110000;
  assign mem[714] = 14'b01110001110110;
  assign mem[715] = 14'b00010110110011;
  assign mem[716] = 14'b10111111110010;
  assign mem[717] = 14'b10011010101000;
  assign mem[718] = 14'b00110110000000;
  assign mem[719] = 14'b00001100100000;
  assign mem[720] = 14'b00010101110101;
  assign mem[721] = 14'b10100110110110;
  assign mem[722] = 14'b00000001100111;
  assign mem[723] = 14'b01110011111100;
  assign mem[724] = 14'b01111100101000;
  assign mem[725] = 14'b00001110101000;
  assign mem[726] = 14'b00001011111100;
  assign mem[727] = 14'b00001001111000;
  assign mem[728] = 14'b01111100111100;
  assign mem[729] = 14'b10000000011111;
  assign mem[730] = 14'b10000011111101;
  assign mem[731] = 14'b01111001001110;
  assign mem[732] = 14'b10101001110110;
  assign mem[733] = 14'b10010101100011;
  assign mem[734] = 14'b00100111001100;
  assign mem[735] = 14'b00011110011010;
  assign mem[736] = 14'b01100101111100;
  assign mem[737] = 14'b10011110101110;
  assign mem[738] = 14'b00010000010100;
  assign mem[739] = 14'b01000011110010;
  assign mem[740] = 14'b00100110011001;
  assign mem[741] = 14'b00111000111001;
  assign mem[742] = 14'b00011001111011;
  assign mem[743] = 14'b01000000101011;
  assign mem[744] = 14'b01001001010000;
  assign mem[745] = 14'b10011000000101;
  assign mem[746] = 14'b10101110001100;
  assign mem[747] = 14'b00111101101010;
  assign mem[748] = 14'b00100000100010;
  assign mem[749] = 14'b01010010001101;
  assign mem[750] = 14'b00011111110100;
  assign mem[751] = 14'b10111001001010;
  assign mem[752] = 14'b01110111010100;
  assign mem[753] = 14'b10111111001100;
  assign mem[754] = 14'b01010011110110;
  assign mem[755] = 14'b00100101001100;
  assign mem[756] = 14'b00010101110111;
  assign mem[757] = 14'b01111000101000;
  assign mem[758] = 14'b00100000110100;
  assign mem[759] = 14'b00110010010001;
  assign mem[760] = 14'b10101010100000;
  assign mem[761] = 14'b10001011000010;
  assign mem[762] = 14'b01110110011010;
  assign mem[763] = 14'b10111011011011;
  assign mem[764] = 14'b00101011100111;
  assign mem[765] = 14'b00010010111111;
  assign mem[766] = 14'b00110100011011;
  assign mem[767] = 14'b00101010010111;
  assign mem[768] = 14'b00100011011011;
  assign mem[769] = 14'b00011111010100;
  assign mem[770] = 14'b10000101111000;
  assign mem[771] = 14'b10011111000000;
  assign mem[772] = 14'b00110010001110;
  assign mem[773] = 14'b00100100100001;
  assign mem[774] = 14'b00011011010110;
  assign mem[775] = 14'b01001001111001;
  assign mem[776] = 14'b01001110000101;
  assign mem[777] = 14'b01110011110111;
  assign mem[778] = 14'b01100010101011;
  assign mem[779] = 14'b10111100001100;
  assign mem[780] = 14'b01000100010110;
  assign mem[781] = 14'b01101111110101;
  assign mem[782] = 14'b01001011101100;
  assign mem[783] = 14'b00000011010011;
  assign mem[784] = 14'b01111101000011;
  assign mem[785] = 14'b10011110101111;
  assign mem[786] = 14'b10010001001010;
  assign mem[787] = 14'b10110011011001;
  assign mem[788] = 14'b00011011000111;
  assign mem[789] = 14'b00100100100000;
  assign mem[790] = 14'b01011010100001;
  assign mem[791] = 14'b10011010010011;
  assign mem[792] = 14'b10000000000000;
  assign mem[793] = 14'b00001111011010;
  assign mem[794] = 14'b01110101100111;
  assign mem[795] = 14'b00010101111001;
  assign mem[796] = 14'b00001101100110;
  assign mem[797] = 14'b00111000011111;
  assign mem[798] = 14'b10000100010001;
  assign mem[799] = 14'b00101011000100;
  assign mem[800] = 14'b10011000101010;
  assign mem[801] = 14'b00011111110010;
  assign mem[802] = 14'b10011110111000;
  assign mem[803] = 14'b00110011000000;
  assign mem[804] = 14'b01011111110100;
  assign mem[805] = 14'b00000000110110;
  assign mem[806] = 14'b00101101000000;
  assign mem[807] = 14'b01001010011011;
  assign mem[808] = 14'b10111000011101;
  assign mem[809] = 14'b00110000000010;
  assign mem[810] = 14'b10000001011110;
  assign mem[811] = 14'b10010011010100;
  assign mem[812] = 14'b01001100010001;
  assign mem[813] = 14'b01101100010101;
  assign mem[814] = 14'b00010001000010;
  assign mem[815] = 14'b10011100110110;
  assign mem[816] = 14'b00101000000111;
  assign mem[817] = 14'b00001011000100;
  assign mem[818] = 14'b00001101111101;
  assign mem[819] = 14'b01100101000001;
  assign mem[820] = 14'b01001101100010;
  assign mem[821] = 14'b10011100101000;
  assign mem[822] = 14'b00100000101010;
  assign mem[823] = 14'b01011001010110;
  assign mem[824] = 14'b10100111110111;
  assign mem[825] = 14'b00001100001100;
  assign mem[826] = 14'b01001001111101;
  assign mem[827] = 14'b01001000001111;
  assign mem[828] = 14'b00100001010110;
  assign mem[829] = 14'b00100000100111;
  assign mem[830] = 14'b01001011000010;
  assign mem[831] = 14'b00001101110100;
  assign mem[832] = 14'b01010011111100;
  assign mem[833] = 14'b01011010100011;
  assign mem[834] = 14'b01011100110010;
  assign mem[835] = 14'b01000011101101;
  assign mem[836] = 14'b01100110011111;
  assign mem[837] = 14'b01110101111101;
  assign mem[838] = 14'b01010010010101;
  assign mem[839] = 14'b10100110101000;
  assign mem[840] = 14'b01000010011100;
  assign mem[841] = 14'b00110010111100;
  assign mem[842] = 14'b01011100011101;
  assign mem[843] = 14'b10101000111110;
  assign mem[844] = 14'b01011010001000;
  assign mem[845] = 14'b10011011111111;
  assign mem[846] = 14'b01111110100000;
  assign mem[847] = 14'b01111001101111;
  assign mem[848] = 14'b01101010010000;
  assign mem[849] = 14'b01110101000011;
  assign mem[850] = 14'b01100010000000;
  assign mem[851] = 14'b00011101110011;
  assign mem[852] = 14'b10101011000011;
  assign mem[853] = 14'b01100010010001;
  assign mem[854] = 14'b10111000011011;
  assign mem[855] = 14'b01011110010000;
  assign mem[856] = 14'b10110010111001;
  assign mem[857] = 14'b00010010010011;
  assign mem[858] = 14'b10001111110001;
  assign mem[859] = 14'b01111011111101;
  assign mem[860] = 14'b00100110101111;
  assign mem[861] = 14'b01111100100010;
  assign mem[862] = 14'b10110001001001;
  assign mem[863] = 14'b01101110010110;
  assign mem[864] = 14'b10001011001111;
  assign mem[865] = 14'b01101001001000;
  assign mem[866] = 14'b01100110001110;
  assign mem[867] = 14'b01111110110010;
  assign mem[868] = 14'b10001001111100;
  assign mem[869] = 14'b01100111000011;
  assign mem[870] = 14'b00110111011001;
  assign mem[871] = 14'b01000011111100;
  assign mem[872] = 14'b01001000000010;
  assign mem[873] = 14'b00100010011101;
  assign mem[874] = 14'b01101101010111;
  assign mem[875] = 14'b01111110101010;
  assign mem[876] = 14'b01010110111000;
  assign mem[877] = 14'b10100010010110;
  assign mem[878] = 14'b10010001101001;
  assign mem[879] = 14'b00100111000011;
  assign mem[880] = 14'b00100101101101;
  assign mem[881] = 14'b01110001101000;
  assign mem[882] = 14'b01101011100001;
  assign mem[883] = 14'b10100101010110;
  assign mem[884] = 14'b10010001011100;
  assign mem[885] = 14'b10010011011101;
  assign mem[886] = 14'b00110111100010;
  assign mem[887] = 14'b00110011111110;
  assign mem[888] = 14'b01011101100111;
  assign mem[889] = 14'b10111011000001;
  assign mem[890] = 14'b00110101010111;
  assign mem[891] = 14'b10111111111011;
  assign mem[892] = 14'b10011001101110;
  assign mem[893] = 14'b10111100011111;
  assign mem[894] = 14'b01000011101100;
  assign mem[895] = 14'b01111010010110;
  assign mem[896] = 14'b10110001000001;
  assign mem[897] = 14'b01100111001101;
  assign mem[898] = 14'b10111111101111;
  assign mem[899] = 14'b00011111111100;
  assign mem[900] = 14'b10110101011011;
  assign mem[901] = 14'b01110010111001;
  assign mem[902] = 14'b10101111000001;
  assign mem[903] = 14'b10110100111110;
  assign mem[904] = 14'b00111010010101;
  assign mem[905] = 14'b10001011101111;
  assign mem[906] = 14'b10011011111010;
  assign mem[907] = 14'b00011001011011;
  assign mem[908] = 14'b01110000000000;
  assign mem[909] = 14'b00111101011111;
  assign mem[910] = 14'b01001110111010;
  assign mem[911] = 14'b00101011001010;
  assign mem[912] = 14'b01110101001000;
  assign mem[913] = 14'b10100010001111;
  assign mem[914] = 14'b00001011110011;
  assign mem[915] = 14'b00011001110110;
  assign mem[916] = 14'b10111100010101;
  assign mem[917] = 14'b01001101011000;
  assign mem[918] = 14'b10011110010110;
  assign mem[919] = 14'b01000100101010;
  assign mem[920] = 14'b01100111000000;
  assign mem[921] = 14'b01111011011010;
  assign mem[922] = 14'b01110101001001;
  assign mem[923] = 14'b10001011001000;
  assign mem[924] = 14'b10111011111101;
  assign mem[925] = 14'b00110111111101;
  assign mem[926] = 14'b10100111111100;
  assign mem[927] = 14'b01011000101010;
  assign mem[928] = 14'b10100001110110;
  assign mem[929] = 14'b01001100100101;
  assign mem[930] = 14'b01110011110110;
  assign mem[931] = 14'b10001001000011;
  assign mem[932] = 14'b00001011000110;
  assign mem[933] = 14'b01101001101100;
  assign mem[934] = 14'b10000100001110;
  assign mem[935] = 14'b01110000011001;
  assign mem[936] = 14'b01010011111011;
  assign mem[937] = 14'b01110001101010;
  assign mem[938] = 14'b10101101001100;
  assign mem[939] = 14'b00000100100010;
  assign mem[940] = 14'b01111010111000;
  assign mem[941] = 14'b01101010101011;
  assign mem[942] = 14'b10111000101110;
  assign mem[943] = 14'b00100111001101;
  assign mem[944] = 14'b01100110110010;
  assign mem[945] = 14'b00111110111010;
  assign mem[946] = 14'b01011010101111;
  assign mem[947] = 14'b00010110110010;
  assign mem[948] = 14'b01011001011001;
  assign mem[949] = 14'b01011010000010;
  assign mem[950] = 14'b01000001010010;
  assign mem[951] = 14'b00100000111001;
  assign mem[952] = 14'b10110101100101;
  assign mem[953] = 14'b01001011110100;
  assign mem[954] = 14'b10001011000001;
  assign mem[955] = 14'b00101100101000;
  assign mem[956] = 14'b10110011110110;
  assign mem[957] = 14'b10010000110000;
  assign mem[958] = 14'b00100111011000;
  assign mem[959] = 14'b10001001001000;
  assign mem[960] = 14'b01101101100011;
  assign mem[961] = 14'b00101001010111;
  assign mem[962] = 14'b00011101101010;
  assign mem[963] = 14'b01101101111111;
  assign mem[964] = 14'b01011100111110;
  assign mem[965] = 14'b10101110011011;
  assign mem[966] = 14'b01010101110000;
  assign mem[967] = 14'b01100010000101;
  assign mem[968] = 14'b10001111011110;
  assign mem[969] = 14'b10110011000000;
  assign mem[970] = 14'b00001001111001;
  assign mem[971] = 14'b10011100111110;
  assign mem[972] = 14'b10110100100010;
  assign mem[973] = 14'b01011000000001;
  assign mem[974] = 14'b10010101110011;
  assign mem[975] = 14'b00100100011101;
  assign mem[976] = 14'b01101101100000;
  assign mem[977] = 14'b01101110101100;
  assign mem[978] = 14'b01001110110111;
  assign mem[979] = 14'b01110000011111;
  assign mem[980] = 14'b10011010001001;
  assign mem[981] = 14'b10001100100101;
  assign mem[982] = 14'b00001000111001;
  assign mem[983] = 14'b01100011110110;
  assign mem[984] = 14'b10101001011101;
  assign mem[985] = 14'b10010111001111;
  assign mem[986] = 14'b10000001001100;
  assign mem[987] = 14'b10110011010000;
  assign mem[988] = 14'b01000001101011;
  assign mem[989] = 14'b00011111001101;
  assign mem[990] = 14'b00000000000010;
  assign mem[991] = 14'b10010001110011;
  assign mem[992] = 14'b00000010100010;
  assign mem[993] = 14'b01100000100110;
  assign mem[994] = 14'b00011111010000;
  assign mem[995] = 14'b00111001000001;
  assign mem[996] = 14'b10011001000000;
  assign mem[997] = 14'b01100011011011;
  assign mem[998] = 14'b01110110000101;
  assign mem[999] = 14'b01100000101011;
  assign mem[1000] = 14'b10000100111110;
  assign mem[1001] = 14'b10011011001111;
  assign mem[1002] = 14'b01010110100000;
  assign mem[1003] = 14'b10001100111011;
  assign mem[1004] = 14'b00111001111010;
  assign mem[1005] = 14'b10111011101001;
  assign mem[1006] = 14'b00010110101100;
  assign mem[1007] = 14'b00101111111011;
  assign mem[1008] = 14'b01010101110110;
  assign mem[1009] = 14'b10010111011100;
  assign mem[1010] = 14'b01001100000001;
  assign mem[1011] = 14'b01011110000011;
  assign mem[1012] = 14'b01101111000010;
  assign mem[1013] = 14'b10010110001010;
  assign mem[1014] = 14'b01000111101100;
  assign mem[1015] = 14'b10011110110101;
  assign mem[1016] = 14'b01100001110101;
  assign mem[1017] = 14'b01011011111111;
  assign mem[1018] = 14'b00101001011100;
  assign mem[1019] = 14'b10011110111100;
  assign mem[1020] = 14'b00011000101100;
  assign mem[1021] = 14'b10100010001011;
  assign mem[1022] = 14'b01001000011110;
  assign mem[1023] = 14'b10011011011101;
  always@(*)
  begin
    data_out_t <= mem[addr_f];
  end
  wire [13:0] data_out_reg [n_outreg:0];
  generate if (n_outreg > 0)
  begin
    for( i=n_outreg-1; i >= 1; i=i-1)
    begin: data_out_reg_stage
      mgc_generic_reg #(
        .width(14),
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_data_out_reg (
        .d(data_out_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(data_out_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(14),
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_data_out_reg_init (
      .d(data_out_t),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(data_out_reg[0])
    );
    assign data_out = data_out_reg[n_outreg-1];
  end
  else
  begin
    assign data_out = data_out_t;
  end
  endgenerate
endmodule
module stagemgc_rom_sync_regout_13_1024_14_1_0_0_1_0_1_0_0_0_1_60 (addr, data_out,
    clk, s_rst, a_rst, en
);
  input [9:0]addr ;
  output [13:0]data_out ;
  input clk ;
  input s_rst ;
  input a_rst ;
  input en ;
  parameter n_width = 14;
  parameter n_size = 1024;
  parameter n_numports = 1;
  parameter n_addr_w = 10;
  parameter n_inreg = 0;
  parameter n_outreg = 1;
  wire [9:0] addr_f;
  wire [9:0] addr_reg [n_inreg:0];
  genvar i;
  generate if (n_inreg > 0)
  begin
    for( i=n_inreg-1; i >= 1; i=i-1)
    begin: addr_reg_stage
      mgc_generic_reg #(
        .width(10),
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_addr_reg (
        .d(addr_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(addr_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(10),
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_addr_reg_init (
      .d(addr),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(addr_reg[0])
    );
    assign addr_f = addr_reg[n_inreg-1];
  end
  else
  begin
    assign addr_f = addr;
  end
  endgenerate
  wire [13:0] mem [1023:0];
  reg [13:0] data_out_t;
  assign mem[0] = 14'b00111111111011;
  assign mem[1] = 14'b01000100110001;
  assign mem[2] = 14'b00010000111001;
  assign mem[3] = 14'b00010011001101;
  assign mem[4] = 14'b00100111100010;
  assign mem[5] = 14'b01011101111110;
  assign mem[6] = 14'b01111100001011;
  assign mem[7] = 14'b01010011010001;
  assign mem[8] = 14'b00101000010011;
  assign mem[9] = 14'b01001010001111;
  assign mem[10] = 14'b01100101000000;
  assign mem[11] = 14'b10110110110111;
  assign mem[12] = 14'b01101101101111;
  assign mem[13] = 14'b00101011111100;
  assign mem[14] = 14'b01011100000010;
  assign mem[15] = 14'b10100111001010;
  assign mem[16] = 14'b00110000100101;
  assign mem[17] = 14'b00100001001101;
  assign mem[18] = 14'b00011110101000;
  assign mem[19] = 14'b10101010101101;
  assign mem[20] = 14'b10100101101001;
  assign mem[21] = 14'b10100010100100;
  assign mem[22] = 14'b01000001011101;
  assign mem[23] = 14'b00011101010011;
  assign mem[24] = 14'b01011011010111;
  assign mem[25] = 14'b10000101100010;
  assign mem[26] = 14'b01001000000111;
  assign mem[27] = 14'b01010001000110;
  assign mem[28] = 14'b10110000111100;
  assign mem[29] = 14'b10100101010010;
  assign mem[30] = 14'b01011011111010;
  assign mem[31] = 14'b10101110010011;
  assign mem[32] = 14'b10000011100001;
  assign mem[33] = 14'b10111111110011;
  assign mem[34] = 14'b10100101100111;
  assign mem[35] = 14'b01110100010110;
  assign mem[36] = 14'b01011001010111;
  assign mem[37] = 14'b00110111110001;
  assign mem[38] = 14'b01011101011101;
  assign mem[39] = 14'b10011101111100;
  assign mem[40] = 14'b01000101001010;
  assign mem[41] = 14'b10000001110010;
  assign mem[42] = 14'b10101000000011;
  assign mem[43] = 14'b01001001000111;
  assign mem[44] = 14'b10101100101100;
  assign mem[45] = 14'b00011000000010;
  assign mem[46] = 14'b10111001010001;
  assign mem[47] = 14'b00000001100100;
  assign mem[48] = 14'b10000000110111;
  assign mem[49] = 14'b01100111100001;
  assign mem[50] = 14'b10010111111101;
  assign mem[51] = 14'b01010000011001;
  assign mem[52] = 14'b00110101010100;
  assign mem[53] = 14'b01111010110010;
  assign mem[54] = 14'b01011011000111;
  assign mem[55] = 14'b10010011110100;
  assign mem[56] = 14'b01010001100001;
  assign mem[57] = 14'b10100111110100;
  assign mem[58] = 14'b01111011001010;
  assign mem[59] = 14'b01110101010010;
  assign mem[60] = 14'b10111110001100;
  assign mem[61] = 14'b10110000011100;
  assign mem[62] = 14'b01011110100001;
  assign mem[63] = 14'b00000001001111;
  assign mem[64] = 14'b00000000001101;
  assign mem[65] = 14'b01101100011010;
  assign mem[66] = 14'b10001010110110;
  assign mem[67] = 14'b01010101001101;
  assign mem[68] = 14'b01000111101010;
  assign mem[69] = 14'b10110010111111;
  assign mem[70] = 14'b00101101010111;
  assign mem[71] = 14'b01001001000100;
  assign mem[72] = 14'b10011001110011;
  assign mem[73] = 14'b01110111000101;
  assign mem[74] = 14'b10001001110110;
  assign mem[75] = 14'b10001110010101;
  assign mem[76] = 14'b00100000100011;
  assign mem[77] = 14'b10000100111011;
  assign mem[78] = 14'b10000111101101;
  assign mem[79] = 14'b00110000100110;
  assign mem[80] = 14'b01101101100111;
  assign mem[81] = 14'b00110011000101;
  assign mem[82] = 14'b00010101010111;
  assign mem[83] = 14'b01100011111101;
  assign mem[84] = 14'b10100000010011;
  assign mem[85] = 14'b10000011110011;
  assign mem[86] = 14'b10100100011111;
  assign mem[87] = 14'b10110100100111;
  assign mem[88] = 14'b10101101010110;
  assign mem[89] = 14'b00100010100011;
  assign mem[90] = 14'b00011100010000;
  assign mem[91] = 14'b01110010010111;
  assign mem[92] = 14'b00000000110000;
  assign mem[93] = 14'b10010101001011;
  assign mem[94] = 14'b00101000000000;
  assign mem[95] = 14'b00010011001100;
  assign mem[96] = 14'b10010011011110;
  assign mem[97] = 14'b10101000100011;
  assign mem[98] = 14'b10111000011000;
  assign mem[99] = 14'b00011100011100;
  assign mem[100] = 14'b10110010001110;
  assign mem[101] = 14'b10001100000110;
  assign mem[102] = 14'b01100000001111;
  assign mem[103] = 14'b00101111000100;
  assign mem[104] = 14'b01011111011101;
  assign mem[105] = 14'b00101011101100;
  assign mem[106] = 14'b00100010011011;
  assign mem[107] = 14'b00011001110100;
  assign mem[108] = 14'b00001011000111;
  assign mem[109] = 14'b01101101011100;
  assign mem[110] = 14'b00010000011101;
  assign mem[111] = 14'b10001100001101;
  assign mem[112] = 14'b01010001111100;
  assign mem[113] = 14'b00010111101101;
  assign mem[114] = 14'b10010001101010;
  assign mem[115] = 14'b10110000000101;
  assign mem[116] = 14'b00001110000100;
  assign mem[117] = 14'b00111100110000;
  assign mem[118] = 14'b10101101111101;
  assign mem[119] = 14'b10100111110000;
  assign mem[120] = 14'b01001101010101;
  assign mem[121] = 14'b01110111000000;
  assign mem[122] = 14'b10011011110110;
  assign mem[123] = 14'b01001010001010;
  assign mem[124] = 14'b10100000011110;
  assign mem[125] = 14'b00000001111110;
  assign mem[126] = 14'b00101101101001;
  assign mem[127] = 14'b01101001000000;
  assign mem[128] = 14'b01100111101011;
  assign mem[129] = 14'b01100110001111;
  assign mem[130] = 14'b00011000101110;
  assign mem[131] = 14'b01001100000100;
  assign mem[132] = 14'b00000000101010;
  assign mem[133] = 14'b00001010100001;
  assign mem[134] = 14'b00100011000000;
  assign mem[135] = 14'b01110000110011;
  assign mem[136] = 14'b00010100010000;
  assign mem[137] = 14'b10111011010101;
  assign mem[138] = 14'b01110111111011;
  assign mem[139] = 14'b10000110000010;
  assign mem[140] = 14'b10111010101101;
  assign mem[141] = 14'b00001111011101;
  assign mem[142] = 14'b10100100101101;
  assign mem[143] = 14'b01111000000111;
  assign mem[144] = 14'b01101110101101;
  assign mem[145] = 14'b10000100100111;
  assign mem[146] = 14'b00001111101100;
  assign mem[147] = 14'b10011111111100;
  assign mem[148] = 14'b01001001011111;
  assign mem[149] = 14'b00000010100011;
  assign mem[150] = 14'b10001110110111;
  assign mem[151] = 14'b01000111110101;
  assign mem[152] = 14'b01100100011111;
  assign mem[153] = 14'b10111100010100;
  assign mem[154] = 14'b00101110101111;
  assign mem[155] = 14'b10111010100010;
  assign mem[156] = 14'b01001000100111;
  assign mem[157] = 14'b00110100100010;
  assign mem[158] = 14'b00100000001100;
  assign mem[159] = 14'b10110001011101;
  assign mem[160] = 14'b10111011101011;
  assign mem[161] = 14'b01101000001000;
  assign mem[162] = 14'b01011000010111;
  assign mem[163] = 14'b01110000111001;
  assign mem[164] = 14'b01011100011010;
  assign mem[165] = 14'b10010001101111;
  assign mem[166] = 14'b00111111111100;
  assign mem[167] = 14'b01011011111000;
  assign mem[168] = 14'b01101100010100;
  assign mem[169] = 14'b00110101001010;
  assign mem[170] = 14'b01010000001101;
  assign mem[171] = 14'b10010010110010;
  assign mem[172] = 14'b10101111011101;
  assign mem[173] = 14'b01010010000100;
  assign mem[174] = 14'b10001100110000;
  assign mem[175] = 14'b00011000010100;
  assign mem[176] = 14'b01101011111100;
  assign mem[177] = 14'b01001010100101;
  assign mem[178] = 14'b00111100001101;
  assign mem[179] = 14'b10001001001100;
  assign mem[180] = 14'b10100001010101;
  assign mem[181] = 14'b01111000111001;
  assign mem[182] = 14'b00011011011110;
  assign mem[183] = 14'b01101110111111;
  assign mem[184] = 14'b10110001101111;
  assign mem[185] = 14'b10111111110001;
  assign mem[186] = 14'b10000110011010;
  assign mem[187] = 14'b00110010101011;
  assign mem[188] = 14'b01100110001000;
  assign mem[189] = 14'b01110110100110;
  assign mem[190] = 14'b10000110001111;
  assign mem[191] = 14'b10110100100000;
  assign mem[192] = 14'b01011111010101;
  assign mem[193] = 14'b00110010110101;
  assign mem[194] = 14'b10011011110001;
  assign mem[195] = 14'b10010110101000;
  assign mem[196] = 14'b01000110011010;
  assign mem[197] = 14'b00111010011000;
  assign mem[198] = 14'b01101010101101;
  assign mem[199] = 14'b10101001000110;
  assign mem[200] = 14'b10001110101010;
  assign mem[201] = 14'b10011011011100;
  assign mem[202] = 14'b00110111101110;
  assign mem[203] = 14'b00100001010101;
  assign mem[204] = 14'b00111100111101;
  assign mem[205] = 14'b01011110010110;
  assign mem[206] = 14'b01110010100101;
  assign mem[207] = 14'b01100111010001;
  assign mem[208] = 14'b00110110001100;
  assign mem[209] = 14'b01001000110011;
  assign mem[210] = 14'b00001001110001;
  assign mem[211] = 14'b00101010001100;
  assign mem[212] = 14'b01111000111010;
  assign mem[213] = 14'b00110101110011;
  assign mem[214] = 14'b00101111110100;
  assign mem[215] = 14'b00110100111100;
  assign mem[216] = 14'b00110111000110;
  assign mem[217] = 14'b01000101000010;
  assign mem[218] = 14'b10111010000111;
  assign mem[219] = 14'b01100001011000;
  assign mem[220] = 14'b00011011000010;
  assign mem[221] = 14'b00100111111110;
  assign mem[222] = 14'b10100001100100;
  assign mem[223] = 14'b01010011100000;
  assign mem[224] = 14'b01010010100110;
  assign mem[225] = 14'b00100010001110;
  assign mem[226] = 14'b10110100101010;
  assign mem[227] = 14'b01100000110111;
  assign mem[228] = 14'b00100110110010;
  assign mem[229] = 14'b10001000110100;
  assign mem[230] = 14'b01010100001011;
  assign mem[231] = 14'b01000000000101;
  assign mem[232] = 14'b01001000000001;
  assign mem[233] = 14'b10000110011101;
  assign mem[234] = 14'b10000000100010;
  assign mem[235] = 14'b00000010010000;
  assign mem[236] = 14'b01011000011000;
  assign mem[237] = 14'b10001000000000;
  assign mem[238] = 14'b00101000111101;
  assign mem[239] = 14'b01010100110000;
  assign mem[240] = 14'b10101000111100;
  assign mem[241] = 14'b00101110001111;
  assign mem[242] = 14'b10110001010010;
  assign mem[243] = 14'b01100001101001;
  assign mem[244] = 14'b00011010110011;
  assign mem[245] = 14'b01001101010111;
  assign mem[246] = 14'b10010101000100;
  assign mem[247] = 14'b00011101100000;
  assign mem[248] = 14'b00111010110100;
  assign mem[249] = 14'b00000000100111;
  assign mem[250] = 14'b10000000011011;
  assign mem[251] = 14'b00100000100000;
  assign mem[252] = 14'b00100111000110;
  assign mem[253] = 14'b00010110111101;
  assign mem[254] = 14'b10100100110110;
  assign mem[255] = 14'b10001000000101;
  assign mem[256] = 14'b01010111100001;
  assign mem[257] = 14'b00010001000101;
  assign mem[258] = 14'b00111011001000;
  assign mem[259] = 14'b01001110110001;
  assign mem[260] = 14'b00100000001010;
  assign mem[261] = 14'b10000011001111;
  assign mem[262] = 14'b10110010111000;
  assign mem[263] = 14'b10010110100111;
  assign mem[264] = 14'b00100000001011;
  assign mem[265] = 14'b10011010010110;
  assign mem[266] = 14'b01110011101101;
  assign mem[267] = 14'b00100111000000;
  assign mem[268] = 14'b01111011101110;
  assign mem[269] = 14'b10110101001010;
  assign mem[270] = 14'b00000101110011;
  assign mem[271] = 14'b01111100111001;
  assign mem[272] = 14'b00110000000001;
  assign mem[273] = 14'b10100001010110;
  assign mem[274] = 14'b00000000101000;
  assign mem[275] = 14'b10011100010100;
  assign mem[276] = 14'b10010000011101;
  assign mem[277] = 14'b01111100110011;
  assign mem[278] = 14'b01010111100011;
  assign mem[279] = 14'b00111111010011;
  assign mem[280] = 14'b01111011010110;
  assign mem[281] = 14'b00001010100100;
  assign mem[282] = 14'b10110001110100;
  assign mem[283] = 14'b01110011010011;
  assign mem[284] = 14'b01100101100101;
  assign mem[285] = 14'b01001101110101;
  assign mem[286] = 14'b00101001000100;
  assign mem[287] = 14'b00110110100000;
  assign mem[288] = 14'b10101011001100;
  assign mem[289] = 14'b01101101101110;
  assign mem[290] = 14'b01101001010001;
  assign mem[291] = 14'b10011011001101;
  assign mem[292] = 14'b01101111100011;
  assign mem[293] = 14'b00100100011010;
  assign mem[294] = 14'b00111100101100;
  assign mem[295] = 14'b01010101100001;
  assign mem[296] = 14'b01111010111001;
  assign mem[297] = 14'b01101100011101;
  assign mem[298] = 14'b01011001101001;
  assign mem[299] = 14'b01010111101101;
  assign mem[300] = 14'b10010100100001;
  assign mem[301] = 14'b10110100110000;
  assign mem[302] = 14'b10110000001101;
  assign mem[303] = 14'b00100111001110;
  assign mem[304] = 14'b01101000100001;
  assign mem[305] = 14'b00000110000010;
  assign mem[306] = 14'b01000101101110;
  assign mem[307] = 14'b00000001101001;
  assign mem[308] = 14'b00100000011100;
  assign mem[309] = 14'b10100011001011;
  assign mem[310] = 14'b00000001110111;
  assign mem[311] = 14'b00111101110011;
  assign mem[312] = 14'b01000100010010;
  assign mem[313] = 14'b10110011110001;
  assign mem[314] = 14'b00111001011000;
  assign mem[315] = 14'b10110010101111;
  assign mem[316] = 14'b00001011101110;
  assign mem[317] = 14'b00110010101000;
  assign mem[318] = 14'b00110000111101;
  assign mem[319] = 14'b00001011110010;
  assign mem[320] = 14'b00111110101101;
  assign mem[321] = 14'b10111010011001;
  assign mem[322] = 14'b10001111111010;
  assign mem[323] = 14'b01010100000010;
  assign mem[324] = 14'b10111001101001;
  assign mem[325] = 14'b10101100001010;
  assign mem[326] = 14'b00101100000010;
  assign mem[327] = 14'b00011100111011;
  assign mem[328] = 14'b01001101100110;
  assign mem[329] = 14'b01111111110101;
  assign mem[330] = 14'b00101010000000;
  assign mem[331] = 14'b01100000111101;
  assign mem[332] = 14'b01101010011110;
  assign mem[333] = 14'b00001110011110;
  assign mem[334] = 14'b00101101111000;
  assign mem[335] = 14'b01000011100111;
  assign mem[336] = 14'b10011110111111;
  assign mem[337] = 14'b01101110110001;
  assign mem[338] = 14'b01011110011111;
  assign mem[339] = 14'b10010011000010;
  assign mem[340] = 14'b10100011111100;
  assign mem[341] = 14'b10001011110110;
  assign mem[342] = 14'b00100110101000;
  assign mem[343] = 14'b01100001101111;
  assign mem[344] = 14'b00001011011000;
  assign mem[345] = 14'b01110110010001;
  assign mem[346] = 14'b01011110101000;
  assign mem[347] = 14'b10100011000000;
  assign mem[348] = 14'b10101100011100;
  assign mem[349] = 14'b00100110010100;
  assign mem[350] = 14'b00101011111011;
  assign mem[351] = 14'b00111011001011;
  assign mem[352] = 14'b00001110110001;
  assign mem[353] = 14'b10001100100110;
  assign mem[354] = 14'b00010011011100;
  assign mem[355] = 14'b10001001101111;
  assign mem[356] = 14'b10101100001001;
  assign mem[357] = 14'b10101111010010;
  assign mem[358] = 14'b01011100000110;
  assign mem[359] = 14'b01000011100101;
  assign mem[360] = 14'b01001000011111;
  assign mem[361] = 14'b00111011101011;
  assign mem[362] = 14'b10011001100010;
  assign mem[363] = 14'b01101110010000;
  assign mem[364] = 14'b01101010000010;
  assign mem[365] = 14'b10000111011110;
  assign mem[366] = 14'b01010110100011;
  assign mem[367] = 14'b01111000011011;
  assign mem[368] = 14'b00010101010001;
  assign mem[369] = 14'b10011001010100;
  assign mem[370] = 14'b00101110000101;
  assign mem[371] = 14'b10110000000001;
  assign mem[372] = 14'b10100000111101;
  assign mem[373] = 14'b10001110010100;
  assign mem[374] = 14'b00000111011110;
  assign mem[375] = 14'b01100101011001;
  assign mem[376] = 14'b00000001100101;
  assign mem[377] = 14'b00011101110111;
  assign mem[378] = 14'b10010100001011;
  assign mem[379] = 14'b00111000011000;
  assign mem[380] = 14'b10111011011101;
  assign mem[381] = 14'b10100100101000;
  assign mem[382] = 14'b00001100101100;
  assign mem[383] = 14'b10001011010011;
  assign mem[384] = 14'b00001001111101;
  assign mem[385] = 14'b01111111011111;
  assign mem[386] = 14'b01010010110011;
  assign mem[387] = 14'b10001110101000;
  assign mem[388] = 14'b00110110111000;
  assign mem[389] = 14'b10000001100010;
  assign mem[390] = 14'b01101110011100;
  assign mem[391] = 14'b01111011110010;
  assign mem[392] = 14'b00101111011100;
  assign mem[393] = 14'b01001010010111;
  assign mem[394] = 14'b00100001110011;
  assign mem[395] = 14'b00111101100001;
  assign mem[396] = 14'b00111010101011;
  assign mem[397] = 14'b10110000101010;
  assign mem[398] = 14'b01111000111011;
  assign mem[399] = 14'b01001100111010;
  assign mem[400] = 14'b10111010011100;
  assign mem[401] = 14'b00000110101000;
  assign mem[402] = 14'b01010110100010;
  assign mem[403] = 14'b01100001010100;
  assign mem[404] = 14'b10101101111011;
  assign mem[405] = 14'b01111001100010;
  assign mem[406] = 14'b10111011000110;
  assign mem[407] = 14'b00010001001001;
  assign mem[408] = 14'b00101101001010;
  assign mem[409] = 14'b10011100101011;
  assign mem[410] = 14'b00101000001001;
  assign mem[411] = 14'b00100011001010;
  assign mem[412] = 14'b00100100110000;
  assign mem[413] = 14'b00001100110101;
  assign mem[414] = 14'b00100111110110;
  assign mem[415] = 14'b10101100001000;
  assign mem[416] = 14'b01111001011001;
  assign mem[417] = 14'b00000010001000;
  assign mem[418] = 14'b00001001101001;
  assign mem[419] = 14'b00110001010101;
  assign mem[420] = 14'b01011100000001;
  assign mem[421] = 14'b10010000000011;
  assign mem[422] = 14'b01101011000111;
  assign mem[423] = 14'b00000001111000;
  assign mem[424] = 14'b01000100110101;
  assign mem[425] = 14'b00011100100001;
  assign mem[426] = 14'b10010110100011;
  assign mem[427] = 14'b01110000101110;
  assign mem[428] = 14'b10100000010101;
  assign mem[429] = 14'b10110010000001;
  assign mem[430] = 14'b00100110001001;
  assign mem[431] = 14'b10010101011010;
  assign mem[432] = 14'b10101110101000;
  assign mem[433] = 14'b00001001010111;
  assign mem[434] = 14'b00100000100101;
  assign mem[435] = 14'b10110011001001;
  assign mem[436] = 14'b01110001000001;
  assign mem[437] = 14'b01100000100001;
  assign mem[438] = 14'b01001011000001;
  assign mem[439] = 14'b10011011000110;
  assign mem[440] = 14'b10001100110010;
  assign mem[441] = 14'b01000110100010;
  assign mem[442] = 14'b10010011101111;
  assign mem[443] = 14'b10110001011000;
  assign mem[444] = 14'b10110110010110;
  assign mem[445] = 14'b01100000011110;
  assign mem[446] = 14'b01111100001110;
  assign mem[447] = 14'b10011000100110;
  assign mem[448] = 14'b01101011110000;
  assign mem[449] = 14'b10110101010011;
  assign mem[450] = 14'b00110010001101;
  assign mem[451] = 14'b10000100011001;
  assign mem[452] = 14'b10011010010001;
  assign mem[453] = 14'b00101100010011;
  assign mem[454] = 14'b10100010110110;
  assign mem[455] = 14'b00111010010100;
  assign mem[456] = 14'b01111100011001;
  assign mem[457] = 14'b00010110110001;
  assign mem[458] = 14'b10101001101001;
  assign mem[459] = 14'b01111110000101;
  assign mem[460] = 14'b00001101000000;
  assign mem[461] = 14'b00011001011100;
  assign mem[462] = 14'b00110101010010;
  assign mem[463] = 14'b01001100100100;
  assign mem[464] = 14'b10101001100111;
  assign mem[465] = 14'b01001111110111;
  assign mem[466] = 14'b10010101000111;
  assign mem[467] = 14'b01100010110101;
  assign mem[468] = 14'b01110100000111;
  assign mem[469] = 14'b00111111110011;
  assign mem[470] = 14'b00110000000000;
  assign mem[471] = 14'b10001010001111;
  assign mem[472] = 14'b10011001111101;
  assign mem[473] = 14'b10011110001010;
  assign mem[474] = 14'b01010010001011;
  assign mem[475] = 14'b10110010010101;
  assign mem[476] = 14'b01100110011100;
  assign mem[477] = 14'b00000100101111;
  assign mem[478] = 14'b00010110111001;
  assign mem[479] = 14'b00111100011111;
  assign mem[480] = 14'b01001100001001;
  assign mem[481] = 14'b01011010110101;
  assign mem[482] = 14'b10011100100001;
  assign mem[483] = 14'b01101011110010;
  assign mem[484] = 14'b00110011101111;
  assign mem[485] = 14'b01011100111011;
  assign mem[486] = 14'b10000110111101;
  assign mem[487] = 14'b01011011011100;
  assign mem[488] = 14'b00111100010000;
  assign mem[489] = 14'b00001110100000;
  assign mem[490] = 14'b01001101000101;
  assign mem[491] = 14'b10000101010010;
  assign mem[492] = 14'b00011101001111;
  assign mem[493] = 14'b00100010001000;
  assign mem[494] = 14'b01010111000011;
  assign mem[495] = 14'b01011011110111;
  assign mem[496] = 14'b00110110011001;
  assign mem[497] = 14'b10110101001101;
  assign mem[498] = 14'b10010100100111;
  assign mem[499] = 14'b01111111011001;
  assign mem[500] = 14'b00000000100011;
  assign mem[501] = 14'b00101000110001;
  assign mem[502] = 14'b01011101001011;
  assign mem[503] = 14'b01111110000000;
  assign mem[504] = 14'b00010000111000;
  assign mem[505] = 14'b10111100000111;
  assign mem[506] = 14'b10000011111100;
  assign mem[507] = 14'b00101111101100;
  assign mem[508] = 14'b00111011100101;
  assign mem[509] = 14'b10101100111001;
  assign mem[510] = 14'b01101001010000;
  assign mem[511] = 14'b10000100000110;
  assign mem[512] = 14'b00100100100100;
  assign mem[513] = 14'b01110111100011;
  assign mem[514] = 14'b00011101110110;
  assign mem[515] = 14'b10100111010101;
  assign mem[516] = 14'b00100001000101;
  assign mem[517] = 14'b10010110100101;
  assign mem[518] = 14'b01100100000010;
  assign mem[519] = 14'b01011110001100;
  assign mem[520] = 14'b00100001001100;
  assign mem[521] = 14'b01111000010101;
  assign mem[522] = 14'b00101001110111;
  assign mem[523] = 14'b01010000111111;
  assign mem[524] = 14'b01100001111110;
  assign mem[525] = 14'b01110100000000;
  assign mem[526] = 14'b00101000100101;
  assign mem[527] = 14'b01101010001011;
  assign mem[528] = 14'b10010000000110;
  assign mem[529] = 14'b10101001010101;
  assign mem[530] = 14'b00000100011000;
  assign mem[531] = 14'b10000110000111;
  assign mem[532] = 14'b00110011000110;
  assign mem[533] = 14'b01101001100001;
  assign mem[534] = 14'b00100100110010;
  assign mem[535] = 14'b00111011000011;
  assign mem[536] = 14'b01011111010110;
  assign mem[537] = 14'b01001001111100;
  assign mem[538] = 14'b01011100100110;
  assign mem[539] = 14'b00100111000001;
  assign mem[540] = 14'b10000111000000;
  assign mem[541] = 14'b10100000110001;
  assign mem[542] = 14'b01011111011011;
  assign mem[543] = 14'b10111101011111;
  assign mem[544] = 14'b00101110001110;
  assign mem[545] = 14'b10111111111111;
  assign mem[546] = 14'b10100000110100;
  assign mem[547] = 14'b01111110010110;
  assign mem[548] = 14'b00001100110001;
  assign mem[549] = 14'b00111110110101;
  assign mem[550] = 14'b00101000110010;
  assign mem[551] = 14'b00010110100100;
  assign mem[552] = 14'b01011100001011;
  assign mem[553] = 14'b10110111001000;
  assign mem[554] = 14'b00110011011100;
  assign mem[555] = 14'b00100101111000;
  assign mem[556] = 14'b01001111100010;
  assign mem[557] = 14'b01110001001010;
  assign mem[558] = 14'b01010001010101;
  assign mem[559] = 14'b01010010100001;
  assign mem[560] = 14'b10011011100100;
  assign mem[561] = 14'b00101010001110;
  assign mem[562] = 14'b01101000000000;
  assign mem[563] = 14'b00001011011111;
  assign mem[564] = 14'b00100011000011;
  assign mem[565] = 14'b10110110001000;
  assign mem[566] = 14'b00001101000001;
  assign mem[567] = 14'b00110000100011;
  assign mem[568] = 14'b01011101111100;
  assign mem[569] = 14'b01101010010001;
  assign mem[570] = 14'b00010001100110;
  assign mem[571] = 14'b01100011000011;
  assign mem[572] = 14'b01010010000010;
  assign mem[573] = 14'b10100010010111;
  assign mem[574] = 14'b10010110101010;
  assign mem[575] = 14'b01010010011110;
  assign mem[576] = 14'b00110110111001;
  assign mem[577] = 14'b10011000101001;
  assign mem[578] = 14'b00101111010001;
  assign mem[579] = 14'b00001100001011;
  assign mem[580] = 14'b10010011011001;
  assign mem[581] = 14'b00110101000000;
  assign mem[582] = 14'b01110100001101;
  assign mem[583] = 14'b00001010011100;
  assign mem[584] = 14'b10011111001000;
  assign mem[585] = 14'b01111110101111;
  assign mem[586] = 14'b01100101111111;
  assign mem[587] = 14'b01100110101000;
  assign mem[588] = 14'b10101001001111;
  assign mem[589] = 14'b01100101010010;
  assign mem[590] = 14'b10000001000111;
  assign mem[591] = 14'b01011001001111;
  assign mem[592] = 14'b10011000110100;
  assign mem[593] = 14'b00000111010011;
  assign mem[594] = 14'b01010101010110;
  assign mem[595] = 14'b01000101001001;
  assign mem[596] = 14'b10111011011111;
  assign mem[597] = 14'b00010010110101;
  assign mem[598] = 14'b01001110010111;
  assign mem[599] = 14'b01101100000110;
  assign mem[600] = 14'b01001111101000;
  assign mem[601] = 14'b00111011110011;
  assign mem[602] = 14'b01010110010101;
  assign mem[603] = 14'b10110100111011;
  assign mem[604] = 14'b00110110111110;
  assign mem[605] = 14'b01001100001011;
  assign mem[606] = 14'b01110011011100;
  assign mem[607] = 14'b00011110001011;
  assign mem[608] = 14'b01100111010111;
  assign mem[609] = 14'b00011000000101;
  assign mem[610] = 14'b10001000000100;
  assign mem[611] = 14'b00000100000100;
  assign mem[612] = 14'b00110100111001;
  assign mem[613] = 14'b01001010111000;
  assign mem[614] = 14'b01000100100111;
  assign mem[615] = 14'b01011001000001;
  assign mem[616] = 14'b01111011010111;
  assign mem[617] = 14'b00100001101011;
  assign mem[618] = 14'b01110010101001;
  assign mem[619] = 14'b00000011101100;
  assign mem[620] = 14'b10100110001011;
  assign mem[621] = 14'b10110100001110;
  assign mem[622] = 14'b00011101110010;
  assign mem[623] = 14'b01001010111001;
  assign mem[624] = 14'b10010100110111;
  assign mem[625] = 14'b01110001000111;
  assign mem[626] = 14'b10000010100010;
  assign mem[627] = 14'b01010000000001;
  assign mem[628] = 14'b10100110100110;
  assign mem[629] = 14'b00100100000111;
  assign mem[630] = 14'b00110100010010;
  assign mem[631] = 14'b10000101101100;
  assign mem[632] = 14'b00001011000011;
  assign mem[633] = 14'b00010001000000;
  assign mem[634] = 14'b01001101001000;
  assign mem[635] = 14'b00001010100110;
  assign mem[636] = 14'b10100000000101;
  assign mem[637] = 14'b00000000010010;
  assign mem[638] = 14'b01011000110100;
  assign mem[639] = 14'b00001111000000;
  assign mem[640] = 14'b01000101101011;
  assign mem[641] = 14'b01111100010101;
  assign mem[642] = 14'b00000011100010;
  assign mem[643] = 14'b00100110010011;
  assign mem[644] = 14'b00000000000110;
  assign mem[645] = 14'b10001010101010;
  assign mem[646] = 14'b00000101000000;
  assign mem[647] = 14'b01100010011010;
  assign mem[648] = 14'b10001100000011;
  assign mem[649] = 14'b10001000011111;
  assign mem[650] = 14'b00101100100100;
  assign mem[651] = 14'b00101110100101;
  assign mem[652] = 14'b00011010101011;
  assign mem[653] = 14'b01010100100000;
  assign mem[654] = 14'b01001110011001;
  assign mem[655] = 14'b10011010010100;
  assign mem[656] = 14'b10011000111110;
  assign mem[657] = 14'b00101110011000;
  assign mem[658] = 14'b00011101101011;
  assign mem[659] = 14'b01101001001001;
  assign mem[660] = 14'b01000001010111;
  assign mem[661] = 14'b01010010101010;
  assign mem[662] = 14'b10011101100100;
  assign mem[663] = 14'b01110111111111;
  assign mem[664] = 14'b01111100000101;
  assign mem[665] = 14'b10001000101000;
  assign mem[666] = 14'b01011000111110;
  assign mem[667] = 14'b00110110000101;
  assign mem[668] = 14'b01000001001111;
  assign mem[669] = 14'b01011001110011;
  assign mem[670] = 14'b01010110111001;
  assign mem[671] = 14'b00110100110010;
  assign mem[672] = 14'b01010001101011;
  assign mem[673] = 14'b00001110111000;
  assign mem[674] = 14'b01000011011111;
  assign mem[675] = 14'b10011001010010;
  assign mem[676] = 14'b01000100000100;
  assign mem[677] = 14'b00110000010000;
  assign mem[678] = 14'b10101101101110;
  assign mem[679] = 14'b00001101001000;
  assign mem[680] = 14'b01100001110001;
  assign mem[681] = 14'b00000111100110;
  assign mem[682] = 14'b01011101110000;
  assign mem[683] = 14'b00010100111110;
  assign mem[684] = 14'b10100010001110;
  assign mem[685] = 14'b01011110000001;
  assign mem[686] = 14'b01001010111110;
  assign mem[687] = 14'b01010101110001;
  assign mem[688] = 14'b01000110010010;
  assign mem[689] = 14'b01000001100001;
  assign mem[690] = 14'b00100100000010;
  assign mem[691] = 14'b01100101111001;
  assign mem[692] = 14'b00010111000011;
  assign mem[693] = 14'b01100011100100;
  assign mem[694] = 14'b10001101000101;
  assign mem[695] = 14'b01111101100101;
  assign mem[696] = 14'b00011001011001;
  assign mem[697] = 14'b01101101101100;
  assign mem[698] = 14'b01001010000100;
  assign mem[699] = 14'b01011001100010;
  assign mem[700] = 14'b01111100010100;
  assign mem[701] = 14'b01100011001111;
  assign mem[702] = 14'b01100101011110;
  assign mem[703] = 14'b01101100000101;
  assign mem[704] = 14'b10110010001101;
  assign mem[705] = 14'b01110100111111;
  assign mem[706] = 14'b10011111011010;
  assign mem[707] = 14'b10011110101011;
  assign mem[708] = 14'b01110111110010;
  assign mem[709] = 14'b01110110000100;
  assign mem[710] = 14'b10110011110101;
  assign mem[711] = 14'b00011000001010;
  assign mem[712] = 14'b01100110101011;
  assign mem[713] = 14'b10011111010111;
  assign mem[714] = 14'b00100011011001;
  assign mem[715] = 14'b01110010011111;
  assign mem[716] = 14'b01011011000000;
  assign mem[717] = 14'b10110010000100;
  assign mem[718] = 14'b10110100111101;
  assign mem[719] = 14'b10010111111010;
  assign mem[720] = 14'b00100011001011;
  assign mem[721] = 14'b10101110111111;
  assign mem[722] = 14'b01010011101100;
  assign mem[723] = 14'b01110011110000;
  assign mem[724] = 14'b00101100101101;
  assign mem[725] = 14'b00111110100011;
  assign mem[726] = 14'b10001111111111;
  assign mem[727] = 14'b00000111100100;
  assign mem[728] = 14'b01110101100110;
  assign mem[729] = 14'b10010011000001;
  assign mem[730] = 14'b10111111001011;
  assign mem[731] = 14'b01100000001101;
  assign mem[732] = 14'b10001101000001;
  assign mem[733] = 14'b00100001001001;
  assign mem[734] = 14'b10100000001111;
  assign mem[735] = 14'b00100111010111;
  assign mem[736] = 14'b10010100111101;
  assign mem[737] = 14'b00111011110000;
  assign mem[738] = 14'b10000111100010;
  assign mem[739] = 14'b10110010011011;
  assign mem[740] = 14'b10101010001000;
  assign mem[741] = 14'b01001010011010;
  assign mem[742] = 14'b10110000100111;
  assign mem[743] = 14'b01000000000001;
  assign mem[744] = 14'b00100101101110;
  assign mem[745] = 14'b01100101100000;
  assign mem[746] = 14'b10011011100001;
  assign mem[747] = 14'b10100100111010;
  assign mem[748] = 14'b00001100101000;
  assign mem[749] = 14'b00101110110111;
  assign mem[750] = 14'b00100001010010;
  assign mem[751] = 14'b01000010111110;
  assign mem[752] = 14'b10111100101110;
  assign mem[753] = 14'b01110100010101;
  assign mem[754] = 14'b01010000001100;
  assign mem[755] = 14'b01111011101011;
  assign mem[756] = 14'b00000011110101;
  assign mem[757] = 14'b01011101010110;
  assign mem[758] = 14'b01001100001010;
  assign mem[759] = 14'b01110001111100;
  assign mem[760] = 14'b01110110001000;
  assign mem[761] = 14'b10100100101011;
  assign mem[762] = 14'b10011011100000;
  assign mem[763] = 14'b10001101110011;
  assign mem[764] = 14'b00100001000001;
  assign mem[765] = 14'b00111010001001;
  assign mem[766] = 14'b10100000101101;
  assign mem[767] = 14'b10011100100110;
  assign mem[768] = 14'b10010101101010;
  assign mem[769] = 14'b10001011100110;
  assign mem[770] = 14'b10101101000010;
  assign mem[771] = 14'b10010100011010;
  assign mem[772] = 14'b00000100100110;
  assign mem[773] = 14'b01001001100111;
  assign mem[774] = 14'b00110100111111;
  assign mem[775] = 14'b00010101100001;
  assign mem[776] = 14'b10001101110000;
  assign mem[777] = 14'b10011111001101;
  assign mem[778] = 14'b01000111011001;
  assign mem[779] = 14'b10101010001010;
  assign mem[780] = 14'b10011010110101;
  assign mem[781] = 14'b01101100001011;
  assign mem[782] = 14'b00000000110101;
  assign mem[783] = 14'b01001000101101;
  assign mem[784] = 14'b00000110110111;
  assign mem[785] = 14'b10100000001101;
  assign mem[786] = 14'b01101101110100;
  assign mem[787] = 14'b10011111011111;
  assign mem[788] = 14'b10000010010111;
  assign mem[789] = 14'b00010001110101;
  assign mem[790] = 14'b00100111111100;
  assign mem[791] = 14'b01110110110001;
  assign mem[792] = 14'b01111111010110;
  assign mem[793] = 14'b10100110000110;
  assign mem[794] = 14'b10000111001000;
  assign mem[795] = 14'b10011001101000;
  assign mem[796] = 14'b01111100001111;
  assign mem[797] = 14'b10101111101101;
  assign mem[798] = 14'b00100001010011;
  assign mem[799] = 14'b01011010000101;
  assign mem[800] = 14'b10100001100111;
  assign mem[801] = 14'b10011000110101;
  assign mem[802] = 14'b00101010011110;
  assign mem[803] = 14'b00010110001011;
  assign mem[804] = 14'b01000110110011;
  assign mem[805] = 14'b00111100000100;
  assign mem[806] = 14'b00111111100010;
  assign mem[807] = 14'b01000011000101;
  assign mem[808] = 14'b10110110001001;
  assign mem[809] = 14'b10110100000101;
  assign mem[810] = 14'b10110001011001;
  assign mem[811] = 14'b01000011011001;
  assign mem[812] = 14'b01001100000101;
  assign mem[813] = 14'b10111110011010;
  assign mem[814] = 14'b00011001001011;
  assign mem[815] = 14'b10101010001100;
  assign mem[816] = 14'b10110011100001;
  assign mem[817] = 14'b10001010000001;
  assign mem[818] = 14'b00100101011001;
  assign mem[819] = 14'b00000000001111;
  assign mem[820] = 14'b10101001001110;
  assign mem[821] = 14'b01001110001011;
  assign mem[822] = 14'b00000000010001;
  assign mem[823] = 14'b00001000110101;
  assign mem[824] = 14'b01011100000011;
  assign mem[825] = 14'b10111110010001;
  assign mem[826] = 14'b10101100110010;
  assign mem[827] = 14'b10100010101100;
  assign mem[828] = 14'b10001010110101;
  assign mem[829] = 14'b00111110000110;
  assign mem[830] = 14'b10101011100101;
  assign mem[831] = 14'b01101111011010;
  assign mem[832] = 14'b01011011010000;
  assign mem[833] = 14'b10100011110010;
  assign mem[834] = 14'b10000010010010;
  assign mem[835] = 14'b01011110010011;
  assign mem[836] = 14'b01101100110100;
  assign mem[837] = 14'b00011000100110;
  assign mem[838] = 14'b10101010111000;
  assign mem[839] = 14'b00011111100100;
  assign mem[840] = 14'b00100110100001;
  assign mem[841] = 14'b01111111111111;
  assign mem[842] = 14'b00000110000000;
  assign mem[843] = 14'b00101001010010;
  assign mem[844] = 14'b00101010101001;
  assign mem[845] = 14'b01010100010111;
  assign mem[846] = 14'b00100001111111;
  assign mem[847] = 14'b10010010110100;
  assign mem[848] = 14'b10111011010011;
  assign mem[849] = 14'b01111101100011;
  assign mem[850] = 14'b01000100010111;
  assign mem[851] = 14'b01100111010011;
  assign mem[852] = 14'b01001110010010;
  assign mem[853] = 14'b10111000100100;
  assign mem[854] = 14'b10001110101011;
  assign mem[855] = 14'b10110010100011;
  assign mem[856] = 14'b00000001101000;
  assign mem[857] = 14'b01100011001100;
  assign mem[858] = 14'b10010110101011;
  assign mem[859] = 14'b01101001100101;
  assign mem[860] = 14'b10111101001110;
  assign mem[861] = 14'b01010111110001;
  assign mem[862] = 14'b10101010110111;
  assign mem[863] = 14'b00001000011101;
  assign mem[864] = 14'b00000010000111;
  assign mem[865] = 14'b00101111100001;
  assign mem[866] = 14'b01110000100000;
  assign mem[867] = 14'b01100101111110;
  assign mem[868] = 14'b01001111011101;
  assign mem[869] = 14'b10111101101000;
  assign mem[870] = 14'b00001101001010;
  assign mem[871] = 14'b01000000100001;
  assign mem[872] = 14'b01111000000101;
  assign mem[873] = 14'b10101101000111;
  assign mem[874] = 14'b10000011101010;
  assign mem[875] = 14'b00001111110000;
  assign mem[876] = 14'b00101010100101;
  assign mem[877] = 14'b10110111111100;
  assign mem[878] = 14'b01011110101010;
  assign mem[879] = 14'b00010001001101;
  assign mem[880] = 14'b00011110011110;
  assign mem[881] = 14'b10000011101000;
  assign mem[882] = 14'b01011000111000;
  assign mem[883] = 14'b01101011011100;
  assign mem[884] = 14'b10111011100101;
  assign mem[885] = 14'b10011101011111;
  assign mem[886] = 14'b01010011010111;
  assign mem[887] = 14'b00001110011111;
  assign mem[888] = 14'b00011011101010;
  assign mem[889] = 14'b00000100010001;
  assign mem[890] = 14'b10000010111001;
  assign mem[891] = 14'b00100011011111;
  assign mem[892] = 14'b01010001101001;
  assign mem[893] = 14'b10100000101011;
  assign mem[894] = 14'b00000001110100;
  assign mem[895] = 14'b10111000011111;
  assign mem[896] = 14'b00000001011011;
  assign mem[897] = 14'b10110110110011;
  assign mem[898] = 14'b00001011110101;
  assign mem[899] = 14'b00010100011000;
  assign mem[900] = 14'b01110101100100;
  assign mem[901] = 14'b01100100110011;
  assign mem[902] = 14'b01111101100000;
  assign mem[903] = 14'b01111111011010;
  assign mem[904] = 14'b01110100100000;
  assign mem[905] = 14'b01000001011111;
  assign mem[906] = 14'b00000100110101;
  assign mem[907] = 14'b00100100001110;
  assign mem[908] = 14'b00100011110100;
  assign mem[909] = 14'b10100010011001;
  assign mem[910] = 14'b10110101110111;
  assign mem[911] = 14'b10010100001001;
  assign mem[912] = 14'b10111111001110;
  assign mem[913] = 14'b10100101100010;
  assign mem[914] = 14'b10010101100001;
  assign mem[915] = 14'b01111011101000;
  assign mem[916] = 14'b10100010000000;
  assign mem[917] = 14'b10011010100001;
  assign mem[918] = 14'b10111111010100;
  assign mem[919] = 14'b01110000001011;
  assign mem[920] = 14'b00111101010100;
  assign mem[921] = 14'b00110001110100;
  assign mem[922] = 14'b00000101101111;
  assign mem[923] = 14'b00100000011101;
  assign mem[924] = 14'b00000101010000;
  assign mem[925] = 14'b01010100001000;
  assign mem[926] = 14'b01010111111111;
  assign mem[927] = 14'b10000110010100;
  assign mem[928] = 14'b01001000001101;
  assign mem[929] = 14'b00011011101111;
  assign mem[930] = 14'b10001010100010;
  assign mem[931] = 14'b00000111000011;
  assign mem[932] = 14'b01011111011100;
  assign mem[933] = 14'b00010100100101;
  assign mem[934] = 14'b01100001100110;
  assign mem[935] = 14'b10001001011011;
  assign mem[936] = 14'b01011100001000;
  assign mem[937] = 14'b01110001110011;
  assign mem[938] = 14'b00110000111100;
  assign mem[939] = 14'b10110100101100;
  assign mem[940] = 14'b01001101110001;
  assign mem[941] = 14'b10111110000001;
  assign mem[942] = 14'b01110011001011;
  assign mem[943] = 14'b00010101010110;
  assign mem[944] = 14'b10111101100010;
  assign mem[945] = 14'b10100101111011;
  assign mem[946] = 14'b00111011100001;
  assign mem[947] = 14'b01010000011101;
  assign mem[948] = 14'b01100010011100;
  assign mem[949] = 14'b00101001001110;
  assign mem[950] = 14'b01000001100101;
  assign mem[951] = 14'b00010110001010;
  assign mem[952] = 14'b10011101010001;
  assign mem[953] = 14'b01000000111100;
  assign mem[954] = 14'b10000010110101;
  assign mem[955] = 14'b10000111000100;
  assign mem[956] = 14'b10100011001101;
  assign mem[957] = 14'b00001101110010;
  assign mem[958] = 14'b01111111011110;
  assign mem[959] = 14'b10011110111101;
  assign mem[960] = 14'b10011000100011;
  assign mem[961] = 14'b10111110011111;
  assign mem[962] = 14'b00000111001011;
  assign mem[963] = 14'b00101110010110;
  assign mem[964] = 14'b00110001011110;
  assign mem[965] = 14'b00000110010101;
  assign mem[966] = 14'b01001110001000;
  assign mem[967] = 14'b10010001011111;
  assign mem[968] = 14'b01100100000100;
  assign mem[969] = 14'b10001100011010;
  assign mem[970] = 14'b00011000001111;
  assign mem[971] = 14'b01111111101111;
  assign mem[972] = 14'b00111000101110;
  assign mem[973] = 14'b10101000001110;
  assign mem[974] = 14'b10010000110001;
  assign mem[975] = 14'b00001010111100;
  assign mem[976] = 14'b10000101111101;
  assign mem[977] = 14'b10010100100100;
  assign mem[978] = 14'b01100111100110;
  assign mem[979] = 14'b10110010101101;
  assign mem[980] = 14'b10110101001011;
  assign mem[981] = 14'b01011011011010;
  assign mem[982] = 14'b00111101101110;
  assign mem[983] = 14'b01001010100111;
  assign mem[984] = 14'b10111010100101;
  assign mem[985] = 14'b00010110100110;
  assign mem[986] = 14'b01011110000010;
  assign mem[987] = 14'b00110100111010;
  assign mem[988] = 14'b10110011001110;
  assign mem[989] = 14'b01010010111110;
  assign mem[990] = 14'b01010101100100;
  assign mem[991] = 14'b00001000101001;
  assign mem[992] = 14'b10010100000010;
  assign mem[993] = 14'b00101000011010;
  assign mem[994] = 14'b00010110010111;
  assign mem[995] = 14'b00101010110101;
  assign mem[996] = 14'b00000111011001;
  assign mem[997] = 14'b10110001110111;
  assign mem[998] = 14'b01001010001001;
  assign mem[999] = 14'b00001101000100;
  assign mem[1000] = 14'b00111111011110;
  assign mem[1001] = 14'b10100110101010;
  assign mem[1002] = 14'b01111000101111;
  assign mem[1003] = 14'b10110111101000;
  assign mem[1004] = 14'b01010110011110;
  assign mem[1005] = 14'b00000100111000;
  assign mem[1006] = 14'b01000011010011;
  assign mem[1007] = 14'b01000011111111;
  assign mem[1008] = 14'b01011010000100;
  assign mem[1009] = 14'b10000111100111;
  assign mem[1010] = 14'b10000010111101;
  assign mem[1011] = 14'b01111111111011;
  assign mem[1012] = 14'b00000000000101;
  assign mem[1013] = 14'b01110011100011;
  assign mem[1014] = 14'b01000100001011;
  assign mem[1015] = 14'b00010010000000;
  assign mem[1016] = 14'b01010100101101;
  assign mem[1017] = 14'b01010001101111;
  assign mem[1018] = 14'b01100101001001;
  assign mem[1019] = 14'b00000110110100;
  assign mem[1020] = 14'b01110110001111;
  assign mem[1021] = 14'b10000110011011;
  assign mem[1022] = 14'b01100001010101;
  assign mem[1023] = 14'b10000000100110;
  always@(*)
  begin
    data_out_t <= mem[addr_f];
  end
  wire [13:0] data_out_reg [n_outreg:0];
  generate if (n_outreg > 0)
  begin
    for( i=n_outreg-1; i >= 1; i=i-1)
    begin: data_out_reg_stage
      mgc_generic_reg #(
        .width(14),
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_data_out_reg (
        .d(data_out_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(data_out_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(14),
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_data_out_reg_init (
      .d(data_out_t),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(data_out_reg[0])
    );
    assign data_out = data_out_reg[n_outreg-1];
  end
  else
  begin
    assign data_out = data_out_t;
  end
  endgenerate
endmodule
module stagemgc_rom_sync_regout_12_1024_14_1_0_0_1_0_1_0_0_0_1_60 (addr, data_out,
    clk, s_rst, a_rst, en
);
  input [9:0]addr ;
  output [13:0]data_out ;
  input clk ;
  input s_rst ;
  input a_rst ;
  input en ;
  parameter n_width = 14;
  parameter n_size = 1024;
  parameter n_numports = 1;
  parameter n_addr_w = 10;
  parameter n_inreg = 0;
  parameter n_outreg = 1;
  wire [9:0] addr_f;
  wire [9:0] addr_reg [n_inreg:0];
  genvar i;
  generate if (n_inreg > 0)
  begin
    for( i=n_inreg-1; i >= 1; i=i-1)
    begin: addr_reg_stage
      mgc_generic_reg #(
        .width(10),
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_addr_reg (
        .d(addr_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(addr_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(10),
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_addr_reg_init (
      .d(addr),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(addr_reg[0])
    );
    assign addr_f = addr_reg[n_inreg-1];
  end
  else
  begin
    assign addr_f = addr;
  end
  endgenerate
  wire [13:0] mem [1023:0];
  reg [13:0] data_out_t;
  assign mem[0] = 14'b00111111111011;
  assign mem[1] = 14'b01111011010000;
  assign mem[2] = 14'b10101100110100;
  assign mem[3] = 14'b10101111001000;
  assign mem[4] = 14'b01101100110000;
  assign mem[5] = 14'b01000011110110;
  assign mem[6] = 14'b01100010000011;
  assign mem[7] = 14'b10011000011111;
  assign mem[8] = 14'b00011000110111;
  assign mem[9] = 14'b01100011111111;
  assign mem[10] = 14'b10010100000101;
  assign mem[11] = 14'b01010010010010;
  assign mem[12] = 14'b00001001001010;
  assign mem[13] = 14'b01011011000001;
  assign mem[14] = 14'b01110101110010;
  assign mem[15] = 14'b10010111101110;
  assign mem[16] = 14'b00010001101110;
  assign mem[17] = 14'b01100100000111;
  assign mem[18] = 14'b00011010101111;
  assign mem[19] = 14'b00001111000101;
  assign mem[20] = 14'b01101110111011;
  assign mem[21] = 14'b01110111111010;
  assign mem[22] = 14'b00111010011111;
  assign mem[23] = 14'b01100100101010;
  assign mem[24] = 14'b10100010101110;
  assign mem[25] = 14'b01111110100100;
  assign mem[26] = 14'b00011101011101;
  assign mem[27] = 14'b00011010011000;
  assign mem[28] = 14'b00010101010100;
  assign mem[29] = 14'b10100001011001;
  assign mem[30] = 14'b10011110110100;
  assign mem[31] = 14'b10001111011100;
  assign mem[32] = 14'b10111110110010;
  assign mem[33] = 14'b01100001100000;
  assign mem[34] = 14'b00001111100101;
  assign mem[35] = 14'b00000001110101;
  assign mem[36] = 14'b01001010101111;
  assign mem[37] = 14'b01000100110111;
  assign mem[38] = 14'b00011000001101;
  assign mem[39] = 14'b01101110100000;
  assign mem[40] = 14'b00101100001101;
  assign mem[41] = 14'b01100100111010;
  assign mem[42] = 14'b01000101001111;
  assign mem[43] = 14'b10001010101101;
  assign mem[44] = 14'b01101111101000;
  assign mem[45] = 14'b00101000000100;
  assign mem[46] = 14'b01011000100000;
  assign mem[47] = 14'b00111111001010;
  assign mem[48] = 14'b10111110011101;
  assign mem[49] = 14'b00000110110000;
  assign mem[50] = 14'b10100111111111;
  assign mem[51] = 14'b00010011010101;
  assign mem[52] = 14'b01110110111010;
  assign mem[53] = 14'b00010111111110;
  assign mem[54] = 14'b00111110001111;
  assign mem[55] = 14'b01111010110111;
  assign mem[56] = 14'b00100010000101;
  assign mem[57] = 14'b01100010100100;
  assign mem[58] = 14'b10001000010000;
  assign mem[59] = 14'b01100110101010;
  assign mem[60] = 14'b01001011101011;
  assign mem[61] = 14'b00011010011010;
  assign mem[62] = 14'b00000000001110;
  assign mem[63] = 14'b00111100100000;
  assign mem[64] = 14'b01010111000001;
  assign mem[65] = 14'b10010010011000;
  assign mem[66] = 14'b10111110000011;
  assign mem[67] = 14'b00011111100011;
  assign mem[68] = 14'b01110101110111;
  assign mem[69] = 14'b00100100001011;
  assign mem[70] = 14'b01001001000001;
  assign mem[71] = 14'b01110010101100;
  assign mem[72] = 14'b00011000010001;
  assign mem[73] = 14'b00010010000100;
  assign mem[74] = 14'b10000011010001;
  assign mem[75] = 14'b10110001111101;
  assign mem[76] = 14'b00001111111100;
  assign mem[77] = 14'b00101110010111;
  assign mem[78] = 14'b10101000010100;
  assign mem[79] = 14'b01101110000101;
  assign mem[80] = 14'b00110011110100;
  assign mem[81] = 14'b10101111100100;
  assign mem[82] = 14'b01010010100101;
  assign mem[83] = 14'b10110100111010;
  assign mem[84] = 14'b10100110001101;
  assign mem[85] = 14'b10011101100110;
  assign mem[86] = 14'b10010100010101;
  assign mem[87] = 14'b01100000100100;
  assign mem[88] = 14'b10010000111101;
  assign mem[89] = 14'b01011111110010;
  assign mem[90] = 14'b00110011111011;
  assign mem[91] = 14'b00001101110011;
  assign mem[92] = 14'b10100011100101;
  assign mem[93] = 14'b00000111101001;
  assign mem[94] = 14'b00010111011110;
  assign mem[95] = 14'b00101100100011;
  assign mem[96] = 14'b10101100110101;
  assign mem[97] = 14'b10011000000001;
  assign mem[98] = 14'b00101010110110;
  assign mem[99] = 14'b10111111010001;
  assign mem[100] = 14'b01001101101010;
  assign mem[101] = 14'b10100011110001;
  assign mem[102] = 14'b10011101011110;
  assign mem[103] = 14'b00010010101011;
  assign mem[104] = 14'b00001011011010;
  assign mem[105] = 14'b00011011100010;
  assign mem[106] = 14'b00111100001110;
  assign mem[107] = 14'b00011111101110;
  assign mem[108] = 14'b01011100000100;
  assign mem[109] = 14'b10101010101010;
  assign mem[110] = 14'b10001100111100;
  assign mem[111] = 14'b01010010011010;
  assign mem[112] = 14'b10001111011011;
  assign mem[113] = 14'b00111000010100;
  assign mem[114] = 14'b00111011000110;
  assign mem[115] = 14'b10011111011110;
  assign mem[116] = 14'b00110001101100;
  assign mem[117] = 14'b00110110001011;
  assign mem[118] = 14'b01001000111100;
  assign mem[119] = 14'b00100110001110;
  assign mem[120] = 14'b01110110111101;
  assign mem[121] = 14'b10010010101010;
  assign mem[122] = 14'b00001101000010;
  assign mem[123] = 14'b01111000010111;
  assign mem[124] = 14'b01101010110100;
  assign mem[125] = 14'b00110101001011;
  assign mem[126] = 14'b01010011100111;
  assign mem[127] = 14'b10111111110100;
  assign mem[128] = 14'b00110111111100;
  assign mem[129] = 14'b00011011001011;
  assign mem[130] = 14'b10101001000100;
  assign mem[131] = 14'b10011000111011;
  assign mem[132] = 14'b10011111100001;
  assign mem[133] = 14'b00111111100110;
  assign mem[134] = 14'b10111111011010;
  assign mem[135] = 14'b10000101001101;
  assign mem[136] = 14'b10100010100001;
  assign mem[137] = 14'b00101010111101;
  assign mem[138] = 14'b01110010101010;
  assign mem[139] = 14'b10100101001110;
  assign mem[140] = 14'b01011110011000;
  assign mem[141] = 14'b00001110101111;
  assign mem[142] = 14'b10010001110010;
  assign mem[143] = 14'b00010111000101;
  assign mem[144] = 14'b01101011010001;
  assign mem[145] = 14'b10010111000100;
  assign mem[146] = 14'b00111000000001;
  assign mem[147] = 14'b01100111101001;
  assign mem[148] = 14'b10111101110001;
  assign mem[149] = 14'b00111111011111;
  assign mem[150] = 14'b00111001100100;
  assign mem[151] = 14'b01111000000000;
  assign mem[152] = 14'b01111111111100;
  assign mem[153] = 14'b01101011110110;
  assign mem[154] = 14'b00110111001101;
  assign mem[155] = 14'b10011001001111;
  assign mem[156] = 14'b01011111001010;
  assign mem[157] = 14'b00001011010111;
  assign mem[158] = 14'b10011101110011;
  assign mem[159] = 14'b01101101011011;
  assign mem[160] = 14'b01101100100001;
  assign mem[161] = 14'b00011110011101;
  assign mem[162] = 14'b10011000000011;
  assign mem[163] = 14'b10100100111111;
  assign mem[164] = 14'b01011110101001;
  assign mem[165] = 14'b00000101111010;
  assign mem[166] = 14'b01111010111111;
  assign mem[167] = 14'b10001000111011;
  assign mem[168] = 14'b10001011000101;
  assign mem[169] = 14'b10010000001101;
  assign mem[170] = 14'b10001010001110;
  assign mem[171] = 14'b01000111000111;
  assign mem[172] = 14'b10010101110101;
  assign mem[173] = 14'b10110110010000;
  assign mem[174] = 14'b01110111001110;
  assign mem[175] = 14'b10001001110101;
  assign mem[176] = 14'b01011000110000;
  assign mem[177] = 14'b01001101011100;
  assign mem[178] = 14'b01100001101011;
  assign mem[179] = 14'b10000011000100;
  assign mem[180] = 14'b10011110101100;
  assign mem[181] = 14'b10001000010011;
  assign mem[182] = 14'b00100100100101;
  assign mem[183] = 14'b00110001010111;
  assign mem[184] = 14'b00010110111011;
  assign mem[185] = 14'b01010101010100;
  assign mem[186] = 14'b10000101101001;
  assign mem[187] = 14'b01111001100111;
  assign mem[188] = 14'b00101001011001;
  assign mem[189] = 14'b00100100010000;
  assign mem[190] = 14'b10001101001100;
  assign mem[191] = 14'b01100000101100;
  assign mem[192] = 14'b00001011100001;
  assign mem[193] = 14'b00111001110010;
  assign mem[194] = 14'b01001001011011;
  assign mem[195] = 14'b01011001111001;
  assign mem[196] = 14'b10001101010110;
  assign mem[197] = 14'b00111001100111;
  assign mem[198] = 14'b00000000010000;
  assign mem[199] = 14'b00001110010010;
  assign mem[200] = 14'b01010001000010;
  assign mem[201] = 14'b10100100100011;
  assign mem[202] = 14'b01000111001000;
  assign mem[203] = 14'b00011110101100;
  assign mem[204] = 14'b00110110110101;
  assign mem[205] = 14'b10000011110100;
  assign mem[206] = 14'b01110101011100;
  assign mem[207] = 14'b01010100000101;
  assign mem[208] = 14'b10100111101101;
  assign mem[209] = 14'b00110011010001;
  assign mem[210] = 14'b01101101111101;
  assign mem[211] = 14'b00010000100100;
  assign mem[212] = 14'b00101101001111;
  assign mem[213] = 14'b01101111110100;
  assign mem[214] = 14'b10001010110111;
  assign mem[215] = 14'b01010011101101;
  assign mem[216] = 14'b01100100001001;
  assign mem[217] = 14'b10000000000101;
  assign mem[218] = 14'b00101110010010;
  assign mem[219] = 14'b01100011100111;
  assign mem[220] = 14'b01001111001000;
  assign mem[221] = 14'b01100111101010;
  assign mem[222] = 14'b01010111111001;
  assign mem[223] = 14'b00000100010110;
  assign mem[224] = 14'b00001110100100;
  assign mem[225] = 14'b10011111110101;
  assign mem[226] = 14'b10001011011111;
  assign mem[227] = 14'b01110111011010;
  assign mem[228] = 14'b00000101011111;
  assign mem[229] = 14'b10010001010010;
  assign mem[230] = 14'b00000011101101;
  assign mem[231] = 14'b01011011100010;
  assign mem[232] = 14'b01111000001100;
  assign mem[233] = 14'b00110001001010;
  assign mem[234] = 14'b10111101011110;
  assign mem[235] = 14'b01110110100010;
  assign mem[236] = 14'b00100000000101;
  assign mem[237] = 14'b10110000010101;
  assign mem[238] = 14'b00111011011010;
  assign mem[239] = 14'b01010001010100;
  assign mem[240] = 14'b01000111111010;
  assign mem[241] = 14'b00011011010100;
  assign mem[242] = 14'b10110000100100;
  assign mem[243] = 14'b00000101010100;
  assign mem[244] = 14'b00111001111111;
  assign mem[245] = 14'b01001000000110;
  assign mem[246] = 14'b00000100101100;
  assign mem[247] = 14'b10101011110001;
  assign mem[248] = 14'b01001111001110;
  assign mem[249] = 14'b10011101000001;
  assign mem[250] = 14'b10110101100000;
  assign mem[251] = 14'b10111111010111;
  assign mem[252] = 14'b01110011111101;
  assign mem[253] = 14'b10100111010011;
  assign mem[254] = 14'b01011001110010;
  assign mem[255] = 14'b01011000010110;
  assign mem[256] = 14'b00111011111011;
  assign mem[257] = 14'b01010110110001;
  assign mem[258] = 14'b00010011001000;
  assign mem[259] = 14'b10000100011100;
  assign mem[260] = 14'b10010000010101;
  assign mem[261] = 14'b00111100000101;
  assign mem[262] = 14'b00000011111010;
  assign mem[263] = 14'b10101111001001;
  assign mem[264] = 14'b01000010000001;
  assign mem[265] = 14'b01100010110110;
  assign mem[266] = 14'b10010111010000;
  assign mem[267] = 14'b10111111011110;
  assign mem[268] = 14'b01000000101000;
  assign mem[269] = 14'b00101011011010;
  assign mem[270] = 14'b00001010110100;
  assign mem[271] = 14'b10001001101000;
  assign mem[272] = 14'b01100100001010;
  assign mem[273] = 14'b01101000111110;
  assign mem[274] = 14'b10011101111001;
  assign mem[275] = 14'b10100010110010;
  assign mem[276] = 14'b00111010101111;
  assign mem[277] = 14'b01110010111100;
  assign mem[278] = 14'b10110001100001;
  assign mem[279] = 14'b10000011110001;
  assign mem[280] = 14'b01100100100101;
  assign mem[281] = 14'b00111001000100;
  assign mem[282] = 14'b01100011000110;
  assign mem[283] = 14'b10001100010010;
  assign mem[284] = 14'b01010100001111;
  assign mem[285] = 14'b00100011100000;
  assign mem[286] = 14'b01100101001100;
  assign mem[287] = 14'b01110011111000;
  assign mem[288] = 14'b10000011100010;
  assign mem[289] = 14'b10101001001000;
  assign mem[290] = 14'b10111011010010;
  assign mem[291] = 14'b01011001100101;
  assign mem[292] = 14'b00001101101100;
  assign mem[293] = 14'b01101101110110;
  assign mem[294] = 14'b00100001110111;
  assign mem[295] = 14'b00100110000100;
  assign mem[296] = 14'b00110101110010;
  assign mem[297] = 14'b10010000000001;
  assign mem[298] = 14'b10000000001110;
  assign mem[299] = 14'b01001011111010;
  assign mem[300] = 14'b01011101001100;
  assign mem[301] = 14'b00101010111010;
  assign mem[302] = 14'b01110000001010;
  assign mem[303] = 14'b00010110011010;
  assign mem[304] = 14'b01110011011101;
  assign mem[305] = 14'b10001010101111;
  assign mem[306] = 14'b10100110100101;
  assign mem[307] = 14'b10110011000001;
  assign mem[308] = 14'b01000001111100;
  assign mem[309] = 14'b00010110011000;
  assign mem[310] = 14'b10101001010000;
  assign mem[311] = 14'b01000011101000;
  assign mem[312] = 14'b10000101101101;
  assign mem[313] = 14'b00011101001011;
  assign mem[314] = 14'b10010011101110;
  assign mem[315] = 14'b00100101110000;
  assign mem[316] = 14'b00111011101000;
  assign mem[317] = 14'b10001101110100;
  assign mem[318] = 14'b00001010101110;
  assign mem[319] = 14'b01010100010001;
  assign mem[320] = 14'b00100111011011;
  assign mem[321] = 14'b01000011110011;
  assign mem[322] = 14'b01011111100011;
  assign mem[323] = 14'b00001001101011;
  assign mem[324] = 14'b00001110101001;
  assign mem[325] = 14'b00101100010010;
  assign mem[326] = 14'b01111001011111;
  assign mem[327] = 14'b00110011001111;
  assign mem[328] = 14'b00100100111011;
  assign mem[329] = 14'b01110101000000;
  assign mem[330] = 14'b01011111100000;
  assign mem[331] = 14'b01001111000000;
  assign mem[332] = 14'b00001100111000;
  assign mem[333] = 14'b10011111011100;
  assign mem[334] = 14'b10110110101010;
  assign mem[335] = 14'b00010001011001;
  assign mem[336] = 14'b00101010100111;
  assign mem[337] = 14'b10011001111000;
  assign mem[338] = 14'b00001110000000;
  assign mem[339] = 14'b00011111101100;
  assign mem[340] = 14'b01001111010011;
  assign mem[341] = 14'b00101001011110;
  assign mem[342] = 14'b10100011100000;
  assign mem[343] = 14'b01111011001100;
  assign mem[344] = 14'b10111110001001;
  assign mem[345] = 14'b01010100111010;
  assign mem[346] = 14'b00101111111110;
  assign mem[347] = 14'b01100100000000;
  assign mem[348] = 14'b10001110101100;
  assign mem[349] = 14'b10110110011000;
  assign mem[350] = 14'b10111101111001;
  assign mem[351] = 14'b01000110101000;
  assign mem[352] = 14'b00010011111001;
  assign mem[353] = 14'b10011000001011;
  assign mem[354] = 14'b10110011001100;
  assign mem[355] = 14'b10011011010001;
  assign mem[356] = 14'b10011100110111;
  assign mem[357] = 14'b10010111111000;
  assign mem[358] = 14'b00100011010110;
  assign mem[359] = 14'b10010010110111;
  assign mem[360] = 14'b10101110111000;
  assign mem[361] = 14'b00000100111011;
  assign mem[362] = 14'b01000110011111;
  assign mem[363] = 14'b00010010000110;
  assign mem[364] = 14'b01011110101101;
  assign mem[365] = 14'b01101001011111;
  assign mem[366] = 14'b10111001011001;
  assign mem[367] = 14'b00000101100101;
  assign mem[368] = 14'b01110011000111;
  assign mem[369] = 14'b01000111000110;
  assign mem[370] = 14'b00001111010111;
  assign mem[371] = 14'b10000101010110;
  assign mem[372] = 14'b10000010100000;
  assign mem[373] = 14'b10011110001110;
  assign mem[374] = 14'b01110101101010;
  assign mem[375] = 14'b10010000100101;
  assign mem[376] = 14'b01000100001111;
  assign mem[377] = 14'b01010001100101;
  assign mem[378] = 14'b00111110011111;
  assign mem[379] = 14'b10001001001001;
  assign mem[380] = 14'b00110001011001;
  assign mem[381] = 14'b01101101001110;
  assign mem[382] = 14'b01000000100010;
  assign mem[383] = 14'b10110110000100;
  assign mem[384] = 14'b00110100101110;
  assign mem[385] = 14'b10110011010101;
  assign mem[386] = 14'b00011011011001;
  assign mem[387] = 14'b00000100100100;
  assign mem[388] = 14'b10000111101001;
  assign mem[389] = 14'b00101011110110;
  assign mem[390] = 14'b10100010001010;
  assign mem[391] = 14'b10111110011100;
  assign mem[392] = 14'b01011010101000;
  assign mem[393] = 14'b10111000100011;
  assign mem[394] = 14'b00110001101101;
  assign mem[395] = 14'b00011111000100;
  assign mem[396] = 14'b00010000000000;
  assign mem[397] = 14'b10010001111100;
  assign mem[398] = 14'b00100110101101;
  assign mem[399] = 14'b10101010110000;
  assign mem[400] = 14'b01000111100110;
  assign mem[401] = 14'b01101001011110;
  assign mem[402] = 14'b00111000100011;
  assign mem[403] = 14'b01010101111111;
  assign mem[404] = 14'b01010001110001;
  assign mem[405] = 14'b00100110011111;
  assign mem[406] = 14'b10000100010110;
  assign mem[407] = 14'b01110111100010;
  assign mem[408] = 14'b01111100011100;
  assign mem[409] = 14'b01100011111011;
  assign mem[410] = 14'b00010000101111;
  assign mem[411] = 14'b00010011111000;
  assign mem[412] = 14'b00110110010010;
  assign mem[413] = 14'b10101100100101;
  assign mem[414] = 14'b00110011011011;
  assign mem[415] = 14'b10110001010000;
  assign mem[416] = 14'b10000100110110;
  assign mem[417] = 14'b10010100000110;
  assign mem[418] = 14'b10011001101101;
  assign mem[419] = 14'b00010011100101;
  assign mem[420] = 14'b00011101000001;
  assign mem[421] = 14'b01100001011001;
  assign mem[422] = 14'b01001001110000;
  assign mem[423] = 14'b10110100101001;
  assign mem[424] = 14'b01011110010010;
  assign mem[425] = 14'b10011001011001;
  assign mem[426] = 14'b00110100001011;
  assign mem[427] = 14'b00011100000101;
  assign mem[428] = 14'b00101100111111;
  assign mem[429] = 14'b01100001100010;
  assign mem[430] = 14'b01010001010000;
  assign mem[431] = 14'b00100001000010;
  assign mem[432] = 14'b01111100011010;
  assign mem[433] = 14'b10010010001001;
  assign mem[434] = 14'b10110001100011;
  assign mem[435] = 14'b01010101100011;
  assign mem[436] = 14'b01011111000100;
  assign mem[437] = 14'b10010110000001;
  assign mem[438] = 14'b01000000001100;
  assign mem[439] = 14'b01110010011011;
  assign mem[440] = 14'b10100011000110;
  assign mem[441] = 14'b10010011111111;
  assign mem[442] = 14'b00010011110111;
  assign mem[443] = 14'b00000110011000;
  assign mem[444] = 14'b01101011111111;
  assign mem[445] = 14'b00110000000111;
  assign mem[446] = 14'b00000101101000;
  assign mem[447] = 14'b10000001010100;
  assign mem[448] = 14'b10110100001111;
  assign mem[449] = 14'b10001111000100;
  assign mem[450] = 14'b10001101011001;
  assign mem[451] = 14'b10110100010011;
  assign mem[452] = 14'b00001101010010;
  assign mem[453] = 14'b10000110101001;
  assign mem[454] = 14'b00001100010000;
  assign mem[455] = 14'b01111011101111;
  assign mem[456] = 14'b10000010001110;
  assign mem[457] = 14'b10111110001010;
  assign mem[458] = 14'b00011100110110;
  assign mem[459] = 14'b10011111100101;
  assign mem[460] = 14'b10111110011000;
  assign mem[461] = 14'b01111010010011;
  assign mem[462] = 14'b10111001111111;
  assign mem[463] = 14'b01010111100000;
  assign mem[464] = 14'b10011000110011;
  assign mem[465] = 14'b00001111110100;
  assign mem[466] = 14'b00001011010001;
  assign mem[467] = 14'b00101011100000;
  assign mem[468] = 14'b01101000010100;
  assign mem[469] = 14'b01100110011000;
  assign mem[470] = 14'b01010011100100;
  assign mem[471] = 14'b01000101001000;
  assign mem[472] = 14'b01101010100000;
  assign mem[473] = 14'b10000011010101;
  assign mem[474] = 14'b10011011100111;
  assign mem[475] = 14'b01010000011110;
  assign mem[476] = 14'b00100100110100;
  assign mem[477] = 14'b01010110110000;
  assign mem[478] = 14'b01010010010011;
  assign mem[479] = 14'b00010100110101;
  assign mem[480] = 14'b10001001100001;
  assign mem[481] = 14'b10010110111101;
  assign mem[482] = 14'b01110010001100;
  assign mem[483] = 14'b01011010011100;
  assign mem[484] = 14'b01001100101110;
  assign mem[485] = 14'b00001110001101;
  assign mem[486] = 14'b10110101011101;
  assign mem[487] = 14'b01000100101011;
  assign mem[488] = 14'b10000000101110;
  assign mem[489] = 14'b01101000011110;
  assign mem[490] = 14'b01000011001110;
  assign mem[491] = 14'b00101111100100;
  assign mem[492] = 14'b00100011101101;
  assign mem[493] = 14'b10111111011001;
  assign mem[494] = 14'b00011110101011;
  assign mem[495] = 14'b10010000000000;
  assign mem[496] = 14'b01000011001000;
  assign mem[497] = 14'b10111010001110;
  assign mem[498] = 14'b00001010110111;
  assign mem[499] = 14'b01000100010011;
  assign mem[500] = 14'b10011001000001;
  assign mem[501] = 14'b01001100010100;
  assign mem[502] = 14'b00100101101011;
  assign mem[503] = 14'b10011111110110;
  assign mem[504] = 14'b00101001011010;
  assign mem[505] = 14'b00001101001001;
  assign mem[506] = 14'b00111100110010;
  assign mem[507] = 14'b10011111110111;
  assign mem[508] = 14'b01110001010000;
  assign mem[509] = 14'b10000100111001;
  assign mem[510] = 14'b10101110111100;
  assign mem[511] = 14'b01101000100000;
  assign mem[512] = 14'b00111111011011;
  assign mem[513] = 14'b01011110101100;
  assign mem[514] = 14'b00111001100110;
  assign mem[515] = 14'b01001001110010;
  assign mem[516] = 14'b10111001001101;
  assign mem[517] = 14'b01011010111000;
  assign mem[518] = 14'b01101110010010;
  assign mem[519] = 14'b01101011010100;
  assign mem[520] = 14'b10101110000001;
  assign mem[521] = 14'b01111011110110;
  assign mem[522] = 14'b01001100011110;
  assign mem[523] = 14'b10111111111100;
  assign mem[524] = 14'b01000000000110;
  assign mem[525] = 14'b00111101000100;
  assign mem[526] = 14'b00111000011010;
  assign mem[527] = 14'b01100101111101;
  assign mem[528] = 14'b01111100000010;
  assign mem[529] = 14'b01111100101110;
  assign mem[530] = 14'b10111011001001;
  assign mem[531] = 14'b01101001100011;
  assign mem[532] = 14'b00001000011001;
  assign mem[533] = 14'b01000111010010;
  assign mem[534] = 14'b00011001010111;
  assign mem[535] = 14'b10000000100011;
  assign mem[536] = 14'b10110010111101;
  assign mem[537] = 14'b01110101111000;
  assign mem[538] = 14'b00001110001010;
  assign mem[539] = 14'b10111000101000;
  assign mem[540] = 14'b10010101001100;
  assign mem[541] = 14'b10101001101010;
  assign mem[542] = 14'b10010111100111;
  assign mem[543] = 14'b00101011111111;
  assign mem[544] = 14'b10110111011000;
  assign mem[545] = 14'b01101010011101;
  assign mem[546] = 14'b01101101000011;
  assign mem[547] = 14'b00001100110011;
  assign mem[548] = 14'b10001011000111;
  assign mem[549] = 14'b01100001111111;
  assign mem[550] = 14'b10101001011011;
  assign mem[551] = 14'b00000101011100;
  assign mem[552] = 14'b01110101011010;
  assign mem[553] = 14'b10000010010011;
  assign mem[554] = 14'b01100100100111;
  assign mem[555] = 14'b00001010110110;
  assign mem[556] = 14'b00001101010100;
  assign mem[557] = 14'b01011000011011;
  assign mem[558] = 14'b00101011011101;
  assign mem[559] = 14'b00111010000100;
  assign mem[560] = 14'b10110101000101;
  assign mem[561] = 14'b00101111010000;
  assign mem[562] = 14'b00010111110011;
  assign mem[563] = 14'b10000111010011;
  assign mem[564] = 14'b01000000010010;
  assign mem[565] = 14'b10100111110010;
  assign mem[566] = 14'b00110011100111;
  assign mem[567] = 14'b01011011111101;
  assign mem[568] = 14'b00101110100010;
  assign mem[569] = 14'b01110001111001;
  assign mem[570] = 14'b10111001101100;
  assign mem[571] = 14'b10001110100011;
  assign mem[572] = 14'b10010001101011;
  assign mem[573] = 14'b10111000110110;
  assign mem[574] = 14'b00000001100010;
  assign mem[575] = 14'b00100111011110;
  assign mem[576] = 14'b00100001000100;
  assign mem[577] = 14'b01000000100011;
  assign mem[578] = 14'b10110010001111;
  assign mem[579] = 14'b00011100110100;
  assign mem[580] = 14'b00111000111101;
  assign mem[581] = 14'b00111101001100;
  assign mem[582] = 14'b01111111000101;
  assign mem[583] = 14'b00100010110000;
  assign mem[584] = 14'b10101001110111;
  assign mem[585] = 14'b01111110011100;
  assign mem[586] = 14'b10010110110011;
  assign mem[587] = 14'b01011101100101;
  assign mem[588] = 14'b01101111100100;
  assign mem[589] = 14'b10000100100000;
  assign mem[590] = 14'b00011010000110;
  assign mem[591] = 14'b00000010011111;
  assign mem[592] = 14'b10101010101011;
  assign mem[593] = 14'b01001100110110;
  assign mem[594] = 14'b00000010000000;
  assign mem[595] = 14'b01110010010000;
  assign mem[596] = 14'b00001011010101;
  assign mem[597] = 14'b10001111000101;
  assign mem[598] = 14'b01001110001110;
  assign mem[599] = 14'b01100011111001;
  assign mem[600] = 14'b00110110100110;
  assign mem[601] = 14'b01011110011011;
  assign mem[602] = 14'b10101011011100;
  assign mem[603] = 14'b01100000100101;
  assign mem[604] = 14'b10111000111110;
  assign mem[605] = 14'b00110101011111;
  assign mem[606] = 14'b10100100010010;
  assign mem[607] = 14'b01110111110100;
  assign mem[608] = 14'b00111001101101;
  assign mem[609] = 14'b01101000000010;
  assign mem[610] = 14'b01101011111001;
  assign mem[611] = 14'b10111010110001;
  assign mem[612] = 14'b10011111100100;
  assign mem[613] = 14'b10111010010010;
  assign mem[614] = 14'b10001110001101;
  assign mem[615] = 14'b10000010101101;
  assign mem[616] = 14'b01001111110110;
  assign mem[617] = 14'b00000000101101;
  assign mem[618] = 14'b00100101100000;
  assign mem[619] = 14'b00011110000001;
  assign mem[620] = 14'b01000100011001;
  assign mem[621] = 14'b00101010100000;
  assign mem[622] = 14'b00011010011111;
  assign mem[623] = 14'b00000000110011;
  assign mem[624] = 14'b00101011111000;
  assign mem[625] = 14'b00001010001010;
  assign mem[626] = 14'b00011101101000;
  assign mem[627] = 14'b10011100001101;
  assign mem[628] = 14'b10011011110011;
  assign mem[629] = 14'b10111011001100;
  assign mem[630] = 14'b01111110100010;
  assign mem[631] = 14'b01001011100001;
  assign mem[632] = 14'b01000000100111;
  assign mem[633] = 14'b01000010100001;
  assign mem[634] = 14'b01011011001110;
  assign mem[635] = 14'b01001010011101;
  assign mem[636] = 14'b10101011101001;
  assign mem[637] = 14'b10110100001100;
  assign mem[638] = 14'b00001001001110;
  assign mem[639] = 14'b10111110100110;
  assign mem[640] = 14'b00000111100010;
  assign mem[641] = 14'b10111110001101;
  assign mem[642] = 14'b00011111010110;
  assign mem[643] = 14'b01101110011000;
  assign mem[644] = 14'b10011100100010;
  assign mem[645] = 14'b00111101001000;
  assign mem[646] = 14'b10111011110000;
  assign mem[647] = 14'b10100100010111;
  assign mem[648] = 14'b10110001100010;
  assign mem[649] = 14'b01101100101010;
  assign mem[650] = 14'b00100010100010;
  assign mem[651] = 14'b00000100011100;
  assign mem[652] = 14'b01010100100101;
  assign mem[653] = 14'b01100111001001;
  assign mem[654] = 14'b00111100011001;
  assign mem[655] = 14'b10100001100011;
  assign mem[656] = 14'b10101110110100;
  assign mem[657] = 14'b01100001010111;
  assign mem[658] = 14'b00001000000101;
  assign mem[659] = 14'b10010101011100;
  assign mem[660] = 14'b10110000010001;
  assign mem[661] = 14'b00111100010111;
  assign mem[662] = 14'b00010010111010;
  assign mem[663] = 14'b01000111111100;
  assign mem[664] = 14'b01111111100000;
  assign mem[665] = 14'b10110010110111;
  assign mem[666] = 14'b00000010011001;
  assign mem[667] = 14'b01110000100100;
  assign mem[668] = 14'b01011010000011;
  assign mem[669] = 14'b01001111100001;
  assign mem[670] = 14'b10010000100000;
  assign mem[671] = 14'b10111101111010;
  assign mem[672] = 14'b10110111100100;
  assign mem[673] = 14'b00010101001010;
  assign mem[674] = 14'b01101000010000;
  assign mem[675] = 14'b00000010110011;
  assign mem[676] = 14'b01010110011100;
  assign mem[677] = 14'b00101001010110;
  assign mem[678] = 14'b01011100110101;
  assign mem[679] = 14'b10111110011001;
  assign mem[680] = 14'b00001101011110;
  assign mem[681] = 14'b00110001010110;
  assign mem[682] = 14'b00000111011101;
  assign mem[683] = 14'b01110001101111;
  assign mem[684] = 14'b01011000101110;
  assign mem[685] = 14'b01111011101010;
  assign mem[686] = 14'b01000010011110;
  assign mem[687] = 14'b00000100101110;
  assign mem[688] = 14'b00101101001101;
  assign mem[689] = 14'b10011110000010;
  assign mem[690] = 14'b01101011101010;
  assign mem[691] = 14'b10010101011000;
  assign mem[692] = 14'b10010110101111;
  assign mem[693] = 14'b10111010000001;
  assign mem[694] = 14'b01000000000010;
  assign mem[695] = 14'b10011001100000;
  assign mem[696] = 14'b10100000011101;
  assign mem[697] = 14'b00010101001001;
  assign mem[698] = 14'b10100111011011;
  assign mem[699] = 14'b01010011001101;
  assign mem[700] = 14'b01100001101110;
  assign mem[701] = 14'b00111101101111;
  assign mem[702] = 14'b00011100001111;
  assign mem[703] = 14'b01100100110001;
  assign mem[704] = 14'b01010000100111;
  assign mem[705] = 14'b00010100011100;
  assign mem[706] = 14'b10000001111011;
  assign mem[707] = 14'b00110101001100;
  assign mem[708] = 14'b00011101010101;
  assign mem[709] = 14'b00010011001111;
  assign mem[710] = 14'b00000001110000;
  assign mem[711] = 14'b01100011111110;
  assign mem[712] = 14'b10110111001100;
  assign mem[713] = 14'b10111111110000;
  assign mem[714] = 14'b01110001110110;
  assign mem[715] = 14'b00010110110011;
  assign mem[716] = 14'b10111111110010;
  assign mem[717] = 14'b10011010101000;
  assign mem[718] = 14'b00110110000000;
  assign mem[719] = 14'b00001100100000;
  assign mem[720] = 14'b00010101110101;
  assign mem[721] = 14'b10100110110110;
  assign mem[722] = 14'b00000001100111;
  assign mem[723] = 14'b01110011111100;
  assign mem[724] = 14'b01111100101000;
  assign mem[725] = 14'b00001110101000;
  assign mem[726] = 14'b00001011111100;
  assign mem[727] = 14'b00001001111000;
  assign mem[728] = 14'b01111100111100;
  assign mem[729] = 14'b10000000011111;
  assign mem[730] = 14'b10000011111101;
  assign mem[731] = 14'b01111001001110;
  assign mem[732] = 14'b10101001110110;
  assign mem[733] = 14'b10010101100011;
  assign mem[734] = 14'b00100111001100;
  assign mem[735] = 14'b00011110011010;
  assign mem[736] = 14'b01100101111100;
  assign mem[737] = 14'b10011110101110;
  assign mem[738] = 14'b00010000010100;
  assign mem[739] = 14'b01000011110010;
  assign mem[740] = 14'b00100110011001;
  assign mem[741] = 14'b00111000111001;
  assign mem[742] = 14'b00011001111011;
  assign mem[743] = 14'b01000000101011;
  assign mem[744] = 14'b01001001010000;
  assign mem[745] = 14'b10011000000101;
  assign mem[746] = 14'b10101110001100;
  assign mem[747] = 14'b00111101101010;
  assign mem[748] = 14'b00100000100010;
  assign mem[749] = 14'b01010010001101;
  assign mem[750] = 14'b00011111110100;
  assign mem[751] = 14'b10111001001010;
  assign mem[752] = 14'b01110111010100;
  assign mem[753] = 14'b10111111001100;
  assign mem[754] = 14'b01010011110110;
  assign mem[755] = 14'b00100101001100;
  assign mem[756] = 14'b00010101110111;
  assign mem[757] = 14'b01111000101000;
  assign mem[758] = 14'b00100000110100;
  assign mem[759] = 14'b00110010010001;
  assign mem[760] = 14'b10101010100000;
  assign mem[761] = 14'b10001011000010;
  assign mem[762] = 14'b01110110011010;
  assign mem[763] = 14'b10111011011011;
  assign mem[764] = 14'b00101011100111;
  assign mem[765] = 14'b00010010111111;
  assign mem[766] = 14'b00110100011011;
  assign mem[767] = 14'b00101010010111;
  assign mem[768] = 14'b00100011011011;
  assign mem[769] = 14'b00011111010100;
  assign mem[770] = 14'b10000101111000;
  assign mem[771] = 14'b10011111000000;
  assign mem[772] = 14'b00110010001110;
  assign mem[773] = 14'b00100100100001;
  assign mem[774] = 14'b00011011010110;
  assign mem[775] = 14'b01001001111001;
  assign mem[776] = 14'b01001110000101;
  assign mem[777] = 14'b01110011110111;
  assign mem[778] = 14'b01100010101011;
  assign mem[779] = 14'b10111100001100;
  assign mem[780] = 14'b01000100010110;
  assign mem[781] = 14'b01101111110101;
  assign mem[782] = 14'b01001011101100;
  assign mem[783] = 14'b00000011010011;
  assign mem[784] = 14'b01111101000011;
  assign mem[785] = 14'b10011110101111;
  assign mem[786] = 14'b10010001001010;
  assign mem[787] = 14'b10110011011001;
  assign mem[788] = 14'b00011011000111;
  assign mem[789] = 14'b00100100100000;
  assign mem[790] = 14'b01011010100001;
  assign mem[791] = 14'b10011010010011;
  assign mem[792] = 14'b10000000000000;
  assign mem[793] = 14'b00001111011010;
  assign mem[794] = 14'b01110101100111;
  assign mem[795] = 14'b00010101111001;
  assign mem[796] = 14'b00001101100110;
  assign mem[797] = 14'b00111000011111;
  assign mem[798] = 14'b10000100010001;
  assign mem[799] = 14'b00101011000100;
  assign mem[800] = 14'b10011000101010;
  assign mem[801] = 14'b00011111110010;
  assign mem[802] = 14'b10011110111000;
  assign mem[803] = 14'b00110011000000;
  assign mem[804] = 14'b01011111110100;
  assign mem[805] = 14'b00000000110110;
  assign mem[806] = 14'b00101101000000;
  assign mem[807] = 14'b01001010011011;
  assign mem[808] = 14'b10111000011101;
  assign mem[809] = 14'b00110000000010;
  assign mem[810] = 14'b10000001011110;
  assign mem[811] = 14'b10010011010100;
  assign mem[812] = 14'b01001100010001;
  assign mem[813] = 14'b01101100010101;
  assign mem[814] = 14'b00010001000010;
  assign mem[815] = 14'b10011100110110;
  assign mem[816] = 14'b00101000000111;
  assign mem[817] = 14'b00001011000100;
  assign mem[818] = 14'b00001101111101;
  assign mem[819] = 14'b01100101000001;
  assign mem[820] = 14'b01001101100010;
  assign mem[821] = 14'b10011100101000;
  assign mem[822] = 14'b00100000101010;
  assign mem[823] = 14'b01011001010110;
  assign mem[824] = 14'b10100111110111;
  assign mem[825] = 14'b00001100001100;
  assign mem[826] = 14'b01001001111101;
  assign mem[827] = 14'b01001000001111;
  assign mem[828] = 14'b00100001010110;
  assign mem[829] = 14'b00100000100111;
  assign mem[830] = 14'b01001011000010;
  assign mem[831] = 14'b00001101110100;
  assign mem[832] = 14'b01010011111100;
  assign mem[833] = 14'b01011010100011;
  assign mem[834] = 14'b01011100110010;
  assign mem[835] = 14'b01000011101101;
  assign mem[836] = 14'b01100110011111;
  assign mem[837] = 14'b01110101111101;
  assign mem[838] = 14'b01010010010101;
  assign mem[839] = 14'b10100110101000;
  assign mem[840] = 14'b01000010011100;
  assign mem[841] = 14'b00110010111100;
  assign mem[842] = 14'b01011100011101;
  assign mem[843] = 14'b10101000111110;
  assign mem[844] = 14'b01011010001000;
  assign mem[845] = 14'b10011011111111;
  assign mem[846] = 14'b01111110100000;
  assign mem[847] = 14'b01111001101111;
  assign mem[848] = 14'b01101010010000;
  assign mem[849] = 14'b01110101000011;
  assign mem[850] = 14'b01100010000000;
  assign mem[851] = 14'b00011101110011;
  assign mem[852] = 14'b10101011000011;
  assign mem[853] = 14'b01100010010001;
  assign mem[854] = 14'b10111000011011;
  assign mem[855] = 14'b01011110010000;
  assign mem[856] = 14'b10110010111001;
  assign mem[857] = 14'b00010010010011;
  assign mem[858] = 14'b10001111110001;
  assign mem[859] = 14'b01111011111101;
  assign mem[860] = 14'b00100110101111;
  assign mem[861] = 14'b01111100100010;
  assign mem[862] = 14'b10110001001001;
  assign mem[863] = 14'b01101110010110;
  assign mem[864] = 14'b10001011001111;
  assign mem[865] = 14'b01101001001000;
  assign mem[866] = 14'b01100110001110;
  assign mem[867] = 14'b01111110110010;
  assign mem[868] = 14'b10001001111100;
  assign mem[869] = 14'b01100111000011;
  assign mem[870] = 14'b00110111011001;
  assign mem[871] = 14'b01000011111100;
  assign mem[872] = 14'b01001000000010;
  assign mem[873] = 14'b00100010011101;
  assign mem[874] = 14'b01101101010111;
  assign mem[875] = 14'b01111110101010;
  assign mem[876] = 14'b01010110111000;
  assign mem[877] = 14'b10100010010110;
  assign mem[878] = 14'b10010001101001;
  assign mem[879] = 14'b00100111000011;
  assign mem[880] = 14'b00100101101101;
  assign mem[881] = 14'b01110001101000;
  assign mem[882] = 14'b01101011100001;
  assign mem[883] = 14'b10100101010110;
  assign mem[884] = 14'b10010001011100;
  assign mem[885] = 14'b10010011011101;
  assign mem[886] = 14'b00110111100010;
  assign mem[887] = 14'b00110011111110;
  assign mem[888] = 14'b01011101100111;
  assign mem[889] = 14'b10111011000001;
  assign mem[890] = 14'b00110101010111;
  assign mem[891] = 14'b10111111111011;
  assign mem[892] = 14'b10011001101110;
  assign mem[893] = 14'b10111100011111;
  assign mem[894] = 14'b01000011101100;
  assign mem[895] = 14'b01111010010110;
  assign mem[896] = 14'b10110001000001;
  assign mem[897] = 14'b01100111001101;
  assign mem[898] = 14'b10111111101111;
  assign mem[899] = 14'b00011111111100;
  assign mem[900] = 14'b10110101011011;
  assign mem[901] = 14'b01110010111001;
  assign mem[902] = 14'b10101111000001;
  assign mem[903] = 14'b10110100111110;
  assign mem[904] = 14'b00111010010101;
  assign mem[905] = 14'b10001011101111;
  assign mem[906] = 14'b10011011111010;
  assign mem[907] = 14'b00011001011011;
  assign mem[908] = 14'b01110000000000;
  assign mem[909] = 14'b00111101011111;
  assign mem[910] = 14'b01001110111010;
  assign mem[911] = 14'b00101011001010;
  assign mem[912] = 14'b01110101001000;
  assign mem[913] = 14'b10100010001111;
  assign mem[914] = 14'b00001011110011;
  assign mem[915] = 14'b00011001110110;
  assign mem[916] = 14'b10111100010101;
  assign mem[917] = 14'b01001101011000;
  assign mem[918] = 14'b10011110010110;
  assign mem[919] = 14'b01000100101010;
  assign mem[920] = 14'b01100111000000;
  assign mem[921] = 14'b01111011011010;
  assign mem[922] = 14'b01110101001001;
  assign mem[923] = 14'b10001011001000;
  assign mem[924] = 14'b10111011111101;
  assign mem[925] = 14'b00110111111101;
  assign mem[926] = 14'b10100111111100;
  assign mem[927] = 14'b01011000101010;
  assign mem[928] = 14'b10100001110110;
  assign mem[929] = 14'b01001100100101;
  assign mem[930] = 14'b01110011110110;
  assign mem[931] = 14'b10001001000011;
  assign mem[932] = 14'b00001011000110;
  assign mem[933] = 14'b01101001101100;
  assign mem[934] = 14'b10000100001110;
  assign mem[935] = 14'b01110000011001;
  assign mem[936] = 14'b01010011111011;
  assign mem[937] = 14'b01110001101010;
  assign mem[938] = 14'b10101101001100;
  assign mem[939] = 14'b00000100100010;
  assign mem[940] = 14'b01111010111000;
  assign mem[941] = 14'b01101010101011;
  assign mem[942] = 14'b10111000101110;
  assign mem[943] = 14'b00100111001101;
  assign mem[944] = 14'b01100110110010;
  assign mem[945] = 14'b00111110111010;
  assign mem[946] = 14'b01011010101111;
  assign mem[947] = 14'b00010110110010;
  assign mem[948] = 14'b01011001011001;
  assign mem[949] = 14'b01011010000010;
  assign mem[950] = 14'b01000001010010;
  assign mem[951] = 14'b00100000111001;
  assign mem[952] = 14'b10110101100101;
  assign mem[953] = 14'b01001011110100;
  assign mem[954] = 14'b10001011000001;
  assign mem[955] = 14'b00101100101000;
  assign mem[956] = 14'b10110011110110;
  assign mem[957] = 14'b10010000110000;
  assign mem[958] = 14'b00100111011000;
  assign mem[959] = 14'b10001001001000;
  assign mem[960] = 14'b01101101100011;
  assign mem[961] = 14'b00101001010111;
  assign mem[962] = 14'b00011101101010;
  assign mem[963] = 14'b01101101111111;
  assign mem[964] = 14'b01011100111110;
  assign mem[965] = 14'b10101110011011;
  assign mem[966] = 14'b01010101110000;
  assign mem[967] = 14'b01100010000101;
  assign mem[968] = 14'b10001111011110;
  assign mem[969] = 14'b10110011000000;
  assign mem[970] = 14'b00001001111001;
  assign mem[971] = 14'b10011100111110;
  assign mem[972] = 14'b10110100100010;
  assign mem[973] = 14'b01011000000001;
  assign mem[974] = 14'b10010101110011;
  assign mem[975] = 14'b00100100011101;
  assign mem[976] = 14'b01101101100000;
  assign mem[977] = 14'b01101110101100;
  assign mem[978] = 14'b01001110110111;
  assign mem[979] = 14'b01110000011111;
  assign mem[980] = 14'b10011010001001;
  assign mem[981] = 14'b10001100100101;
  assign mem[982] = 14'b00001000111001;
  assign mem[983] = 14'b01100011110110;
  assign mem[984] = 14'b10101001011101;
  assign mem[985] = 14'b10010111001111;
  assign mem[986] = 14'b10000001001100;
  assign mem[987] = 14'b10110011010000;
  assign mem[988] = 14'b01000001101011;
  assign mem[989] = 14'b00011111001101;
  assign mem[990] = 14'b00000000000010;
  assign mem[991] = 14'b10010001110011;
  assign mem[992] = 14'b00000010100010;
  assign mem[993] = 14'b01100000100110;
  assign mem[994] = 14'b00011111010000;
  assign mem[995] = 14'b00111001000001;
  assign mem[996] = 14'b10011001000000;
  assign mem[997] = 14'b01100011011011;
  assign mem[998] = 14'b01110110000101;
  assign mem[999] = 14'b01100000101011;
  assign mem[1000] = 14'b10000100111110;
  assign mem[1001] = 14'b10011011001111;
  assign mem[1002] = 14'b01010110100000;
  assign mem[1003] = 14'b10001100111011;
  assign mem[1004] = 14'b00111001111010;
  assign mem[1005] = 14'b10111011101001;
  assign mem[1006] = 14'b00010110101100;
  assign mem[1007] = 14'b00101111111011;
  assign mem[1008] = 14'b01010101110110;
  assign mem[1009] = 14'b10010111011100;
  assign mem[1010] = 14'b01001100000001;
  assign mem[1011] = 14'b01011110000011;
  assign mem[1012] = 14'b01101111000010;
  assign mem[1013] = 14'b10010110001010;
  assign mem[1014] = 14'b01000111101100;
  assign mem[1015] = 14'b10011110110101;
  assign mem[1016] = 14'b01100001110101;
  assign mem[1017] = 14'b01011011111111;
  assign mem[1018] = 14'b00101001011100;
  assign mem[1019] = 14'b10011110111100;
  assign mem[1020] = 14'b00011000101100;
  assign mem[1021] = 14'b10100010001011;
  assign mem[1022] = 14'b01001000011110;
  assign mem[1023] = 14'b10011011011101;
  always@(*)
  begin
    data_out_t <= mem[addr_f];
  end
  wire [13:0] data_out_reg [n_outreg:0];
  generate if (n_outreg > 0)
  begin
    for( i=n_outreg-1; i >= 1; i=i-1)
    begin: data_out_reg_stage
      mgc_generic_reg #(
        .width(14),
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_data_out_reg (
        .d(data_out_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(data_out_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(14),
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_data_out_reg_init (
      .d(data_out_t),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(data_out_reg[0])
    );
    assign data_out = data_out_reg[n_outreg-1];
  end
  else
  begin
    assign data_out = data_out_t;
  end
  endgenerate
endmodule
module stagemgc_rom_sync_regout_11_1024_14_1_0_0_1_0_1_0_0_0_1_60 (addr, data_out,
    clk, s_rst, a_rst, en
);
  input [9:0]addr ;
  output [13:0]data_out ;
  input clk ;
  input s_rst ;
  input a_rst ;
  input en ;
  parameter n_width = 14;
  parameter n_size = 1024;
  parameter n_numports = 1;
  parameter n_addr_w = 10;
  parameter n_inreg = 0;
  parameter n_outreg = 1;
  wire [9:0] addr_f;
  wire [9:0] addr_reg [n_inreg:0];
  genvar i;
  generate if (n_inreg > 0)
  begin
    for( i=n_inreg-1; i >= 1; i=i-1)
    begin: addr_reg_stage
      mgc_generic_reg #(
        .width(10),
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_addr_reg (
        .d(addr_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(addr_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(10),
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_addr_reg_init (
      .d(addr),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(addr_reg[0])
    );
    assign addr_f = addr_reg[n_inreg-1];
  end
  else
  begin
    assign addr_f = addr;
  end
  endgenerate
  wire [13:0] mem [1023:0];
  reg [13:0] data_out_t;
  assign mem[0] = 14'b00111111111011;
  assign mem[1] = 14'b01000100110001;
  assign mem[2] = 14'b00010000111001;
  assign mem[3] = 14'b00010011001101;
  assign mem[4] = 14'b00100111100010;
  assign mem[5] = 14'b01011101111110;
  assign mem[6] = 14'b01111100001011;
  assign mem[7] = 14'b01010011010001;
  assign mem[8] = 14'b00101000010011;
  assign mem[9] = 14'b01001010001111;
  assign mem[10] = 14'b01100101000000;
  assign mem[11] = 14'b10110110110111;
  assign mem[12] = 14'b01101101101111;
  assign mem[13] = 14'b00101011111100;
  assign mem[14] = 14'b01011100000010;
  assign mem[15] = 14'b10100111001010;
  assign mem[16] = 14'b00110000100101;
  assign mem[17] = 14'b00100001001101;
  assign mem[18] = 14'b00011110101000;
  assign mem[19] = 14'b10101010101101;
  assign mem[20] = 14'b10100101101001;
  assign mem[21] = 14'b10100010100100;
  assign mem[22] = 14'b01000001011101;
  assign mem[23] = 14'b00011101010011;
  assign mem[24] = 14'b01011011010111;
  assign mem[25] = 14'b10000101100010;
  assign mem[26] = 14'b01001000000111;
  assign mem[27] = 14'b01010001000110;
  assign mem[28] = 14'b10110000111100;
  assign mem[29] = 14'b10100101010010;
  assign mem[30] = 14'b01011011111010;
  assign mem[31] = 14'b10101110010011;
  assign mem[32] = 14'b10000011100001;
  assign mem[33] = 14'b10111111110011;
  assign mem[34] = 14'b10100101100111;
  assign mem[35] = 14'b01110100010110;
  assign mem[36] = 14'b01011001010111;
  assign mem[37] = 14'b00110111110001;
  assign mem[38] = 14'b01011101011101;
  assign mem[39] = 14'b10011101111100;
  assign mem[40] = 14'b01000101001010;
  assign mem[41] = 14'b10000001110010;
  assign mem[42] = 14'b10101000000011;
  assign mem[43] = 14'b01001001000111;
  assign mem[44] = 14'b10101100101100;
  assign mem[45] = 14'b00011000000010;
  assign mem[46] = 14'b10111001010001;
  assign mem[47] = 14'b00000001100100;
  assign mem[48] = 14'b10000000110111;
  assign mem[49] = 14'b01100111100001;
  assign mem[50] = 14'b10010111111101;
  assign mem[51] = 14'b01010000011001;
  assign mem[52] = 14'b00110101010100;
  assign mem[53] = 14'b01111010110010;
  assign mem[54] = 14'b01011011000111;
  assign mem[55] = 14'b10010011110100;
  assign mem[56] = 14'b01010001100001;
  assign mem[57] = 14'b10100111110100;
  assign mem[58] = 14'b01111011001010;
  assign mem[59] = 14'b01110101010010;
  assign mem[60] = 14'b10111110001100;
  assign mem[61] = 14'b10110000011100;
  assign mem[62] = 14'b01011110100001;
  assign mem[63] = 14'b00000001001111;
  assign mem[64] = 14'b00000000001101;
  assign mem[65] = 14'b01101100011010;
  assign mem[66] = 14'b10001010110110;
  assign mem[67] = 14'b01010101001101;
  assign mem[68] = 14'b01000111101010;
  assign mem[69] = 14'b10110010111111;
  assign mem[70] = 14'b00101101010111;
  assign mem[71] = 14'b01001001000100;
  assign mem[72] = 14'b10011001110011;
  assign mem[73] = 14'b01110111000101;
  assign mem[74] = 14'b10001001110110;
  assign mem[75] = 14'b10001110010101;
  assign mem[76] = 14'b00100000100011;
  assign mem[77] = 14'b10000100111011;
  assign mem[78] = 14'b10000111101101;
  assign mem[79] = 14'b00110000100110;
  assign mem[80] = 14'b01101101100111;
  assign mem[81] = 14'b00110011000101;
  assign mem[82] = 14'b00010101010111;
  assign mem[83] = 14'b01100011111101;
  assign mem[84] = 14'b10100000010011;
  assign mem[85] = 14'b10000011110011;
  assign mem[86] = 14'b10100100011111;
  assign mem[87] = 14'b10110100100111;
  assign mem[88] = 14'b10101101010110;
  assign mem[89] = 14'b00100010100011;
  assign mem[90] = 14'b00011100010000;
  assign mem[91] = 14'b01110010010111;
  assign mem[92] = 14'b00000000110000;
  assign mem[93] = 14'b10010101001011;
  assign mem[94] = 14'b00101000000000;
  assign mem[95] = 14'b00010011001100;
  assign mem[96] = 14'b10010011011110;
  assign mem[97] = 14'b10101000100011;
  assign mem[98] = 14'b10111000011000;
  assign mem[99] = 14'b00011100011100;
  assign mem[100] = 14'b10110010001110;
  assign mem[101] = 14'b10001100000110;
  assign mem[102] = 14'b01100000001111;
  assign mem[103] = 14'b00101111000100;
  assign mem[104] = 14'b01011111011101;
  assign mem[105] = 14'b00101011101100;
  assign mem[106] = 14'b00100010011011;
  assign mem[107] = 14'b00011001110100;
  assign mem[108] = 14'b00001011000111;
  assign mem[109] = 14'b01101101011100;
  assign mem[110] = 14'b00010000011101;
  assign mem[111] = 14'b10001100001101;
  assign mem[112] = 14'b01010001111100;
  assign mem[113] = 14'b00010111101101;
  assign mem[114] = 14'b10010001101010;
  assign mem[115] = 14'b10110000000101;
  assign mem[116] = 14'b00001110000100;
  assign mem[117] = 14'b00111100110000;
  assign mem[118] = 14'b10101101111101;
  assign mem[119] = 14'b10100111110000;
  assign mem[120] = 14'b01001101010101;
  assign mem[121] = 14'b01110111000000;
  assign mem[122] = 14'b10011011110110;
  assign mem[123] = 14'b01001010001010;
  assign mem[124] = 14'b10100000011110;
  assign mem[125] = 14'b00000001111110;
  assign mem[126] = 14'b00101101101001;
  assign mem[127] = 14'b01101001000000;
  assign mem[128] = 14'b01100111101011;
  assign mem[129] = 14'b01100110001111;
  assign mem[130] = 14'b00011000101110;
  assign mem[131] = 14'b01001100000100;
  assign mem[132] = 14'b00000000101010;
  assign mem[133] = 14'b00001010100001;
  assign mem[134] = 14'b00100011000000;
  assign mem[135] = 14'b01110000110011;
  assign mem[136] = 14'b00010100010000;
  assign mem[137] = 14'b10111011010101;
  assign mem[138] = 14'b01110111111011;
  assign mem[139] = 14'b10000110000010;
  assign mem[140] = 14'b10111010101101;
  assign mem[141] = 14'b00001111011101;
  assign mem[142] = 14'b10100100101101;
  assign mem[143] = 14'b01111000000111;
  assign mem[144] = 14'b01101110101101;
  assign mem[145] = 14'b10000100100111;
  assign mem[146] = 14'b00001111101100;
  assign mem[147] = 14'b10011111111100;
  assign mem[148] = 14'b01001001011111;
  assign mem[149] = 14'b00000010100011;
  assign mem[150] = 14'b10001110110111;
  assign mem[151] = 14'b01000111110101;
  assign mem[152] = 14'b01100100011111;
  assign mem[153] = 14'b10111100010100;
  assign mem[154] = 14'b00101110101111;
  assign mem[155] = 14'b10111010100010;
  assign mem[156] = 14'b01001000100111;
  assign mem[157] = 14'b00110100100010;
  assign mem[158] = 14'b00100000001100;
  assign mem[159] = 14'b10110001011101;
  assign mem[160] = 14'b10111011101011;
  assign mem[161] = 14'b01101000001000;
  assign mem[162] = 14'b01011000010111;
  assign mem[163] = 14'b01110000111001;
  assign mem[164] = 14'b01011100011010;
  assign mem[165] = 14'b10010001101111;
  assign mem[166] = 14'b00111111111100;
  assign mem[167] = 14'b01011011111000;
  assign mem[168] = 14'b01101100010100;
  assign mem[169] = 14'b00110101001010;
  assign mem[170] = 14'b01010000001101;
  assign mem[171] = 14'b10010010110010;
  assign mem[172] = 14'b10101111011101;
  assign mem[173] = 14'b01010010000100;
  assign mem[174] = 14'b10001100110000;
  assign mem[175] = 14'b00011000010100;
  assign mem[176] = 14'b01101011111100;
  assign mem[177] = 14'b01001010100101;
  assign mem[178] = 14'b00111100001101;
  assign mem[179] = 14'b10001001001100;
  assign mem[180] = 14'b10100001010101;
  assign mem[181] = 14'b01111000111001;
  assign mem[182] = 14'b00011011011110;
  assign mem[183] = 14'b01101110111111;
  assign mem[184] = 14'b10110001101111;
  assign mem[185] = 14'b10111111110001;
  assign mem[186] = 14'b10000110011010;
  assign mem[187] = 14'b00110010101011;
  assign mem[188] = 14'b01100110001000;
  assign mem[189] = 14'b01110110100110;
  assign mem[190] = 14'b10000110001111;
  assign mem[191] = 14'b10110100100000;
  assign mem[192] = 14'b01011111010101;
  assign mem[193] = 14'b00110010110101;
  assign mem[194] = 14'b10011011110001;
  assign mem[195] = 14'b10010110101000;
  assign mem[196] = 14'b01000110011010;
  assign mem[197] = 14'b00111010011000;
  assign mem[198] = 14'b01101010101101;
  assign mem[199] = 14'b10101001000110;
  assign mem[200] = 14'b10001110101010;
  assign mem[201] = 14'b10011011011100;
  assign mem[202] = 14'b00110111101110;
  assign mem[203] = 14'b00100001010101;
  assign mem[204] = 14'b00111100111101;
  assign mem[205] = 14'b01011110010110;
  assign mem[206] = 14'b01110010100101;
  assign mem[207] = 14'b01100111010001;
  assign mem[208] = 14'b00110110001100;
  assign mem[209] = 14'b01001000110011;
  assign mem[210] = 14'b00001001110001;
  assign mem[211] = 14'b00101010001100;
  assign mem[212] = 14'b01111000111010;
  assign mem[213] = 14'b00110101110011;
  assign mem[214] = 14'b00101111110100;
  assign mem[215] = 14'b00110100111100;
  assign mem[216] = 14'b00110111000110;
  assign mem[217] = 14'b01000101000010;
  assign mem[218] = 14'b10111010000111;
  assign mem[219] = 14'b01100001011000;
  assign mem[220] = 14'b00011011000010;
  assign mem[221] = 14'b00100111111110;
  assign mem[222] = 14'b10100001100100;
  assign mem[223] = 14'b01010011100000;
  assign mem[224] = 14'b01010010100110;
  assign mem[225] = 14'b00100010001110;
  assign mem[226] = 14'b10110100101010;
  assign mem[227] = 14'b01100000110111;
  assign mem[228] = 14'b00100110110010;
  assign mem[229] = 14'b10001000110100;
  assign mem[230] = 14'b01010100001011;
  assign mem[231] = 14'b01000000000101;
  assign mem[232] = 14'b01001000000001;
  assign mem[233] = 14'b10000110011101;
  assign mem[234] = 14'b10000000100010;
  assign mem[235] = 14'b00000010010000;
  assign mem[236] = 14'b01011000011000;
  assign mem[237] = 14'b10001000000000;
  assign mem[238] = 14'b00101000111101;
  assign mem[239] = 14'b01010100110000;
  assign mem[240] = 14'b10101000111100;
  assign mem[241] = 14'b00101110001111;
  assign mem[242] = 14'b10110001010010;
  assign mem[243] = 14'b01100001101001;
  assign mem[244] = 14'b00011010110011;
  assign mem[245] = 14'b01001101010111;
  assign mem[246] = 14'b10010101000100;
  assign mem[247] = 14'b00011101100000;
  assign mem[248] = 14'b00111010110100;
  assign mem[249] = 14'b00000000100111;
  assign mem[250] = 14'b10000000011011;
  assign mem[251] = 14'b00100000100000;
  assign mem[252] = 14'b00100111000110;
  assign mem[253] = 14'b00010110111101;
  assign mem[254] = 14'b10100100110110;
  assign mem[255] = 14'b10001000000101;
  assign mem[256] = 14'b01010111100001;
  assign mem[257] = 14'b00010001000101;
  assign mem[258] = 14'b00111011001000;
  assign mem[259] = 14'b01001110110001;
  assign mem[260] = 14'b00100000001010;
  assign mem[261] = 14'b10000011001111;
  assign mem[262] = 14'b10110010111000;
  assign mem[263] = 14'b10010110100111;
  assign mem[264] = 14'b00100000001011;
  assign mem[265] = 14'b10011010010110;
  assign mem[266] = 14'b01110011101101;
  assign mem[267] = 14'b00100111000000;
  assign mem[268] = 14'b01111011101110;
  assign mem[269] = 14'b10110101001010;
  assign mem[270] = 14'b00000101110011;
  assign mem[271] = 14'b01111100111001;
  assign mem[272] = 14'b00110000000001;
  assign mem[273] = 14'b10100001010110;
  assign mem[274] = 14'b00000000101000;
  assign mem[275] = 14'b10011100010100;
  assign mem[276] = 14'b10010000011101;
  assign mem[277] = 14'b01111100110011;
  assign mem[278] = 14'b01010111100011;
  assign mem[279] = 14'b00111111010011;
  assign mem[280] = 14'b01111011010110;
  assign mem[281] = 14'b00001010100100;
  assign mem[282] = 14'b10110001110100;
  assign mem[283] = 14'b01110011010011;
  assign mem[284] = 14'b01100101100101;
  assign mem[285] = 14'b01001101110101;
  assign mem[286] = 14'b00101001000100;
  assign mem[287] = 14'b00110110100000;
  assign mem[288] = 14'b10101011001100;
  assign mem[289] = 14'b01101101101110;
  assign mem[290] = 14'b01101001010001;
  assign mem[291] = 14'b10011011001101;
  assign mem[292] = 14'b01101111100011;
  assign mem[293] = 14'b00100100011010;
  assign mem[294] = 14'b00111100101100;
  assign mem[295] = 14'b01010101100001;
  assign mem[296] = 14'b01111010111001;
  assign mem[297] = 14'b01101100011101;
  assign mem[298] = 14'b01011001101001;
  assign mem[299] = 14'b01010111101101;
  assign mem[300] = 14'b10010100100001;
  assign mem[301] = 14'b10110100110000;
  assign mem[302] = 14'b10110000001101;
  assign mem[303] = 14'b00100111001110;
  assign mem[304] = 14'b01101000100001;
  assign mem[305] = 14'b00000110000010;
  assign mem[306] = 14'b01000101101110;
  assign mem[307] = 14'b00000001101001;
  assign mem[308] = 14'b00100000011100;
  assign mem[309] = 14'b10100011001011;
  assign mem[310] = 14'b00000001110111;
  assign mem[311] = 14'b00111101110011;
  assign mem[312] = 14'b01000100010010;
  assign mem[313] = 14'b10110011110001;
  assign mem[314] = 14'b00111001011000;
  assign mem[315] = 14'b10110010101111;
  assign mem[316] = 14'b00001011101110;
  assign mem[317] = 14'b00110010101000;
  assign mem[318] = 14'b00110000111101;
  assign mem[319] = 14'b00001011110010;
  assign mem[320] = 14'b00111110101101;
  assign mem[321] = 14'b10111010011001;
  assign mem[322] = 14'b10001111111010;
  assign mem[323] = 14'b01010100000010;
  assign mem[324] = 14'b10111001101001;
  assign mem[325] = 14'b10101100001010;
  assign mem[326] = 14'b00101100000010;
  assign mem[327] = 14'b00011100111011;
  assign mem[328] = 14'b01001101100110;
  assign mem[329] = 14'b01111111110101;
  assign mem[330] = 14'b00101010000000;
  assign mem[331] = 14'b01100000111101;
  assign mem[332] = 14'b01101010011110;
  assign mem[333] = 14'b00001110011110;
  assign mem[334] = 14'b00101101111000;
  assign mem[335] = 14'b01000011100111;
  assign mem[336] = 14'b10011110111111;
  assign mem[337] = 14'b01101110110001;
  assign mem[338] = 14'b01011110011111;
  assign mem[339] = 14'b10010011000010;
  assign mem[340] = 14'b10100011111100;
  assign mem[341] = 14'b10001011110110;
  assign mem[342] = 14'b00100110101000;
  assign mem[343] = 14'b01100001101111;
  assign mem[344] = 14'b00001011011000;
  assign mem[345] = 14'b01110110010001;
  assign mem[346] = 14'b01011110101000;
  assign mem[347] = 14'b10100011000000;
  assign mem[348] = 14'b10101100011100;
  assign mem[349] = 14'b00100110010100;
  assign mem[350] = 14'b00101011111011;
  assign mem[351] = 14'b00111011001011;
  assign mem[352] = 14'b00001110110001;
  assign mem[353] = 14'b10001100100110;
  assign mem[354] = 14'b00010011011100;
  assign mem[355] = 14'b10001001101111;
  assign mem[356] = 14'b10101100001001;
  assign mem[357] = 14'b10101111010010;
  assign mem[358] = 14'b01011100000110;
  assign mem[359] = 14'b01000011100101;
  assign mem[360] = 14'b01001000011111;
  assign mem[361] = 14'b00111011101011;
  assign mem[362] = 14'b10011001100010;
  assign mem[363] = 14'b01101110010000;
  assign mem[364] = 14'b01101010000010;
  assign mem[365] = 14'b10000111011110;
  assign mem[366] = 14'b01010110100011;
  assign mem[367] = 14'b01111000011011;
  assign mem[368] = 14'b00010101010001;
  assign mem[369] = 14'b10011001010100;
  assign mem[370] = 14'b00101110000101;
  assign mem[371] = 14'b10110000000001;
  assign mem[372] = 14'b10100000111101;
  assign mem[373] = 14'b10001110010100;
  assign mem[374] = 14'b00000111011110;
  assign mem[375] = 14'b01100101011001;
  assign mem[376] = 14'b00000001100101;
  assign mem[377] = 14'b00011101110111;
  assign mem[378] = 14'b10010100001011;
  assign mem[379] = 14'b00111000011000;
  assign mem[380] = 14'b10111011011101;
  assign mem[381] = 14'b10100100101000;
  assign mem[382] = 14'b00001100101100;
  assign mem[383] = 14'b10001011010011;
  assign mem[384] = 14'b00001001111101;
  assign mem[385] = 14'b01111111011111;
  assign mem[386] = 14'b01010010110011;
  assign mem[387] = 14'b10001110101000;
  assign mem[388] = 14'b00110110111000;
  assign mem[389] = 14'b10000001100010;
  assign mem[390] = 14'b01101110011100;
  assign mem[391] = 14'b01111011110010;
  assign mem[392] = 14'b00101111011100;
  assign mem[393] = 14'b01001010010111;
  assign mem[394] = 14'b00100001110011;
  assign mem[395] = 14'b00111101100001;
  assign mem[396] = 14'b00111010101011;
  assign mem[397] = 14'b10110000101010;
  assign mem[398] = 14'b01111000111011;
  assign mem[399] = 14'b01001100111010;
  assign mem[400] = 14'b10111010011100;
  assign mem[401] = 14'b00000110101000;
  assign mem[402] = 14'b01010110100010;
  assign mem[403] = 14'b01100001010100;
  assign mem[404] = 14'b10101101111011;
  assign mem[405] = 14'b01111001100010;
  assign mem[406] = 14'b10111011000110;
  assign mem[407] = 14'b00010001001001;
  assign mem[408] = 14'b00101101001010;
  assign mem[409] = 14'b10011100101011;
  assign mem[410] = 14'b00101000001001;
  assign mem[411] = 14'b00100011001010;
  assign mem[412] = 14'b00100100110000;
  assign mem[413] = 14'b00001100110101;
  assign mem[414] = 14'b00100111110110;
  assign mem[415] = 14'b10101100001000;
  assign mem[416] = 14'b01111001011001;
  assign mem[417] = 14'b00000010001000;
  assign mem[418] = 14'b00001001101001;
  assign mem[419] = 14'b00110001010101;
  assign mem[420] = 14'b01011100000001;
  assign mem[421] = 14'b10010000000011;
  assign mem[422] = 14'b01101011000111;
  assign mem[423] = 14'b00000001111000;
  assign mem[424] = 14'b01000100110101;
  assign mem[425] = 14'b00011100100001;
  assign mem[426] = 14'b10010110100011;
  assign mem[427] = 14'b01110000101110;
  assign mem[428] = 14'b10100000010101;
  assign mem[429] = 14'b10110010000001;
  assign mem[430] = 14'b00100110001001;
  assign mem[431] = 14'b10010101011010;
  assign mem[432] = 14'b10101110101000;
  assign mem[433] = 14'b00001001010111;
  assign mem[434] = 14'b00100000100101;
  assign mem[435] = 14'b10110011001001;
  assign mem[436] = 14'b01110001000001;
  assign mem[437] = 14'b01100000100001;
  assign mem[438] = 14'b01001011000001;
  assign mem[439] = 14'b10011011000110;
  assign mem[440] = 14'b10001100110010;
  assign mem[441] = 14'b01000110100010;
  assign mem[442] = 14'b10010011101111;
  assign mem[443] = 14'b10110001011000;
  assign mem[444] = 14'b10110110010110;
  assign mem[445] = 14'b01100000011110;
  assign mem[446] = 14'b01111100001110;
  assign mem[447] = 14'b10011000100110;
  assign mem[448] = 14'b01101011110000;
  assign mem[449] = 14'b10110101010011;
  assign mem[450] = 14'b00110010001101;
  assign mem[451] = 14'b10000100011001;
  assign mem[452] = 14'b10011010010001;
  assign mem[453] = 14'b00101100010011;
  assign mem[454] = 14'b10100010110110;
  assign mem[455] = 14'b00111010010100;
  assign mem[456] = 14'b01111100011001;
  assign mem[457] = 14'b00010110110001;
  assign mem[458] = 14'b10101001101001;
  assign mem[459] = 14'b01111110000101;
  assign mem[460] = 14'b00001101000000;
  assign mem[461] = 14'b00011001011100;
  assign mem[462] = 14'b00110101010010;
  assign mem[463] = 14'b01001100100100;
  assign mem[464] = 14'b10101001100111;
  assign mem[465] = 14'b01001111110111;
  assign mem[466] = 14'b10010101000111;
  assign mem[467] = 14'b01100010110101;
  assign mem[468] = 14'b01110100000111;
  assign mem[469] = 14'b00111111110011;
  assign mem[470] = 14'b00110000000000;
  assign mem[471] = 14'b10001010001111;
  assign mem[472] = 14'b10011001111101;
  assign mem[473] = 14'b10011110001010;
  assign mem[474] = 14'b01010010001011;
  assign mem[475] = 14'b10110010010101;
  assign mem[476] = 14'b01100110011100;
  assign mem[477] = 14'b00000100101111;
  assign mem[478] = 14'b00010110111001;
  assign mem[479] = 14'b00111100011111;
  assign mem[480] = 14'b01001100001001;
  assign mem[481] = 14'b01011010110101;
  assign mem[482] = 14'b10011100100001;
  assign mem[483] = 14'b01101011110010;
  assign mem[484] = 14'b00110011101111;
  assign mem[485] = 14'b01011100111011;
  assign mem[486] = 14'b10000110111101;
  assign mem[487] = 14'b01011011011100;
  assign mem[488] = 14'b00111100010000;
  assign mem[489] = 14'b00001110100000;
  assign mem[490] = 14'b01001101000101;
  assign mem[491] = 14'b10000101010010;
  assign mem[492] = 14'b00011101001111;
  assign mem[493] = 14'b00100010001000;
  assign mem[494] = 14'b01010111000011;
  assign mem[495] = 14'b01011011110111;
  assign mem[496] = 14'b00110110011001;
  assign mem[497] = 14'b10110101001101;
  assign mem[498] = 14'b10010100100111;
  assign mem[499] = 14'b01111111011001;
  assign mem[500] = 14'b00000000100011;
  assign mem[501] = 14'b00101000110001;
  assign mem[502] = 14'b01011101001011;
  assign mem[503] = 14'b01111110000000;
  assign mem[504] = 14'b00010000111000;
  assign mem[505] = 14'b10111100000111;
  assign mem[506] = 14'b10000011111100;
  assign mem[507] = 14'b00101111101100;
  assign mem[508] = 14'b00111011100101;
  assign mem[509] = 14'b10101100111001;
  assign mem[510] = 14'b01101001010000;
  assign mem[511] = 14'b10000100000110;
  assign mem[512] = 14'b00100100100100;
  assign mem[513] = 14'b01110111100011;
  assign mem[514] = 14'b00011101110110;
  assign mem[515] = 14'b10100111010101;
  assign mem[516] = 14'b00100001000101;
  assign mem[517] = 14'b10010110100101;
  assign mem[518] = 14'b01100100000010;
  assign mem[519] = 14'b01011110001100;
  assign mem[520] = 14'b00100001001100;
  assign mem[521] = 14'b01111000010101;
  assign mem[522] = 14'b00101001110111;
  assign mem[523] = 14'b01010000111111;
  assign mem[524] = 14'b01100001111110;
  assign mem[525] = 14'b01110100000000;
  assign mem[526] = 14'b00101000100101;
  assign mem[527] = 14'b01101010001011;
  assign mem[528] = 14'b10010000000110;
  assign mem[529] = 14'b10101001010101;
  assign mem[530] = 14'b00000100011000;
  assign mem[531] = 14'b10000110000111;
  assign mem[532] = 14'b00110011000110;
  assign mem[533] = 14'b01101001100001;
  assign mem[534] = 14'b00100100110010;
  assign mem[535] = 14'b00111011000011;
  assign mem[536] = 14'b01011111010110;
  assign mem[537] = 14'b01001001111100;
  assign mem[538] = 14'b01011100100110;
  assign mem[539] = 14'b00100111000001;
  assign mem[540] = 14'b10000111000000;
  assign mem[541] = 14'b10100000110001;
  assign mem[542] = 14'b01011111011011;
  assign mem[543] = 14'b10111101011111;
  assign mem[544] = 14'b00101110001110;
  assign mem[545] = 14'b10111111111111;
  assign mem[546] = 14'b10100000110100;
  assign mem[547] = 14'b01111110010110;
  assign mem[548] = 14'b00001100110001;
  assign mem[549] = 14'b00111110110101;
  assign mem[550] = 14'b00101000110010;
  assign mem[551] = 14'b00010110100100;
  assign mem[552] = 14'b01011100001011;
  assign mem[553] = 14'b10110111001000;
  assign mem[554] = 14'b00110011011100;
  assign mem[555] = 14'b00100101111000;
  assign mem[556] = 14'b01001111100010;
  assign mem[557] = 14'b01110001001010;
  assign mem[558] = 14'b01010001010101;
  assign mem[559] = 14'b01010010100001;
  assign mem[560] = 14'b10011011100100;
  assign mem[561] = 14'b00101010001110;
  assign mem[562] = 14'b01101000000000;
  assign mem[563] = 14'b00001011011111;
  assign mem[564] = 14'b00100011000011;
  assign mem[565] = 14'b10110110001000;
  assign mem[566] = 14'b00001101000001;
  assign mem[567] = 14'b00110000100011;
  assign mem[568] = 14'b01011101111100;
  assign mem[569] = 14'b01101010010001;
  assign mem[570] = 14'b00010001100110;
  assign mem[571] = 14'b01100011000011;
  assign mem[572] = 14'b01010010000010;
  assign mem[573] = 14'b10100010010111;
  assign mem[574] = 14'b10010110101010;
  assign mem[575] = 14'b01010010011110;
  assign mem[576] = 14'b00110110111001;
  assign mem[577] = 14'b10011000101001;
  assign mem[578] = 14'b00101111010001;
  assign mem[579] = 14'b00001100001011;
  assign mem[580] = 14'b10010011011001;
  assign mem[581] = 14'b00110101000000;
  assign mem[582] = 14'b01110100001101;
  assign mem[583] = 14'b00001010011100;
  assign mem[584] = 14'b10011111001000;
  assign mem[585] = 14'b01111110101111;
  assign mem[586] = 14'b01100101111111;
  assign mem[587] = 14'b01100110101000;
  assign mem[588] = 14'b10101001001111;
  assign mem[589] = 14'b01100101010010;
  assign mem[590] = 14'b10000001000111;
  assign mem[591] = 14'b01011001001111;
  assign mem[592] = 14'b10011000110100;
  assign mem[593] = 14'b00000111010011;
  assign mem[594] = 14'b01010101010110;
  assign mem[595] = 14'b01000101001001;
  assign mem[596] = 14'b10111011011111;
  assign mem[597] = 14'b00010010110101;
  assign mem[598] = 14'b01001110010111;
  assign mem[599] = 14'b01101100000110;
  assign mem[600] = 14'b01001111101000;
  assign mem[601] = 14'b00111011110011;
  assign mem[602] = 14'b01010110010101;
  assign mem[603] = 14'b10110100111011;
  assign mem[604] = 14'b00110110111110;
  assign mem[605] = 14'b01001100001011;
  assign mem[606] = 14'b01110011011100;
  assign mem[607] = 14'b00011110001011;
  assign mem[608] = 14'b01100111010111;
  assign mem[609] = 14'b00011000000101;
  assign mem[610] = 14'b10001000000100;
  assign mem[611] = 14'b00000100000100;
  assign mem[612] = 14'b00110100111001;
  assign mem[613] = 14'b01001010111000;
  assign mem[614] = 14'b01000100100111;
  assign mem[615] = 14'b01011001000001;
  assign mem[616] = 14'b01111011010111;
  assign mem[617] = 14'b00100001101011;
  assign mem[618] = 14'b01110010101001;
  assign mem[619] = 14'b00000011101100;
  assign mem[620] = 14'b10100110001011;
  assign mem[621] = 14'b10110100001110;
  assign mem[622] = 14'b00011101110010;
  assign mem[623] = 14'b01001010111001;
  assign mem[624] = 14'b10010100110111;
  assign mem[625] = 14'b01110001000111;
  assign mem[626] = 14'b10000010100010;
  assign mem[627] = 14'b01010000000001;
  assign mem[628] = 14'b10100110100110;
  assign mem[629] = 14'b00100100000111;
  assign mem[630] = 14'b00110100010010;
  assign mem[631] = 14'b10000101101100;
  assign mem[632] = 14'b00001011000011;
  assign mem[633] = 14'b00010001000000;
  assign mem[634] = 14'b01001101001000;
  assign mem[635] = 14'b00001010100110;
  assign mem[636] = 14'b10100000000101;
  assign mem[637] = 14'b00000000010010;
  assign mem[638] = 14'b01011000110100;
  assign mem[639] = 14'b00001111000000;
  assign mem[640] = 14'b01000101101011;
  assign mem[641] = 14'b01111100010101;
  assign mem[642] = 14'b00000011100010;
  assign mem[643] = 14'b00100110010011;
  assign mem[644] = 14'b00000000000110;
  assign mem[645] = 14'b10001010101010;
  assign mem[646] = 14'b00000101000000;
  assign mem[647] = 14'b01100010011010;
  assign mem[648] = 14'b10001100000011;
  assign mem[649] = 14'b10001000011111;
  assign mem[650] = 14'b00101100100100;
  assign mem[651] = 14'b00101110100101;
  assign mem[652] = 14'b00011010101011;
  assign mem[653] = 14'b01010100100000;
  assign mem[654] = 14'b01001110011001;
  assign mem[655] = 14'b10011010010100;
  assign mem[656] = 14'b10011000111110;
  assign mem[657] = 14'b00101110011000;
  assign mem[658] = 14'b00011101101011;
  assign mem[659] = 14'b01101001001001;
  assign mem[660] = 14'b01000001010111;
  assign mem[661] = 14'b01010010101010;
  assign mem[662] = 14'b10011101100100;
  assign mem[663] = 14'b01110111111111;
  assign mem[664] = 14'b01111100000101;
  assign mem[665] = 14'b10001000101000;
  assign mem[666] = 14'b01011000111110;
  assign mem[667] = 14'b00110110000101;
  assign mem[668] = 14'b01000001001111;
  assign mem[669] = 14'b01011001110011;
  assign mem[670] = 14'b01010110111001;
  assign mem[671] = 14'b00110100110010;
  assign mem[672] = 14'b01010001101011;
  assign mem[673] = 14'b00001110111000;
  assign mem[674] = 14'b01000011011111;
  assign mem[675] = 14'b10011001010010;
  assign mem[676] = 14'b01000100000100;
  assign mem[677] = 14'b00110000010000;
  assign mem[678] = 14'b10101101101110;
  assign mem[679] = 14'b00001101001000;
  assign mem[680] = 14'b01100001110001;
  assign mem[681] = 14'b00000111100110;
  assign mem[682] = 14'b01011101110000;
  assign mem[683] = 14'b00010100111110;
  assign mem[684] = 14'b10100010001110;
  assign mem[685] = 14'b01011110000001;
  assign mem[686] = 14'b01001010111110;
  assign mem[687] = 14'b01010101110001;
  assign mem[688] = 14'b01000110010010;
  assign mem[689] = 14'b01000001100001;
  assign mem[690] = 14'b00100100000010;
  assign mem[691] = 14'b01100101111001;
  assign mem[692] = 14'b00010111000011;
  assign mem[693] = 14'b01100011100100;
  assign mem[694] = 14'b10001101000101;
  assign mem[695] = 14'b01111101100101;
  assign mem[696] = 14'b00011001011001;
  assign mem[697] = 14'b01101101101100;
  assign mem[698] = 14'b01001010000100;
  assign mem[699] = 14'b01011001100010;
  assign mem[700] = 14'b01111100010100;
  assign mem[701] = 14'b01100011001111;
  assign mem[702] = 14'b01100101011110;
  assign mem[703] = 14'b01101100000101;
  assign mem[704] = 14'b10110010001101;
  assign mem[705] = 14'b01110100111111;
  assign mem[706] = 14'b10011111011010;
  assign mem[707] = 14'b10011110101011;
  assign mem[708] = 14'b01110111110010;
  assign mem[709] = 14'b01110110000100;
  assign mem[710] = 14'b10110011110101;
  assign mem[711] = 14'b00011000001010;
  assign mem[712] = 14'b01100110101011;
  assign mem[713] = 14'b10011111010111;
  assign mem[714] = 14'b00100011011001;
  assign mem[715] = 14'b01110010011111;
  assign mem[716] = 14'b01011011000000;
  assign mem[717] = 14'b10110010000100;
  assign mem[718] = 14'b10110100111101;
  assign mem[719] = 14'b10010111111010;
  assign mem[720] = 14'b00100011001011;
  assign mem[721] = 14'b10101110111111;
  assign mem[722] = 14'b01010011101100;
  assign mem[723] = 14'b01110011110000;
  assign mem[724] = 14'b00101100101101;
  assign mem[725] = 14'b00111110100011;
  assign mem[726] = 14'b10001111111111;
  assign mem[727] = 14'b00000111100100;
  assign mem[728] = 14'b01110101100110;
  assign mem[729] = 14'b10010011000001;
  assign mem[730] = 14'b10111111001011;
  assign mem[731] = 14'b01100000001101;
  assign mem[732] = 14'b10001101000001;
  assign mem[733] = 14'b00100001001001;
  assign mem[734] = 14'b10100000001111;
  assign mem[735] = 14'b00100111010111;
  assign mem[736] = 14'b10010100111101;
  assign mem[737] = 14'b00111011110000;
  assign mem[738] = 14'b10000111100010;
  assign mem[739] = 14'b10110010011011;
  assign mem[740] = 14'b10101010001000;
  assign mem[741] = 14'b01001010011010;
  assign mem[742] = 14'b10110000100111;
  assign mem[743] = 14'b01000000000001;
  assign mem[744] = 14'b00100101101110;
  assign mem[745] = 14'b01100101100000;
  assign mem[746] = 14'b10011011100001;
  assign mem[747] = 14'b10100100111010;
  assign mem[748] = 14'b00001100101000;
  assign mem[749] = 14'b00101110110111;
  assign mem[750] = 14'b00100001010010;
  assign mem[751] = 14'b01000010111110;
  assign mem[752] = 14'b10111100101110;
  assign mem[753] = 14'b01110100010101;
  assign mem[754] = 14'b01010000001100;
  assign mem[755] = 14'b01111011101011;
  assign mem[756] = 14'b00000011110101;
  assign mem[757] = 14'b01011101010110;
  assign mem[758] = 14'b01001100001010;
  assign mem[759] = 14'b01110001111100;
  assign mem[760] = 14'b01110110001000;
  assign mem[761] = 14'b10100100101011;
  assign mem[762] = 14'b10011011100000;
  assign mem[763] = 14'b10001101110011;
  assign mem[764] = 14'b00100001000001;
  assign mem[765] = 14'b00111010001001;
  assign mem[766] = 14'b10100000101101;
  assign mem[767] = 14'b10011100100110;
  assign mem[768] = 14'b10010101101010;
  assign mem[769] = 14'b10001011100110;
  assign mem[770] = 14'b10101101000010;
  assign mem[771] = 14'b10010100011010;
  assign mem[772] = 14'b00000100100110;
  assign mem[773] = 14'b01001001100111;
  assign mem[774] = 14'b00110100111111;
  assign mem[775] = 14'b00010101100001;
  assign mem[776] = 14'b10001101110000;
  assign mem[777] = 14'b10011111001101;
  assign mem[778] = 14'b01000111011001;
  assign mem[779] = 14'b10101010001010;
  assign mem[780] = 14'b10011010110101;
  assign mem[781] = 14'b01101100001011;
  assign mem[782] = 14'b00000000110101;
  assign mem[783] = 14'b01001000101101;
  assign mem[784] = 14'b00000110110111;
  assign mem[785] = 14'b10100000001101;
  assign mem[786] = 14'b01101101110100;
  assign mem[787] = 14'b10011111011111;
  assign mem[788] = 14'b10000010010111;
  assign mem[789] = 14'b00010001110101;
  assign mem[790] = 14'b00100111111100;
  assign mem[791] = 14'b01110110110001;
  assign mem[792] = 14'b01111111010110;
  assign mem[793] = 14'b10100110000110;
  assign mem[794] = 14'b10000111001000;
  assign mem[795] = 14'b10011001101000;
  assign mem[796] = 14'b01111100001111;
  assign mem[797] = 14'b10101111101101;
  assign mem[798] = 14'b00100001010011;
  assign mem[799] = 14'b01011010000101;
  assign mem[800] = 14'b10100001100111;
  assign mem[801] = 14'b10011000110101;
  assign mem[802] = 14'b00101010011110;
  assign mem[803] = 14'b00010110001011;
  assign mem[804] = 14'b01000110110011;
  assign mem[805] = 14'b00111100000100;
  assign mem[806] = 14'b00111111100010;
  assign mem[807] = 14'b01000011000101;
  assign mem[808] = 14'b10110110001001;
  assign mem[809] = 14'b10110100000101;
  assign mem[810] = 14'b10110001011001;
  assign mem[811] = 14'b01000011011001;
  assign mem[812] = 14'b01001100000101;
  assign mem[813] = 14'b10111110011010;
  assign mem[814] = 14'b00011001001011;
  assign mem[815] = 14'b10101010001100;
  assign mem[816] = 14'b10110011100001;
  assign mem[817] = 14'b10001010000001;
  assign mem[818] = 14'b00100101011001;
  assign mem[819] = 14'b00000000001111;
  assign mem[820] = 14'b10101001001110;
  assign mem[821] = 14'b01001110001011;
  assign mem[822] = 14'b00000000010001;
  assign mem[823] = 14'b00001000110101;
  assign mem[824] = 14'b01011100000011;
  assign mem[825] = 14'b10111110010001;
  assign mem[826] = 14'b10101100110010;
  assign mem[827] = 14'b10100010101100;
  assign mem[828] = 14'b10001010110101;
  assign mem[829] = 14'b00111110000110;
  assign mem[830] = 14'b10101011100101;
  assign mem[831] = 14'b01101111011010;
  assign mem[832] = 14'b01011011010000;
  assign mem[833] = 14'b10100011110010;
  assign mem[834] = 14'b10000010010010;
  assign mem[835] = 14'b01011110010011;
  assign mem[836] = 14'b01101100110100;
  assign mem[837] = 14'b00011000100110;
  assign mem[838] = 14'b10101010111000;
  assign mem[839] = 14'b00011111100100;
  assign mem[840] = 14'b00100110100001;
  assign mem[841] = 14'b01111111111111;
  assign mem[842] = 14'b00000110000000;
  assign mem[843] = 14'b00101001010010;
  assign mem[844] = 14'b00101010101001;
  assign mem[845] = 14'b01010100010111;
  assign mem[846] = 14'b00100001111111;
  assign mem[847] = 14'b10010010110100;
  assign mem[848] = 14'b10111011010011;
  assign mem[849] = 14'b01111101100011;
  assign mem[850] = 14'b01000100010111;
  assign mem[851] = 14'b01100111010011;
  assign mem[852] = 14'b01001110010010;
  assign mem[853] = 14'b10111000100100;
  assign mem[854] = 14'b10001110101011;
  assign mem[855] = 14'b10110010100011;
  assign mem[856] = 14'b00000001101000;
  assign mem[857] = 14'b01100011001100;
  assign mem[858] = 14'b10010110101011;
  assign mem[859] = 14'b01101001100101;
  assign mem[860] = 14'b10111101001110;
  assign mem[861] = 14'b01010111110001;
  assign mem[862] = 14'b10101010110111;
  assign mem[863] = 14'b00001000011101;
  assign mem[864] = 14'b00000010000111;
  assign mem[865] = 14'b00101111100001;
  assign mem[866] = 14'b01110000100000;
  assign mem[867] = 14'b01100101111110;
  assign mem[868] = 14'b01001111011101;
  assign mem[869] = 14'b10111101101000;
  assign mem[870] = 14'b00001101001010;
  assign mem[871] = 14'b01000000100001;
  assign mem[872] = 14'b01111000000101;
  assign mem[873] = 14'b10101101000111;
  assign mem[874] = 14'b10000011101010;
  assign mem[875] = 14'b00001111110000;
  assign mem[876] = 14'b00101010100101;
  assign mem[877] = 14'b10110111111100;
  assign mem[878] = 14'b01011110101010;
  assign mem[879] = 14'b00010001001101;
  assign mem[880] = 14'b00011110011110;
  assign mem[881] = 14'b10000011101000;
  assign mem[882] = 14'b01011000111000;
  assign mem[883] = 14'b01101011011100;
  assign mem[884] = 14'b10111011100101;
  assign mem[885] = 14'b10011101011111;
  assign mem[886] = 14'b01010011010111;
  assign mem[887] = 14'b00001110011111;
  assign mem[888] = 14'b00011011101010;
  assign mem[889] = 14'b00000100010001;
  assign mem[890] = 14'b10000010111001;
  assign mem[891] = 14'b00100011011111;
  assign mem[892] = 14'b01010001101001;
  assign mem[893] = 14'b10100000101011;
  assign mem[894] = 14'b00000001110100;
  assign mem[895] = 14'b10111000011111;
  assign mem[896] = 14'b00000001011011;
  assign mem[897] = 14'b10110110110011;
  assign mem[898] = 14'b00001011110101;
  assign mem[899] = 14'b00010100011000;
  assign mem[900] = 14'b01110101100100;
  assign mem[901] = 14'b01100100110011;
  assign mem[902] = 14'b01111101100000;
  assign mem[903] = 14'b01111111011010;
  assign mem[904] = 14'b01110100100000;
  assign mem[905] = 14'b01000001011111;
  assign mem[906] = 14'b00000100110101;
  assign mem[907] = 14'b00100100001110;
  assign mem[908] = 14'b00100011110100;
  assign mem[909] = 14'b10100010011001;
  assign mem[910] = 14'b10110101110111;
  assign mem[911] = 14'b10010100001001;
  assign mem[912] = 14'b10111111001110;
  assign mem[913] = 14'b10100101100010;
  assign mem[914] = 14'b10010101100001;
  assign mem[915] = 14'b01111011101000;
  assign mem[916] = 14'b10100010000000;
  assign mem[917] = 14'b10011010100001;
  assign mem[918] = 14'b10111111010100;
  assign mem[919] = 14'b01110000001011;
  assign mem[920] = 14'b00111101010100;
  assign mem[921] = 14'b00110001110100;
  assign mem[922] = 14'b00000101101111;
  assign mem[923] = 14'b00100000011101;
  assign mem[924] = 14'b00000101010000;
  assign mem[925] = 14'b01010100001000;
  assign mem[926] = 14'b01010111111111;
  assign mem[927] = 14'b10000110010100;
  assign mem[928] = 14'b01001000001101;
  assign mem[929] = 14'b00011011101111;
  assign mem[930] = 14'b10001010100010;
  assign mem[931] = 14'b00000111000011;
  assign mem[932] = 14'b01011111011100;
  assign mem[933] = 14'b00010100100101;
  assign mem[934] = 14'b01100001100110;
  assign mem[935] = 14'b10001001011011;
  assign mem[936] = 14'b01011100001000;
  assign mem[937] = 14'b01110001110011;
  assign mem[938] = 14'b00110000111100;
  assign mem[939] = 14'b10110100101100;
  assign mem[940] = 14'b01001101110001;
  assign mem[941] = 14'b10111110000001;
  assign mem[942] = 14'b01110011001011;
  assign mem[943] = 14'b00010101010110;
  assign mem[944] = 14'b10111101100010;
  assign mem[945] = 14'b10100101111011;
  assign mem[946] = 14'b00111011100001;
  assign mem[947] = 14'b01010000011101;
  assign mem[948] = 14'b01100010011100;
  assign mem[949] = 14'b00101001001110;
  assign mem[950] = 14'b01000001100101;
  assign mem[951] = 14'b00010110001010;
  assign mem[952] = 14'b10011101010001;
  assign mem[953] = 14'b01000000111100;
  assign mem[954] = 14'b10000010110101;
  assign mem[955] = 14'b10000111000100;
  assign mem[956] = 14'b10100011001101;
  assign mem[957] = 14'b00001101110010;
  assign mem[958] = 14'b01111111011110;
  assign mem[959] = 14'b10011110111101;
  assign mem[960] = 14'b10011000100011;
  assign mem[961] = 14'b10111110011111;
  assign mem[962] = 14'b00000111001011;
  assign mem[963] = 14'b00101110010110;
  assign mem[964] = 14'b00110001011110;
  assign mem[965] = 14'b00000110010101;
  assign mem[966] = 14'b01001110001000;
  assign mem[967] = 14'b10010001011111;
  assign mem[968] = 14'b01100100000100;
  assign mem[969] = 14'b10001100011010;
  assign mem[970] = 14'b00011000001111;
  assign mem[971] = 14'b01111111101111;
  assign mem[972] = 14'b00111000101110;
  assign mem[973] = 14'b10101000001110;
  assign mem[974] = 14'b10010000110001;
  assign mem[975] = 14'b00001010111100;
  assign mem[976] = 14'b10000101111101;
  assign mem[977] = 14'b10010100100100;
  assign mem[978] = 14'b01100111100110;
  assign mem[979] = 14'b10110010101101;
  assign mem[980] = 14'b10110101001011;
  assign mem[981] = 14'b01011011011010;
  assign mem[982] = 14'b00111101101110;
  assign mem[983] = 14'b01001010100111;
  assign mem[984] = 14'b10111010100101;
  assign mem[985] = 14'b00010110100110;
  assign mem[986] = 14'b01011110000010;
  assign mem[987] = 14'b00110100111010;
  assign mem[988] = 14'b10110011001110;
  assign mem[989] = 14'b01010010111110;
  assign mem[990] = 14'b01010101100100;
  assign mem[991] = 14'b00001000101001;
  assign mem[992] = 14'b10010100000010;
  assign mem[993] = 14'b00101000011010;
  assign mem[994] = 14'b00010110010111;
  assign mem[995] = 14'b00101010110101;
  assign mem[996] = 14'b00000111011001;
  assign mem[997] = 14'b10110001110111;
  assign mem[998] = 14'b01001010001001;
  assign mem[999] = 14'b00001101000100;
  assign mem[1000] = 14'b00111111011110;
  assign mem[1001] = 14'b10100110101010;
  assign mem[1002] = 14'b01111000101111;
  assign mem[1003] = 14'b10110111101000;
  assign mem[1004] = 14'b01010110011110;
  assign mem[1005] = 14'b00000100111000;
  assign mem[1006] = 14'b01000011010011;
  assign mem[1007] = 14'b01000011111111;
  assign mem[1008] = 14'b01011010000100;
  assign mem[1009] = 14'b10000111100111;
  assign mem[1010] = 14'b10000010111101;
  assign mem[1011] = 14'b01111111111011;
  assign mem[1012] = 14'b00000000000101;
  assign mem[1013] = 14'b01110011100011;
  assign mem[1014] = 14'b01000100001011;
  assign mem[1015] = 14'b00010010000000;
  assign mem[1016] = 14'b01010100101101;
  assign mem[1017] = 14'b01010001101111;
  assign mem[1018] = 14'b01100101001001;
  assign mem[1019] = 14'b00000110110100;
  assign mem[1020] = 14'b01110110001111;
  assign mem[1021] = 14'b10000110011011;
  assign mem[1022] = 14'b01100001010101;
  assign mem[1023] = 14'b10000000100110;
  always@(*)
  begin
    data_out_t <= mem[addr_f];
  end
  wire [13:0] data_out_reg [n_outreg:0];
  generate if (n_outreg > 0)
  begin
    for( i=n_outreg-1; i >= 1; i=i-1)
    begin: data_out_reg_stage
      mgc_generic_reg #(
        .width(14),
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_data_out_reg (
        .d(data_out_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(data_out_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(14),
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_data_out_reg_init (
      .d(data_out_t),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(data_out_reg[0])
    );
    assign data_out = data_out_reg[n_outreg-1];
  end
  else
  begin
    assign data_out = data_out_t;
  end
  endgenerate
endmodule
module stagemgc_rom_sync_regout_10_1024_62_1_0_0_1_0_1_0_0_0_1_60 (addr, data_out,
    clk, s_rst, a_rst, en
);
  input [9:0]addr ;
  output [61:0]data_out ;
  input clk ;
  input s_rst ;
  input a_rst ;
  input en ;
  parameter n_width = 62;
  parameter n_size = 1024;
  parameter n_numports = 1;
  parameter n_addr_w = 10;
  parameter n_inreg = 0;
  parameter n_outreg = 1;
  wire [9:0] addr_f;
  wire [9:0] addr_reg [n_inreg:0];
  genvar i;
  generate if (n_inreg > 0)
  begin
    for( i=n_inreg-1; i >= 1; i=i-1)
    begin: addr_reg_stage
      mgc_generic_reg #(
        .width(10),
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_addr_reg (
        .d(addr_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(addr_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(10),
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_addr_reg_init (
      .d(addr),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(addr_reg[0])
    );
    assign addr_f = addr_reg[n_inreg-1];
  end
  else
  begin
    assign addr_f = addr;
  end
  endgenerate
  wire [61:0] mem [1023:0];
  reg [61:0] data_out_t;
  assign mem[0] = 62'b00000000000000000000000000000000000000000000000000000000000000;
  assign mem[1] = 62'b11111111110000000000000000000000000000000000000000000000000000;
  assign mem[2] = 62'b11111111100110101000001001111001100110011111110011101111001101;
  assign mem[3] = 62'b11111111100110101000001001111001100110011111110011101111001101;
  assign mem[4] = 62'b11111111011000011111011110001010100110101011101010100101100011;
  assign mem[5] = 62'b11111111101101100100000110101111001111001100101000110101000110;
  assign mem[6] = 62'b11111111101101100100000110101111001111001100101000110101000110;
  assign mem[7] = 62'b11111111011000011111011110001010100110101011101010100101100011;
  assign mem[8] = 62'b11111111001000111110001011100000111100011010011010011000001011;
  assign mem[9] = 62'b11111111101111011000101001011111001111111101110101110010110000;
  assign mem[10] = 62'b11111111101010100110110110011000101001000011101010000110100011;
  assign mem[11] = 62'b11111111100001110001110011101100111001101011100110100011001000;
  assign mem[12] = 62'b11111111100001110001110011101100111001101011100110100011001000;
  assign mem[13] = 62'b11111111101010100110110110011000101001000011101010000110100011;
  assign mem[14] = 62'b11111111101111011000101001011111001111111101110101110010110000;
  assign mem[15] = 62'b11111111001000111110001011100000111100011010011010011000001011;
  assign mem[16] = 62'b11111110111001000101111010011010111100001010011011010000101100;
  assign mem[17] = 62'b11111111101111110110001000110110100011110100010010010100100110;
  assign mem[18] = 62'b11111111101000101111001000000001101011000101010001011101000001;
  assign mem[19] = 62'b11111111100100010011001111001100100101000010010001110111010110;
  assign mem[20] = 62'b11111111011110001010110101110100111000000001101111011000111011;
  assign mem[21] = 62'b11111111101100001110001011001011110001100000001011110110110001;
  assign mem[22] = 62'b11111111101110100111110100000101010110110001100010110111011010;
  assign mem[23] = 62'b11111111010010100101000000011000101110110101011001111100000110;
  assign mem[24] = 62'b11111111010010100101000000011000101110110101011001111100000110;
  assign mem[25] = 62'b11111111101110100111110100000101010110110001100010110111011010;
  assign mem[26] = 62'b11111111101100001110001011001011110001100000001011110110110001;
  assign mem[27] = 62'b11111111011110001010110101110100111000000001101111011000111011;
  assign mem[28] = 62'b11111111100100010011001111001100100101000010010001110111010110;
  assign mem[29] = 62'b11111111101000101111001000000001101011000101010001011101000001;
  assign mem[30] = 62'b11111111101111110110001000110110100011110100010010010100100110;
  assign mem[31] = 62'b11111110111001000101111010011010111100001010011011010000101100;
  assign mem[32] = 62'b11111110101001000111110110010111110001000011011101100000010100;
  assign mem[33] = 62'b11111111101111111101100010000111100011011110010110110101111110;
  assign mem[34] = 62'b11111111100111101101011101111100100010011010101010111110101111;
  assign mem[35] = 62'b11111111100101011111010110100100110100100011001110110010100000;
  assign mem[36] = 62'b11111111011011010111010001000000001001111000010101110011000000;
  assign mem[37] = 62'b11111111101100111011010111101011110100001111001100011101110011;
  assign mem[38] = 62'b11111111101110001000010010000100000100111101101000011011100101;
  assign mem[39] = 62'b11111111010101100011111001101001110101101010110001111111011101;
  assign mem[40] = 62'b11111111001111000110011111100101111011001000010101111100011011;
  assign mem[41] = 62'b11111111101111000010100111111011111011100100100011000011010111;
  assign mem[42] = 62'b11111111101011011100101000001101000101000110010110111000111110;
  assign mem[43] = 62'b11111111100000011100111000011110011001001000101111111111101110;
  assign mem[44] = 62'b11111111100011000011111111011111111100111000010111000000110101;
  assign mem[45] = 62'b11111111101001101100111110000001000111111100111000011101000001;
  assign mem[46] = 62'b11111111101111101001110101010101111111000010001010010100010111;
  assign mem[47] = 62'b11111111000010110010000001000001101110100011100110000100111010;
  assign mem[48] = 62'b11111111000010110010000001000001101110100011100110000100111010;
  assign mem[49] = 62'b11111111101111101001110101010101111111000010001010010100010111;
  assign mem[50] = 62'b11111111101001101100111110000001000111111100111000011101000001;
  assign mem[51] = 62'b11111111100011000011111111011111111100111000010111000000110101;
  assign mem[52] = 62'b11111111100000011100111000011110011001001000101111111111101110;
  assign mem[53] = 62'b11111111101011011100101000001101000101000110010110111000111110;
  assign mem[54] = 62'b11111111101111000010100111111011111011100100100011000011010111;
  assign mem[55] = 62'b11111111001111000110011111100101111011001000010101111100011011;
  assign mem[56] = 62'b11111111010101100011111001101001110101101010110001111111011101;
  assign mem[57] = 62'b11111111101110001000010010000100000100111101101000011011100101;
  assign mem[58] = 62'b11111111101100111011010111101011110100001111001100011101110011;
  assign mem[59] = 62'b11111111011011010111010001000000001001111000010101110011000000;
  assign mem[60] = 62'b11111111100101011111010110100100110100100011001110110010100000;
  assign mem[61] = 62'b11111111100111101101011101111100100010011010101010111110101111;
  assign mem[62] = 62'b11111111101111111101100010000111100011011110010110110101111110;
  assign mem[63] = 62'b11111110101001000111110110010111110001000011011101100000010100;
  assign mem[64] = 62'b11111110011001001000010101010111110111101000110110011001111110;
  assign mem[65] = 62'b11111111101111111111011000100001100000100001001100110100001101;
  assign mem[66] = 62'b11111111100111001011010000100000110111111011111111111110010110;
  assign mem[67] = 62'b11111111100110000100001011011101010101000111010010110011011111;
  assign mem[68] = 62'b11111111011001111011110111100101000011101010001110110110001010;
  assign mem[69] = 62'b11111111101101010000010011010011010001010011011100100100111010;
  assign mem[70] = 62'b11111111101101110110110001001110110110110011001100001000111100;
  assign mem[71] = 62'b11111111010111000010001000010100110000111110100100010110011111;
  assign mem[72] = 62'b11111111001100000010111000001001101010011111100100111101100011;
  assign mem[73] = 62'b11111111101111001110001111001110101100011001001110010110001001;
  assign mem[74] = 62'b11111111101011000010010000101001011000000101010000001000000000;
  assign mem[75] = 62'b11111111100001000111101011001101010100000110110100101100100011;
  assign mem[76] = 62'b11111111100010011011010000010101001100110111010001001011011111;
  assign mem[77] = 62'b11111111101010001010011010011110100000010001100010011110000010;
  assign mem[78] = 62'b11111111101111100001110110010011111010011100010100101110101001;
  assign mem[79] = 62'b11111111000101111000100001010001000100100010110011111111000110;
  assign mem[80] = 62'b11111110111111010101100100111001010110101010010111001100001110;
  assign mem[81] = 62'b11111111101111110000100110010001110000111000011001111111010011;
  assign mem[82] = 62'b11111111101001001110100010001001001001100100100110001111111011;
  assign mem[83] = 62'b11111111100011101011111111101000101001001000000101000010111001;
  assign mem[84] = 62'b11111111011111100010111010010011011011111110001001101010111010;
  assign mem[85] = 62'b11111111101011110101111100000010101100011011111001010100101010;
  assign mem[86] = 62'b11111111101110110101110100000011100111011010000100100101100011;
  assign mem[87] = 62'b11111111010001000100011101001001100010101100011111011001110111;
  assign mem[88] = 62'b11111111010100000100110101110010010100000101110110011000000001;
  assign mem[89] = 62'b11111111101110011000101000100011101100010010001110000100010010;
  assign mem[90] = 62'b11111111101100100101010100101100100001001101000001000111110101;
  assign mem[91] = 62'b11111111011100110001100110111010011001001100011100010001011110;
  assign mem[92] = 62'b11111111100100111001101100101010111011111000111110010111101001;
  assign mem[93] = 62'b11111111101000001110110000111000001011111111111001011101101110;
  assign mem[94] = 62'b11111111101111111010011100110110101101000000011000100000111010;
  assign mem[95] = 62'b11111110110010110101010010000010010010110011100001100111110110;
  assign mem[96] = 62'b11111110110010110101010010000010010010110011100001100111110110;
  assign mem[97] = 62'b11111111101111111010011100110110101101000000011000100000111010;
  assign mem[98] = 62'b11111111101000001110110000111000001011111111111001011101101110;
  assign mem[99] = 62'b11111111100100111001101100101010111011111000111110010111101001;
  assign mem[100] = 62'b11111111011100110001100110111010011001001100011100010001011110;
  assign mem[101] = 62'b11111111101100100101010100101100100001001101000001000111110101;
  assign mem[102] = 62'b11111111101110011000101000100011101100010010001110000100010010;
  assign mem[103] = 62'b11111111010100000100110101110010010100000101110110011000000001;
  assign mem[104] = 62'b11111111010001000100011101001001100010101100011111011001110111;
  assign mem[105] = 62'b11111111101110110101110100000011100111011010000100100101100011;
  assign mem[106] = 62'b11111111101011110101111100000010101100011011111001010100101010;
  assign mem[107] = 62'b11111111011111100010111010010011011011111110001001101010111010;
  assign mem[108] = 62'b11111111100011101011111111101000101001001000000101000010111001;
  assign mem[109] = 62'b11111111101001001110100010001001001001100100100110001111111011;
  assign mem[110] = 62'b11111111101111110000100110010001110000111000011001111111010011;
  assign mem[111] = 62'b11111110111111010101100100111001010110101010010111001100001110;
  assign mem[112] = 62'b11111111000101111000100001010001000100100010110011111111000110;
  assign mem[113] = 62'b11111111101111100001110110010011111010011100010100101110101001;
  assign mem[114] = 62'b11111111101010001010011010011110100000010001100010011110000010;
  assign mem[115] = 62'b11111111100010011011010000010101001100110111010001001011011111;
  assign mem[116] = 62'b11111111100001000111101011001101010100000110110100101100100011;
  assign mem[117] = 62'b11111111101011000010010000101001011000000101010000001000000000;
  assign mem[118] = 62'b11111111101111001110001111001110101100011001001110010110001001;
  assign mem[119] = 62'b11111111001100000010111000001001101010011111100100111101100011;
  assign mem[120] = 62'b11111111010111000010001000010100110000111110100100010110011111;
  assign mem[121] = 62'b11111111101101110110110001001110110110110011001100001000111100;
  assign mem[122] = 62'b11111111101101010000010011010011010001010011011100100100111010;
  assign mem[123] = 62'b11111111011001111011110111100101000011101010001110110110001010;
  assign mem[124] = 62'b11111111100110000100001011011101010101000111010010110011011111;
  assign mem[125] = 62'b11111111100111001011010000100000110111111011111111111110010110;
  assign mem[126] = 62'b11111111101111111111011000100001100000100001001100110100001101;
  assign mem[127] = 62'b11111110011001001000010101010111110111101000110110011001111110;
  assign mem[128] = 62'b11111110001001001000011101000111111100110111101100011110000100;
  assign mem[129] = 62'b11111111101111111111110110001000010110100110111001001011011011;
  assign mem[130] = 62'b11111111100110111001110100010001010100111010101010100010101111;
  assign mem[131] = 62'b11111111100110010110010001100100100101111100000111100000111101;
  assign mem[132] = 62'b11111111011001001101110010101001100011101111001001001111010111;
  assign mem[133] = 62'b11111111101101011010010110000101110011110010011110011010001011;
  assign mem[134] = 62'b11111111101101101101100101001001100010001110001010000010011011;
  assign mem[135] = 62'b11111111010111110000111010100100110001000111011100110011100111;
  assign mem[136] = 62'b11111111001010100000101010000000100101101100000000010001010001;
  assign mem[137] = 62'b11111111101111010011100110000000111011000010110010111100101101;
  assign mem[138] = 62'b11111111101010110100101011110010011110001000011101010100010001;
  assign mem[139] = 62'b11111111100001011100110100110101100011110111101101101101001001;
  assign mem[140] = 62'b11111111100010000110100111100110011001001100111110101101011001;
  assign mem[141] = 62'b11111111101010011000110000100100011011000000101111101011100010;
  assign mem[142] = 62'b11111111101111011101011001100110100011101000010010000001110111;
  assign mem[143] = 62'b11111111000111011011011101100111011110010100001011111100110001;
  assign mem[144] = 62'b11111110111100001101111000010111000111100111101100001011010101;
  assign mem[145] = 62'b11111111101111110011100001010111111101011011011010011001111011;
  assign mem[146] = 62'b11111111101000111110111100110010100011111011111001010000001101;
  assign mem[147] = 62'b11111111100011111111101101100101010011010001010101011011010100;
  assign mem[148] = 62'b11111111011110110111000001100101010010111011110111100011010110;
  assign mem[149] = 62'b11111111101100000010001100010000100110011100100101010101001001;
  assign mem[150] = 62'b11111111101110101110111101100011001000110111110000101101110100;
  assign mem[151] = 62'b11111111010001110100110100010000111111010011001101101100111110;
  assign mem[152] = 62'b11111111010011010101000001000011000010111000011000000101010010;
  assign mem[153] = 62'b11111111101110100000010111101110101011010011001101000100001101;
  assign mem[154] = 62'b11111111101100011001111000101100110100100010000111001110011011;
  assign mem[155] = 62'b11111111011101011110010111011101011011100001101110001110001001;
  assign mem[156] = 62'b11111111100100100110100100010010011011100110110000100100111001;
  assign mem[157] = 62'b11111111101000011111000100000000001111101110100010111010111111;
  assign mem[158] = 62'b11111111101111111000011100101011111100101111010101101100001001;
  assign mem[159] = 62'b11111110110101111101101101000000001010100110101010010000011001;
  assign mem[160] = 62'b11111110101111011001010110111001111001111110000010000011100000;
  assign mem[161] = 62'b11111111101111111100001001010101100101100011100111000110101101;
  assign mem[162] = 62'b11111111100111111110001110110011100011010101110001011101110001;
  assign mem[163] = 62'b11111111100101001100101000001010010010101000110101010110010110;
  assign mem[164] = 62'b11111111011100000100100100100111011000000000010001111011100111;
  assign mem[165] = 62'b11111111101100110000011111000011110011111111001111110001011100;
  assign mem[166] = 62'b11111111101110010000100110101001001011001010111100000101111110;
  assign mem[167] = 62'b11111111010100110100011110001001000010011110001110011101101010;
  assign mem[168] = 62'b11111111010000010011111011100000001110001101111111110110101110;
  assign mem[169] = 62'b11111111101110111100010111100010100011111001000111001111000010;
  assign mem[170] = 62'b11111111101011101001011010101001100111001101011001000011010010;
  assign mem[171] = 62'b11111111100000000111001111110010000111010011000011111010110111;
  assign mem[172] = 62'b11111111100011011000000101100010110001000001100101100111110011;
  assign mem[173] = 62'b11111111101001011101110111111011110100110001111101011101000010;
  assign mem[174] = 62'b11111111101111101101010111100101110001100101011101011101000001;
  assign mem[175] = 62'b11111111000001001110011111000011001110110110101111010101110111;
  assign mem[176] = 62'b11111111000100010101010111011010110001001010010011111001011010;
  assign mem[177] = 62'b11111111101111100101111111100100100100110010010000100110011011;
  assign mem[178] = 62'b11111111101001111011110100001111101111001010011010111110010100;
  assign mem[179] = 62'b11111111100010101111101101101100100101111110101111001111101010;
  assign mem[180] = 62'b11111111100000110010010111000001001101010111011000100110001111;
  assign mem[181] = 62'b11111111101011001111100100110100111110111101010101011100010010;
  assign mem[182] = 62'b11111111101111001000100101001011110111011101100011101011011010;
  assign mem[183] = 62'b11111111001101100100110100111111100101010001010100001100010001;
  assign mem[184] = 62'b11111111010110010011000111110111011101001111110010011111000110;
  assign mem[185] = 62'b11111111101101111111101010111001100010001011011011111000101011;
  assign mem[186] = 62'b11111111101101000101111110011101110100001111100011010111011100;
  assign mem[187] = 62'b11111111011010101001101100100000101011011011010011111111001010;
  assign mem[188] = 62'b11111111100101110001110111101110111110011001010000000110001100;
  assign mem[189] = 62'b11111111100111011100011110011101011111000000110111001001100001;
  assign mem[190] = 62'b11111111101111111110100111001011101111111111101111011101011101;
  assign mem[191] = 62'b11111110100010110110000110010101110101100101000101010111001101;
  assign mem[192] = 62'b11111110100010110110000110010101110101100101000101010111001101;
  assign mem[193] = 62'b11111111101111111110100111001011101111111111101111011101011101;
  assign mem[194] = 62'b11111111100111011100011110011101011111000000110111001001100001;
  assign mem[195] = 62'b11111111100101110001110111101110111110011001010000000110001100;
  assign mem[196] = 62'b11111111011010101001101100100000101011011011010011111111001010;
  assign mem[197] = 62'b11111111101101000101111110011101110100001111100011010111011100;
  assign mem[198] = 62'b11111111101101111111101010111001100010001011011011111000101011;
  assign mem[199] = 62'b11111111010110010011000111110111011101001111110010011111000110;
  assign mem[200] = 62'b11111111001101100100110100111111100101010001010100001100010001;
  assign mem[201] = 62'b11111111101111001000100101001011110111011101100011101011011010;
  assign mem[202] = 62'b11111111101011001111100100110100111110111101010101011100010010;
  assign mem[203] = 62'b11111111100000110010010111000001001101010111011000100110001111;
  assign mem[204] = 62'b11111111100010101111101101101100100101111110101111001111101010;
  assign mem[205] = 62'b11111111101001111011110100001111101111001010011010111110010100;
  assign mem[206] = 62'b11111111101111100101111111100100100100110010010000100110011011;
  assign mem[207] = 62'b11111111000100010101010111011010110001001010010011111001011010;
  assign mem[208] = 62'b11111111000001001110011111000011001110110110101111010101110111;
  assign mem[209] = 62'b11111111101111101101010111100101110001100101011101011101000001;
  assign mem[210] = 62'b11111111101001011101110111111011110100110001111101011101000010;
  assign mem[211] = 62'b11111111100011011000000101100010110001000001100101100111110011;
  assign mem[212] = 62'b11111111100000000111001111110010000111010011000011111010110111;
  assign mem[213] = 62'b11111111101011101001011010101001100111001101011001000011010010;
  assign mem[214] = 62'b11111111101110111100010111100010100011111001000111001111000010;
  assign mem[215] = 62'b11111111010000010011111011100000001110001101111111110110101110;
  assign mem[216] = 62'b11111111010100110100011110001001000010011110001110011101101010;
  assign mem[217] = 62'b11111111101110010000100110101001001011001010111100000101111110;
  assign mem[218] = 62'b11111111101100110000011111000011110011111111001111110001011100;
  assign mem[219] = 62'b11111111011100000100100100100111011000000000010001111011100111;
  assign mem[220] = 62'b11111111100101001100101000001010010010101000110101010110010110;
  assign mem[221] = 62'b11111111100111111110001110110011100011010101110001011101110001;
  assign mem[222] = 62'b11111111101111111100001001010101100101100011100111000110101101;
  assign mem[223] = 62'b11111110101111011001010110111001111001111110000010000011100000;
  assign mem[224] = 62'b11111110110101111101101101000000001010100110101010010000011001;
  assign mem[225] = 62'b11111111101111111000011100101011111100101111010101101100001001;
  assign mem[226] = 62'b11111111101000011111000100000000001111101110100010111010111111;
  assign mem[227] = 62'b11111111100100100110100100010010011011100110110000100100111001;
  assign mem[228] = 62'b11111111011101011110010111011101011011100001101110001110001001;
  assign mem[229] = 62'b11111111101100011001111000101100110100100010000111001110011011;
  assign mem[230] = 62'b11111111101110100000010111101110101011010011001101000100001101;
  assign mem[231] = 62'b11111111010011010101000001000011000010111000011000000101010010;
  assign mem[232] = 62'b11111111010001110100110100010000111111010011001101101100111110;
  assign mem[233] = 62'b11111111101110101110111101100011001000110111110000101101110100;
  assign mem[234] = 62'b11111111101100000010001100010000100110011100100101010101001001;
  assign mem[235] = 62'b11111111011110110111000001100101010010111011110111100011010110;
  assign mem[236] = 62'b11111111100011111111101101100101010011010001010101011011010100;
  assign mem[237] = 62'b11111111101000111110111100110010100011111011111001010000001101;
  assign mem[238] = 62'b11111111101111110011100001010111111101011011011010011001111011;
  assign mem[239] = 62'b11111110111100001101111000010111000111100111101100001011010101;
  assign mem[240] = 62'b11111111000111011011011101100111011110010100001011111100110001;
  assign mem[241] = 62'b11111111101111011101011001100110100011101000010010000001110111;
  assign mem[242] = 62'b11111111101010011000110000100100011011000000101111101011100010;
  assign mem[243] = 62'b11111111100010000110100111100110011001001100111110101101011001;
  assign mem[244] = 62'b11111111100001011100110100110101100011110111101101101101001001;
  assign mem[245] = 62'b11111111101010110100101011110010011110001000011101010100010001;
  assign mem[246] = 62'b11111111101111010011100110000000111011000010110010111100101101;
  assign mem[247] = 62'b11111111001010100000101010000000100101101100000000010001010001;
  assign mem[248] = 62'b11111111010111110000111010100100110001000111011100110011100111;
  assign mem[249] = 62'b11111111101101101101100101001001100010001110001010000010011011;
  assign mem[250] = 62'b11111111101101011010010110000101110011110010011110011010001011;
  assign mem[251] = 62'b11111111011001001101110010101001100011101111001001001111010111;
  assign mem[252] = 62'b11111111100110010110010001100100100101111100000111100000111101;
  assign mem[253] = 62'b11111111100110111001110100010001010100111010101010100010101111;
  assign mem[254] = 62'b11111111101111111111110110001000010110100110111001001011011011;
  assign mem[255] = 62'b11111110001001001000011101000111111100110111101100011110000100;
  assign mem[256] = 62'b11111101111001001000011111000011111110011001110000000001110001;
  assign mem[257] = 62'b11111111101111111111111101100010000101100011101000101010010010;
  assign mem[258] = 62'b11111111100110110001000000110101110011110000011000001001110101;
  assign mem[259] = 62'b11111111100110011111001111011110000100100100011010111100010000;
  assign mem[260] = 62'b11111111011000110110101010010100101110110010001010010010110000;
  assign mem[261] = 62'b11111111101101011111010000101100000010101110001110110011111001;
  assign mem[262] = 62'b11111111101101101000111000001110101001011001101000100110001000;
  assign mem[263] = 62'b11111111011000001000001110001110110000010011101010101011000100;
  assign mem[264] = 62'b11111111001001101111011100101111110010110111000100001101100110;
  assign mem[265] = 62'b11111111101111010110001010001010110001011110001001111010000100;
  assign mem[266] = 62'b11111111101010101101110011001001011001000101101100000011010100;
  assign mem[267] = 62'b11111111100001100111010101101000001001111100101011100110111000;
  assign mem[268] = 62'b11111111100001111100001111000010001011101111001000011000011011;
  assign mem[269] = 62'b11111111101010011111110101100001010010100111111110011010011101;
  assign mem[270] = 62'b11111111101111011011000011111101111101111101011011101110110111;
  assign mem[271] = 62'b11111111001000001100110110011011101000100111000110010011000110;
  assign mem[272] = 62'b11111110111010101001111011011100100100010010010101110000000011;
  assign mem[273] = 62'b11111111101111110100110111100100010100001000100000101110000100;
  assign mem[274] = 62'b11111111101000110111000100010100110011000101101001100011001100;
  assign mem[275] = 62'b11111111100100001001011111111100010111100011100110101110110001;
  assign mem[276] = 62'b11111111011110100000111110000011101010111110000101000100010100;
  assign mem[277] = 62'b11111111101100001000001101111000111111101010010111000110110000;
  assign mem[278] = 62'b11111111101110101011011011001011101000111001111010100010001110;
  assign mem[279] = 62'b11111111010010001100111011101110101011110000111011101101110001;
  assign mem[280] = 62'b11111111010010111101000010001011011010111011000000001110000111;
  assign mem[281] = 62'b11111111101110100100001000010000110110000111011111011111110010;
  assign mem[282] = 62'b11111111101100010100000100001000000001001010110110100100000111;
  assign mem[283] = 62'b11111111011101110100101000111100010100100000011100110001011000;
  assign mem[284] = 62'b11111111100100011100111011010100011011100110000111001101000111;
  assign mem[285] = 62'b11111111101000100111000111111010011010010011011101010010101010;
  assign mem[286] = 62'b11111111101111110111010101001110011111111100011111010001010110;
  assign mem[287] = 62'b11111110110111100001110101100001101010010111010101101100100001;
  assign mem[288] = 62'b11111110101100010000101000110100010010110000001101011111100011;
  assign mem[289] = 62'b11111111101111111100111000001100001111100011010101011101011100;
  assign mem[290] = 62'b11111111100111110101111000001101101100110000110011110110110010;
  assign mem[291] = 62'b11111111100101010110000001000000111000100101110101000100110111;
  assign mem[292] = 62'b11111111011011101101111100111100100011000001001011110100000001;
  assign mem[293] = 62'b11111111101100110101111101100110001001100010110011001011110110;
  assign mem[294] = 62'b11111111101110001100011110101011101000011100001100111000100101;
  assign mem[295] = 62'b11111111010101001100001101100010000000101011110011110000100100;
  assign mem[296] = 62'b11111111001111110111001101110000011010110111111110110111111001;
  assign mem[297] = 62'b11111111101110111111100010001000001100000010111001010111101100;
  assign mem[298] = 62'b11111111101011100011000011100011010010011101010000010011101001;
  assign mem[299] = 62'b11111111100000010010000101011000100110101011100010001000011010;
  assign mem[300] = 62'b11111111100011001110000100000000001101000011001000111001010111;
  assign mem[301] = 62'b11111111101001100101011100111100101110110110000000110100100010;
  assign mem[302] = 62'b11111111101111101011101000111010001110010001101100111110111011;
  assign mem[303] = 62'b11111111000010000000010001011011010100111011000111101111001111;
  assign mem[304] = 62'b11111111000011100011101101101110110000110011011000110100010100;
  assign mem[305] = 62'b11111111101111100111111100111001010101101011011011001011001000;
  assign mem[306] = 62'b11111111101001110100011011000111110101111010101000000011010101;
  assign mem[307] = 62'b11111111100010111001111000000011100011111010001110101000010111;
  assign mem[308] = 62'b11111111100000100111101001000001110100000101111100010111100001;
  assign mem[309] = 62'b11111111101011010110001000100111111110100100100001010000000101;
  assign mem[310] = 62'b11111111101111000101101000111101010011111101110010000001011101;
  assign mem[311] = 62'b11111111001110010101101100101000011110000100000001101000011011;
  assign mem[312] = 62'b11111111010101111011100010011100110111100111101010011010010011;
  assign mem[313] = 62'b11111111101110000100000000110011001010001010011000000010101100;
  assign mem[314] = 62'b11111111101101000000101101010011111110101100101011110110010010;
  assign mem[315] = 62'b11111111011011000000100000110101101100011111110100000000001001;
  assign mem[316] = 62'b11111111100101101000101000110100101010010111010111001001010000;
  assign mem[317] = 62'b11111111100111100101000000000001010111010011110101010111100101;
  assign mem[318] = 62'b11111111101111111110000111000111011010110110111000000111011111;
  assign mem[319] = 62'b11111110100101111111000000000011010010100100001100110101000011;
  assign mem[320] = 62'b11111110011111011010010011011100110001110100011100111100000001;
  assign mem[321] = 62'b11111111101111111111000010010100011101111100011101001111111000;
  assign mem[322] = 62'b11111111100111010011111001010010001101101010001101001010001101;
  assign mem[323] = 62'b11111111100101111011000011010010010101100000110111000001110100;
  assign mem[324] = 62'b11111111011010010010110100000100100111110111101010000111100101;
  assign mem[325] = 62'b11111111101101001011001011001000100000111000001110111110011111;
  assign mem[326] = 62'b11111111101101111011010000010111110111110111100100011111011010;
  assign mem[327] = 62'b11111111010110101010101001110101111101110001110111111000010111;
  assign mem[328] = 62'b11111111001100110011111000110010110011000100101011001010000110;
  assign mem[329] = 62'b11111111101111001011011100100111001001000010001001101010011101;
  assign mem[330] = 62'b11111111101011001000111100110101000111000000000001001110110100;
  assign mem[331] = 62'b11111111100000111101000010011010111011001010101000111001111110;
  assign mem[332] = 62'b11111111100010100101100000011100100111011000101001110010101000;
  assign mem[333] = 62'b11111111101010000011001001010111101010101110101111100100110111;
  assign mem[334] = 62'b11111111101111100011111101010111111111101011100100000111011011;
  assign mem[335] = 62'b11111111000101000110111101111110000101100101111100010111110010;
  assign mem[336] = 62'b11111111000000011100101010000001000111101110101000001100011101;
  assign mem[337] = 62'b11111111101111101111000001011000010111111001000100000110000110;
  assign mem[338] = 62'b11111111101001010110001110111111100100100011100110110111010111;
  assign mem[339] = 62'b11111111100011100010000100000110000101110111111110101100100010;
  assign mem[340] = 62'b11111111011111111000101111011001001011111001110001001000010000;
  assign mem[341] = 62'b11111111101011101111101101011111000100100100111000000011101010;
  assign mem[342] = 62'b11111111101110111001001000001011100010010110101001110110111100;
  assign mem[343] = 62'b11111111010000101100001101100111001111110110111101101110010000;
  assign mem[344] = 62'b11111111010100011100101011100010100101010101110001000001010100;
  assign mem[345] = 62'b11111111101110010100101001111100000100011100101001111111111100;
  assign mem[346] = 62'b11111111101100101010111100000101101001101000001011100100000000;
  assign mem[347] = 62'b11111111011100011011000111111101001001100101110000000000001011;
  assign mem[348] = 62'b11111111100101000011001100000010011111010110011010000010011011;
  assign mem[349] = 62'b11111111101000000110100001101100110011101101010111101011001100;
  assign mem[350] = 62'b11111111101111111011010101100011101100101101100111001111000100;
  assign mem[351] = 62'b11111110110001010001000000000100110100110101110000100110110011;
  assign mem[352] = 62'b11111110110100011001100001000101111001001001110010000010010110;
  assign mem[353] = 62'b11111111101111111001011111001110101111001011100011100101000000;
  assign mem[354] = 62'b11111111101000010110111100010100011010111010010101100011001100;
  assign mem[355] = 62'b11111111100100110000001010000101000101111011000000000000000100;
  assign mem[356] = 62'b11111111011101001000000001011011101000111010011101101101011011;
  assign mem[357] = 62'b11111111101100011111101000111001010010001000110011110011110011;
  assign mem[358] = 62'b11111111101110011100100010011111011011011010101001011101000100;
  assign mem[359] = 62'b11111111010011101100111100111011111010000001000001010010110111;
  assign mem[360] = 62'b11111111010001011100101010000011010111011101100101000101110111;
  assign mem[361] = 62'b11111111101110110010011011001011010011110000111011111110000100;
  assign mem[362] = 62'b11111111101011111100000110010011100001010100110111011111011101;
  assign mem[363] = 62'b11111111011111001101000000010110010110001111111101000001100111;
  assign mem[364] = 62'b11111111100011110101111000001000111000110001011000001101000100;
  assign mem[365] = 62'b11111111101001000110110001011001101111110101001001110110100010;
  assign mem[366] = 62'b11111111101111110010000110010001101100111111101011011100100001;
  assign mem[367] = 62'b11111110111101110001110000111011001011101011101001111111001001;
  assign mem[368] = 62'b11111111000110101010000001001100000100111101100100101010110010;
  assign mem[369] = 62'b11111111101111011111101010011000101001111001100011110101101110;
  assign mem[370] = 62'b11111111101010010001100111100011001000000100011001101011001000;
  assign mem[371] = 62'b11111111100010010000111101010111111011100110001010110000011111;
  assign mem[372] = 62'b11111111100001010010010001010110101111001100110110110011101011;
  assign mem[373] = 62'b11111111101010111011100000010010110100001111000001010001110100;
  assign mem[374] = 62'b11111111101111010000111101000010000101111111111001001011011101;
  assign mem[375] = 62'b11111111001011010001110011001011101111001111010110011100100010;
  assign mem[376] = 62'b11111111010111011001100011010000001111001001000001100011110110;
  assign mem[377] = 62'b11111111101101110010001101011111001011010000010000001001100000;
  assign mem[378] = 62'b11111111101101010101010110111101010010111010010011111010110001;
  assign mem[379] = 62'b11111111011001100100110111000101100001010000011011110111111111;
  assign mem[380] = 62'b11111111100110001101010000001110100011000111000001101111101001;
  assign mem[381] = 62'b11111111100111000010100100001010110011000101110110110101111010;
  assign mem[382] = 62'b11111111101111111111101001110010110100010010110101000110100001;
  assign mem[383] = 62'b11111110010010110110010011011010111011111000110000111011111101;
  assign mem[384] = 62'b11111110010010110110010011011010111011111000110000111011111101;
  assign mem[385] = 62'b11111111101111111111101001110010110100010010110101000110100001;
  assign mem[386] = 62'b11111111100111000010100100001010110011000101110110110101111010;
  assign mem[387] = 62'b11111111100110001101010000001110100011000111000001101111101001;
  assign mem[388] = 62'b11111111011001100100110111000101100001010000011011110111111111;
  assign mem[389] = 62'b11111111101101010101010110111101010010111010010011111010110001;
  assign mem[390] = 62'b11111111101101110010001101011111001011010000010000001001100000;
  assign mem[391] = 62'b11111111010111011001100011010000001111001001000001100011110110;
  assign mem[392] = 62'b11111111001011010001110011001011101111001111010110011100100010;
  assign mem[393] = 62'b11111111101111010000111101000010000101111111111001001011011101;
  assign mem[394] = 62'b11111111101010111011100000010010110100001111000001010001110100;
  assign mem[395] = 62'b11111111100001010010010001010110101111001100110110110011101011;
  assign mem[396] = 62'b11111111100010010000111101010111111011100110001010110000011111;
  assign mem[397] = 62'b11111111101010010001100111100011001000000100011001101011001000;
  assign mem[398] = 62'b11111111101111011111101010011000101001111001100011110101101110;
  assign mem[399] = 62'b11111111000110101010000001001100000100111101100100101010110010;
  assign mem[400] = 62'b11111110111101110001110000111011001011101011101001111111001001;
  assign mem[401] = 62'b11111111101111110010000110010001101100111111101011011100100001;
  assign mem[402] = 62'b11111111101001000110110001011001101111110101001001110110100010;
  assign mem[403] = 62'b11111111100011110101111000001000111000110001011000001101000100;
  assign mem[404] = 62'b11111111011111001101000000010110010110001111111101000001100111;
  assign mem[405] = 62'b11111111101011111100000110010011100001010100110111011111011101;
  assign mem[406] = 62'b11111111101110110010011011001011010011110000111011111110000100;
  assign mem[407] = 62'b11111111010001011100101010000011010111011101100101000101110111;
  assign mem[408] = 62'b11111111010011101100111100111011111010000001000001010010110111;
  assign mem[409] = 62'b11111111101110011100100010011111011011011010101001011101000100;
  assign mem[410] = 62'b11111111101100011111101000111001010010001000110011110011110011;
  assign mem[411] = 62'b11111111011101001000000001011011101000111010011101101101011011;
  assign mem[412] = 62'b11111111100100110000001010000101000101111011000000000000000100;
  assign mem[413] = 62'b11111111101000010110111100010100011010111010010101100011001100;
  assign mem[414] = 62'b11111111101111111001011111001110101111001011100011100101000000;
  assign mem[415] = 62'b11111110110100011001100001000101111001001001110010000010010110;
  assign mem[416] = 62'b11111110110001010001000000000100110100110101110000100110110011;
  assign mem[417] = 62'b11111111101111111011010101100011101100101101100111001111000100;
  assign mem[418] = 62'b11111111101000000110100001101100110011101101010111101011001100;
  assign mem[419] = 62'b11111111100101000011001100000010011111010110011010000010011011;
  assign mem[420] = 62'b11111111011100011011000111111101001001100101110000000000001011;
  assign mem[421] = 62'b11111111101100101010111100000101101001101000001011100100000000;
  assign mem[422] = 62'b11111111101110010100101001111100000100011100101001111111111100;
  assign mem[423] = 62'b11111111010100011100101011100010100101010101110001000001010100;
  assign mem[424] = 62'b11111111010000101100001101100111001111110110111101101110010000;
  assign mem[425] = 62'b11111111101110111001001000001011100010010110101001110110111100;
  assign mem[426] = 62'b11111111101011101111101101011111000100100100111000000011101010;
  assign mem[427] = 62'b11111111011111111000101111011001001011111001110001001000010000;
  assign mem[428] = 62'b11111111100011100010000100000110000101110111111110101100100010;
  assign mem[429] = 62'b11111111101001010110001110111111100100100011100110110111010111;
  assign mem[430] = 62'b11111111101111101111000001011000010111111001000100000110000110;
  assign mem[431] = 62'b11111111000000011100101010000001000111101110101000001100011101;
  assign mem[432] = 62'b11111111000101000110111101111110000101100101111100010111110010;
  assign mem[433] = 62'b11111111101111100011111101010111111111101011100100000111011011;
  assign mem[434] = 62'b11111111101010000011001001010111101010101110101111100100110111;
  assign mem[435] = 62'b11111111100010100101100000011100100111011000101001110010101000;
  assign mem[436] = 62'b11111111100000111101000010011010111011001010101000111001111110;
  assign mem[437] = 62'b11111111101011001000111100110101000111000000000001001110110100;
  assign mem[438] = 62'b11111111101111001011011100100111001001000010001001101010011101;
  assign mem[439] = 62'b11111111001100110011111000110010110011000100101011001010000110;
  assign mem[440] = 62'b11111111010110101010101001110101111101110001110111111000010111;
  assign mem[441] = 62'b11111111101101111011010000010111110111110111100100011111011010;
  assign mem[442] = 62'b11111111101101001011001011001000100000111000001110111110011111;
  assign mem[443] = 62'b11111111011010010010110100000100100111110111101010000111100101;
  assign mem[444] = 62'b11111111100101111011000011010010010101100000110111000001110100;
  assign mem[445] = 62'b11111111100111010011111001010010001101101010001101001010001101;
  assign mem[446] = 62'b11111111101111111111000010010100011101111100011101001111111000;
  assign mem[447] = 62'b11111110011111011010010011011100110001110100011100111100000001;
  assign mem[448] = 62'b11111110100101111111000000000011010010100100001100110101000011;
  assign mem[449] = 62'b11111111101111111110000111000111011010110110111000000111011111;
  assign mem[450] = 62'b11111111100111100101000000000001010111010011110101010111100101;
  assign mem[451] = 62'b11111111100101101000101000110100101010010111010111001001010000;
  assign mem[452] = 62'b11111111011011000000100000110101101100011111110100000000001001;
  assign mem[453] = 62'b11111111101101000000101101010011111110101100101011110110010010;
  assign mem[454] = 62'b11111111101110000100000000110011001010001010011000000010101100;
  assign mem[455] = 62'b11111111010101111011100010011100110111100111101010011010010011;
  assign mem[456] = 62'b11111111001110010101101100101000011110000100000001101000011011;
  assign mem[457] = 62'b11111111101111000101101000111101010011111101110010000001011101;
  assign mem[458] = 62'b11111111101011010110001000100111111110100100100001010000000101;
  assign mem[459] = 62'b11111111100000100111101001000001110100000101111100010111100001;
  assign mem[460] = 62'b11111111100010111001111000000011100011111010001110101000010111;
  assign mem[461] = 62'b11111111101001110100011011000111110101111010101000000011010101;
  assign mem[462] = 62'b11111111101111100111111100111001010101101011011011001011001000;
  assign mem[463] = 62'b11111111000011100011101101101110110000110011011000110100010100;
  assign mem[464] = 62'b11111111000010000000010001011011010100111011000111101111001111;
  assign mem[465] = 62'b11111111101111101011101000111010001110010001101100111110111011;
  assign mem[466] = 62'b11111111101001100101011100111100101110110110000000110100100010;
  assign mem[467] = 62'b11111111100011001110000100000000001101000011001000111001010111;
  assign mem[468] = 62'b11111111100000010010000101011000100110101011100010001000011010;
  assign mem[469] = 62'b11111111101011100011000011100011010010011101010000010011101001;
  assign mem[470] = 62'b11111111101110111111100010001000001100000010111001010111101100;
  assign mem[471] = 62'b11111111001111110111001101110000011010110111111110110111111001;
  assign mem[472] = 62'b11111111010101001100001101100010000000101011110011110000100100;
  assign mem[473] = 62'b11111111101110001100011110101011101000011100001100111000100101;
  assign mem[474] = 62'b11111111101100110101111101100110001001100010110011001011110110;
  assign mem[475] = 62'b11111111011011101101111100111100100011000001001011110100000001;
  assign mem[476] = 62'b11111111100101010110000001000000111000100101110101000100110111;
  assign mem[477] = 62'b11111111100111110101111000001101101100110000110011110110110010;
  assign mem[478] = 62'b11111111101111111100111000001100001111100011010101011101011100;
  assign mem[479] = 62'b11111110101100010000101000110100010010110000001101011111100011;
  assign mem[480] = 62'b11111110110111100001110101100001101010010111010101101100100001;
  assign mem[481] = 62'b11111111101111110111010101001110011111111100011111010001010110;
  assign mem[482] = 62'b11111111101000100111000111111010011010010011011101010010101010;
  assign mem[483] = 62'b11111111100100011100111011010100011011100110000111001101000111;
  assign mem[484] = 62'b11111111011101110100101000111100010100100000011100110001011000;
  assign mem[485] = 62'b11111111101100010100000100001000000001001010110110100100000111;
  assign mem[486] = 62'b11111111101110100100001000010000110110000111011111011111110010;
  assign mem[487] = 62'b11111111010010111101000010001011011010111011000000001110000111;
  assign mem[488] = 62'b11111111010010001100111011101110101011110000111011101101110001;
  assign mem[489] = 62'b11111111101110101011011011001011101000111001111010100010001110;
  assign mem[490] = 62'b11111111101100001000001101111000111111101010010111000110110000;
  assign mem[491] = 62'b11111111011110100000111110000011101010111110000101000100010100;
  assign mem[492] = 62'b11111111100100001001011111111100010111100011100110101110110001;
  assign mem[493] = 62'b11111111101000110111000100010100110011000101101001100011001100;
  assign mem[494] = 62'b11111111101111110100110111100100010100001000100000101110000100;
  assign mem[495] = 62'b11111110111010101001111011011100100100010010010101110000000011;
  assign mem[496] = 62'b11111111001000001100110110011011101000100111000110010011000110;
  assign mem[497] = 62'b11111111101111011011000011111101111101111101011011101110110111;
  assign mem[498] = 62'b11111111101010011111110101100001010010100111111110011010011101;
  assign mem[499] = 62'b11111111100001111100001111000010001011101111001000011000011011;
  assign mem[500] = 62'b11111111100001100111010101101000001001111100101011100110111000;
  assign mem[501] = 62'b11111111101010101101110011001001011001000101101100000011010100;
  assign mem[502] = 62'b11111111101111010110001010001010110001011110001001111010000100;
  assign mem[503] = 62'b11111111001001101111011100101111110010110111000100001101100110;
  assign mem[504] = 62'b11111111011000001000001110001110110000010011101010101011000100;
  assign mem[505] = 62'b11111111101101101000111000001110101001011001101000100110001000;
  assign mem[506] = 62'b11111111101101011111010000101100000010101110001110110011111001;
  assign mem[507] = 62'b11111111011000110110101010010100101110110010001010010010110000;
  assign mem[508] = 62'b11111111100110011111001111011110000100100100011010111100010000;
  assign mem[509] = 62'b11111111100110110001000000110101110011110000011000001001110101;
  assign mem[510] = 62'b11111111101111111111111101100010000101100011101000101010010010;
  assign mem[511] = 62'b11111101111001001000011111000011111110011001110000000001110001;
  assign mem[512] = 62'b11111101101001001000011111100010111110110011001010010010111010;
  assign mem[513] = 62'b11111111101111111111111111011000100001011000100001110100000010;
  assign mem[514] = 62'b11111111100110101100100101110011101101001011111110001010011100;
  assign mem[515] = 62'b11111111100110100011101101000111101010101000011001110001110001;
  assign mem[516] = 62'b11111111011000101011000100101110000110110101011110110101000100;
  assign mem[517] = 62'b11111111101101100001101100010010000100010001011010010001001111;
  assign mem[518] = 62'b11111111101101100110100000000011011101100010110011110101000110;
  assign mem[519] = 62'b11111111011000010011110110101010101010111100111001000000111111;
  assign mem[520] = 62'b11111111001001010110110100100111101001101101100010101011111010;
  assign mem[521] = 62'b11111111101111010111011010011011101101010000110110100001011101;
  assign mem[522] = 62'b11111111101010101010010101010001111010001011001011100110001110;
  assign mem[523] = 62'b11111111100001101100100101000000010111000100110111001110111111;
  assign mem[524] = 62'b11111111100001110111000001101101100100110111000100100001110010;
  assign mem[525] = 62'b11111111101010100011010110011101101110010101000101101011010010;
  assign mem[526] = 62'b11111111101111011001110111010101010110100010000011110011101110;
  assign mem[527] = 62'b11111111001000100101100001011100100111110001000001100000000100;
  assign mem[528] = 62'b11111110111001110111111011011011101011001001001010100001011100;
  assign mem[529] = 62'b11111111101111110101100000110100101101101001110101110010011110;
  assign mem[530] = 62'b11111111101000110011000110101001110101000110000100011001010101;
  assign mem[531] = 62'b11111111100100001110010111111101011011001010100100001110000000;
  assign mem[532] = 62'b11111111011110010101111010100001101101001111001101100000100101;
  assign mem[533] = 62'b11111111101100001011001101000101001001001100011110001111110001;
  assign mem[534] = 62'b11111111101110101001101000001110010011111001100101100000000000;
  assign mem[535] = 62'b11111111010010011000111110011010011001010101010101010010111010;
  assign mem[536] = 62'b11111111010010110001000001101001001110100101010100010100100000;
  assign mem[537] = 62'b11111111101110100101111110110000110110000000010110101100110000;
  assign mem[538] = 62'b11111111101100010001001000001100110001010000011100000000000100;
  assign mem[539] = 62'b11111111011101111111101111111101100110101010010100000111011110;
  assign mem[540] = 62'b11111111100100011000000101101001101001001010110011001010100010;
  assign mem[541] = 62'b11111111101000101011001000011100011110110111100001110110001000;
  assign mem[542] = 62'b11111111101111110110101111101001110101000101000101001110001100;
  assign mem[543] = 62'b11111110111000010011111000011100010010110000010011000010100001;
  assign mem[544] = 62'b11111110101010101100010000000110111101010111111000001100010111;
  assign mem[545] = 62'b11111111101111111101001101110001010100101100011011111011010011;
  assign mem[546] = 62'b11111111100111110001101011100010011100111000101101001100110011;
  assign mem[547] = 62'b11111111100101011010101100001101010001100101110110010010011111;
  assign mem[548] = 62'b11111111011011100010100111100000010100111111010101011010010011;
  assign mem[549] = 62'b11111111101100111000101011001100100111100110011010000001100000;
  assign mem[550] = 62'b11111111101110001010011000111101000100001110010001100101111010;
  assign mem[551] = 62'b11111111010101011000000100000000010010111101000110011110110100;
  assign mem[552] = 62'b11111111001111011110110111010010000000101111010011100000000010;
  assign mem[553] = 62'b11111111101111000001000101101000010100110011110111001110001100;
  assign mem[554] = 62'b11111111101011011111110110011010000110111001111001001011101001;
  assign mem[555] = 62'b11111111100000010111011111001111101100001100011011100010110111;
  assign mem[556] = 62'b11111111100011001001000010000111101100010010011010011000011111;
  assign mem[557] = 62'b11111111101001101001001101111110100100001010110000011010110010;
  assign mem[558] = 62'b11111111101111101010101111101111001011000011001111110111011100;
  assign mem[559] = 62'b11111111000010011001001001100101001101111111010011010000001001;
  assign mem[560] = 62'b11111111000011001010110111101111111001010001010001011010100111;
  assign mem[561] = 62'b11111111101111101000111001101110101100011110100001011110010001;
  assign mem[562] = 62'b11111111101001110000101101000100010000111100000111010111000010;
  assign mem[563] = 62'b11111111100010111110111100001001001011010001000001000000010101;
  assign mem[564] = 62'b11111111100000100010010001000100100000001100101011000010001100;
  assign mem[565] = 62'b11111111101011011001011000111100010100111111011011110001000111;
  assign mem[566] = 62'b11111111101111000100001001000010111100100010011000111101011111;
  assign mem[567] = 62'b11111111001110101110000110101101000110001011011110001101001000;
  assign mem[568] = 62'b11111111010101101111101110011110001011100111011011001110110110;
  assign mem[569] = 62'b11111111101110000110001010000000101111110111000110011011011001;
  assign mem[570] = 62'b11111111101100111110000011000011101000110011100100011001111011;
  assign mem[571] = 62'b11111111011011001011111001011100011101101100110001100101110010;
  assign mem[572] = 62'b11111111100101100100000000000111010101111101110010001111011111;
  assign mem[573] = 62'b11111111100111101001001111011100000111101111111001011111010010;
  assign mem[574] = 62'b11111111101111111101110101001110111011000110111001000101100100;
  assign mem[575] = 62'b11111110100111100011011011101010100101100001110100011010000110;
  assign mem[576] = 62'b11111110011100010001010100111101001100111001010011101100011101;
  assign mem[577] = 62'b11111111101111111111001110000010011100111000101010011001111001;
  assign mem[578] = 62'b11111111100111001111100101010110001110000001111001100101000010;
  assign mem[579] = 62'b11111111100101111111100111110010111101111001010110101000010000;
  assign mem[580] = 62'b11111111011010000111010110010101000011101101010000101011000000;
  assign mem[581] = 62'b11111111101101001101101111110001111011110010111111101111011100;
  assign mem[582] = 62'b11111111101101111001000001011000001111011011011000110110000001;
  assign mem[583] = 62'b11111111010110110110011001100001100011100010100000110010110110;
  assign mem[584] = 62'b11111111001100011011011001000001010011010111010111010011011101;
  assign mem[585] = 62'b11111111101111001100110110100001011010001110101010111011110000;
  assign mem[586] = 62'b11111111101011000101100111010000101010010011001010001011110101;
  assign mem[587] = 62'b11111111100001000010010111001001001000110100001010100101010111;
  assign mem[588] = 62'b11111111100010100000011000101111101111010011010011110010111010;
  assign mem[589] = 62'b11111111101010000110110010011011010010110000001010011101011110;
  assign mem[590] = 62'b11111111101111100010111010011100110111110010110100101101111000;
  assign mem[591] = 62'b11111111000101011111110000000010000110010101001100101111011110;
  assign mem[592] = 62'b11111111000000000011101110100010101101011011111011100001011011;
  assign mem[593] = 62'b11111111101111101111110100011100001111000010101000110110001000;
  assign mem[594] = 62'b11111111101001010010011001000011100011101011000100101001101100;
  assign mem[595] = 62'b11111111100011100111000010001111100011110101100011000000101001;
  assign mem[596] = 62'b11111111011111101101110101011101011100001001001101001011011110;
  assign mem[597] = 62'b11111111101011110010110101010011001011000011010010001100100111;
  assign mem[598] = 62'b11111111101110110111011110101101101010000001111000011001010001;
  assign mem[599] = 62'b11111111010000111000010101101101001110000101110100100111001110;
  assign mem[600] = 62'b11111111010100010000110001000011011100100010010011011011110000;
  assign mem[601] = 62'b11111111101110010110101001110101010101000001000110011111010011;
  assign mem[602] = 62'b11111111101100101000001000111100011001101110011100010001001001;
  assign mem[603] = 62'b11111111011100100110010111111111000011100001100101001110001001;
  assign mem[604] = 62'b11111111100100111110011100110000100101110011001010010010000110;
  assign mem[605] = 62'b11111111101000001010101001110000010011111101010100010111111111;
  assign mem[606] = 62'b11111111101111111010111001110100100101001100000100000100001111;
  assign mem[607] = 62'b11111110110010000011001001011001110100111011010100010001001101;
  assign mem[608] = 62'b11111110110011100111011001111100010010110001011010001010011001;
  assign mem[609] = 62'b11111111101111111001111110101010000101010010000010110101100000;
  assign mem[610] = 62'b11111111101000010010110111000100010001101011111000001111111010;
  assign mem[611] = 62'b11111111100100110100111011110001101101010110001001111101111111;
  assign mem[612] = 62'b11111111011100111100110100101110101110111000011100110100100001;
  assign mem[613] = 62'b11111111101100100010011111010110000111000000101001110000010011;
  assign mem[614] = 62'b11111111101110011010100110000111000101010111010101001110100111;
  assign mem[615] = 62'b11111111010011111000111001101111101001011011101100001001110001;
  assign mem[616] = 62'b11111111010001010000100011111011101111110001101001001101111000;
  assign mem[617] = 62'b11111111101110110100001000001101011110100110011001000000001001;
  assign mem[618] = 62'b11111111101011111001000001101101100001000100010101010011000001;
  assign mem[619] = 62'b11111111011111010111111101111011100110010101101100110110100011;
  assign mem[620] = 62'b11111111100011110000111100010001001001100000011100010100011000;
  assign mem[621] = 62'b11111111101001001010101010010000011111110001011010100000010101;
  assign mem[622] = 62'b11111111101111110001010110111000111011011111011001101011110110;
  assign mem[623] = 62'b11111110111110100011101011011111111101111001001010101000111111;
  assign mem[624] = 62'b11111111000110010001010001101010000011000111011000001100001101;
  assign mem[625] = 62'b11111111101111100000110000111101001010010000001100011000001100;
  assign mem[626] = 62'b11111111101010001110000001100001001010010110010011101111000110;
  assign mem[627] = 62'b11111111100010010110000111001101001100101110110111000100010000;
  assign mem[628] = 62'b11111111100001001100111110100111001111111011100010010101001111;
  assign mem[629] = 62'b11111111101010111110111000111111011000100111110101011110110110;
  assign mem[630] = 62'b11111111101111001111100110101110111100000110111011110001100101;
  assign mem[631] = 62'b11111111001011101010010110001100110100111100010101110110101101;
  assign mem[632] = 62'b11111111010111001101110110001111001001001001100001000010010010;
  assign mem[633] = 62'b11111111101101110100011111111011110011100010101001000101011010;
  assign mem[634] = 62'b11111111101101010010110101101100011011000110000111010100100100;
  assign mem[635] = 62'b11111111011001110000010111110101000100000011011111100111110010;
  assign mem[636] = 62'b11111111100110001000101110010001001111111011000010001011111111;
  assign mem[637] = 62'b11111111100111000110111010110010010110000011100100000110111111;
  assign mem[638] = 62'b11111111101111111111100001110001101000011100001100101101110111;
  assign mem[639] = 62'b11111110010101111111010100110100100001111110101011001000100110;
  assign mem[640] = 62'b11111110001111011010100010100101101010101110011001011111001011;
  assign mem[641] = 62'b11111111101111111111110000100101000011110001010011101111010001;
  assign mem[642] = 62'b11111111100110111110001100101010011001110010010101101101110101;
  assign mem[643] = 62'b11111111100110010001110001010101000011011111110101001101011011;
  assign mem[644] = 62'b11111111011001011001010101010110110111101010111001010010001111;
  assign mem[645] = 62'b11111111101101010111110111000101110010100010001000101001111111;
  assign mem[646] = 62'b11111111101101101111111001111001000011100101010111010110011010;
  assign mem[647] = 62'b11111111010111100101001111010111100110000100111101111110101110;
  assign mem[648] = 62'b11111111001010111001001111000111010101111100111011100110101011;
  assign mem[649] = 62'b11111111101111010010010010001000000110101111001010101110110100;
  assign mem[650] = 62'b11111111101010111000000110100011110011010001011110110011101111;
  assign mem[651] = 62'b11111111100001010111100011011011100100110110111110001010111100;
  assign mem[652] = 62'b11111111100010001011110010110101100110001011000001001111100010;
  assign mem[653] = 62'b11111111101010010101001100100100010000100100001111010100100011;
  assign mem[654] = 62'b11111111101111011110100010100110011100000110100011001000101010;
  assign mem[655] = 62'b11111111000111000010101111110110001101000010001100010011111111;
  assign mem[656] = 62'b11111110111100111111110101001100111011001100000111110111000001;
  assign mem[657] = 62'b11111111101111110010110100011100000011100100010100001101010100;
  assign mem[658] = 62'b11111111101001000010110111100101000011010101110101111011111110;
  assign mem[659] = 62'b11111111100011111010110011001111101010101111100000011010000000;
  assign mem[660] = 62'b11111111011111000010000001100100000110101111111111011111111110;
  assign mem[661] = 62'b11111111101011111111001001110100100101101000011011000101000111;
  assign mem[662] = 62'b11111111101110110000101100111101001011000110101111011010110010;
  assign mem[663] = 62'b11111111010001101000101111011111111011111010001111001001000011;
  assign mem[664] = 62'b11111111010011100000111111010111100011010100111011011010101011;
  assign mem[665] = 62'b11111111101110011110011101101100101001101001010001011001011010;
  assign mem[666] = 62'b11111111101100011100110001010110001001100111101010101011010111;
  assign mem[667] = 62'b11111111011101010011001101000000101011101010000110000010011101;
  assign mem[668] = 62'b11111111100100101011010111100101010001011001110010001011110001;
  assign mem[669] = 62'b11111111101000011011000000101000011101100110101010000110010101;
  assign mem[670] = 62'b11111111101111111000111110100100101011111010011101100010000110;
  assign mem[671] = 62'b11111110110101001011100111011101001010010011010100110100001010;
  assign mem[672] = 62'b11111110110000011110110110000101001110010001100011000001100100;
  assign mem[673] = 62'b11111111101111111011110000000100000010100000100110000110010001;
  assign mem[674] = 62'b11111111101000000010011000101101110101011011100101001011111010;
  assign mem[675] = 62'b11111111100101000111111010100000011100110110011001101010100110;
  assign mem[676] = 62'b11111111011100001111110110110101000111001001100011000100101001;
  assign mem[677] = 62'b11111111101100101101101110001000001010000000001101101010011001;
  assign mem[678] = 62'b11111111101110010010101000110111111111100000011100111001011110;
  assign mem[679] = 62'b11111111010100101000100101001111010001000110111000001011110011;
  assign mem[680] = 62'b11111111010000100000000100111000000101111010110110011000011110;
  assign mem[681] = 62'b11111111101110111010110000011101001100010100001010010101000100;
  assign mem[682] = 62'b11111111101011101100100100100110100000101101101100010000001101;
  assign mem[683] = 62'b11111111100000000001110100000011001000001010111000001011100001;
  assign mem[684] = 62'b11111111100011011101000101001100011011100000010111111110001101;
  assign mem[685] = 62'b11111111101001011010000011111101000010101111010111111111100001;
  assign mem[686] = 62'b11111111101111101110001101000110001101011001101010110110110111;
  assign mem[687] = 62'b11111111000000110101100100110110111100101100100110011110000110;
  assign mem[688] = 62'b11111111000100101110001011000101111111011110011111101010001000;
  assign mem[689] = 62'b11111111101111100100111111000101001111100001011010110000001000;
  assign mem[690] = 62'b11111111101001111111011111010011110001001100010100100111011110;
  assign mem[691] = 62'b11111111100010101010100111011011101000011110101110101101011000;
  assign mem[692] = 62'b11111111100000110111101101000010111000010010111100010010110110;
  assign mem[693] = 62'b11111111101011001100010001010110100101111100110111101111110011;
  assign mem[694] = 62'b11111111101111001010000001011111111100010001100000100111001110;
  assign mem[695] = 62'b11111111001101001100010111011101001101001011001011110111101110;
  assign mem[696] = 62'b11111111010110011110111001010010011100101011010110001111001011;
  assign mem[697] = 62'b11111111101101111101011110001101101010100110111010010110011100;
  assign mem[698] = 62'b11111111101101001000100101010111000110111001011010010011100001;
  assign mem[699] = 62'b11111111011010011110010000110011010011110110111111001100011011;
  assign mem[700] = 62'b11111111100101110110011101111011100111001111100011010001011100;
  assign mem[701] = 62'b11111111100111011000001100010100101100001100000100011101100100;
  assign mem[702] = 62'b11111111101111111110110101010111100100001001011111110110101110;
  assign mem[703] = 62'b11111110100001010001101000010111011011010000101100000101111111;
  assign mem[704] = 62'b11111110100100011010100011100101101111111110000110000101111001;
  assign mem[705] = 62'b11111111101111111110010111110001000010000010001100000000010100;
  assign mem[706] = 62'b11111111100111100000101111101100011011100100001011001101011011;
  assign mem[707] = 62'b11111111100101101101010000101100100110010011110111010001001000;
  assign mem[708] = 62'b11111111011010110101000111001100010010010111001101110000001001;
  assign mem[709] = 62'b11111111101101000011010110011100101111010110011101001010111001;
  assign mem[710] = 62'b11111111101110000001110110011011011001001010000000111101010100;
  assign mem[711] = 62'b11111111010110000111010101100101011100100010001100001000000010;
  assign mem[712] = 62'b11111111001101111101010001011000111111000000010000100110011010;
  assign mem[713] = 62'b11111111101111000111000111101010111110001010000100011100001000;
  assign mem[714] = 62'b11111111101011010010110111010000001001110111100111100100100101;
  assign mem[715] = 62'b11111111100000101101000000010110000111100011111000010111101100;
  assign mem[716] = 62'b11111111100010110100110011001111010011010011101001101110111000;
  assign mem[717] = 62'b11111111101001111000001000001011101101101101000010010001110010;
  assign mem[718] = 62'b11111111101111100110111110110101111100111110111101111000101001;
  assign mem[719] = 62'b11111111000011111100100010111101010111110110110100100010010011;
  assign mem[720] = 62'b11111111000001100111011000100101000000101111100010010011100111;
  assign mem[721] = 62'b11111111101111101100100000110111000110100000011101010101001101;
  assign mem[722] = 62'b11111111101001100001101010111011110001010001010111010110010100;
  assign mem[723] = 62'b11111111100011010011000101001001010010110000010100110111100001;
  assign mem[724] = 62'b11111111100000001100101010111001010101111011011011110110010110;
  assign mem[725] = 62'b11111111101011100110001111101000011111110110010001010101011110;
  assign mem[726] = 62'b11111111101110111101111101011011100101000111001010001111000000;
  assign mem[727] = 62'b11111111010000000111110001100000000110101110011111110111010010;
  assign mem[728] = 62'b11111111010101000000010110001111011100000110010111000001001000;
  assign mem[729] = 62'b11111111101110001110100011001111101100011101011100111010000101;
  assign mem[730] = 62'b11111111101100110011001110111000100000110000101101111010100000;
  assign mem[731] = 62'b11111111011011111001010001010100010111111111111100000011011001;
  assign mem[732] = 62'b11111111100101010001010100111111110101000101011001110111111100;
  assign mem[733] = 62'b11111111100111111010000011111110000111101100000011011010000110;
  assign mem[734] = 62'b11111111101111111100100001011000010100111000010011000111101101;
  assign mem[735] = 62'b11111110101101110101000000011011111001100000001000111011001001;
  assign mem[736] = 62'b11111110110110101111110001101100111110011110011011000100101001;
  assign mem[737] = 62'b11111111101111110111111001100100100010111101110011001100000111;
  assign mem[738] = 62'b11111111101000100011000110011011100111010010000001101110100001;
  assign mem[739] = 62'b11111111100100100001110000001100110000011000001001000111111111;
  assign mem[740] = 62'b11111111011101101001100000110001011100111110100001000011011001;
  assign mem[741] = 62'b11111111101100010110111110111101011001111111101111100001011010;
  assign mem[742] = 62'b11111111101110100010010000100101011011101011010110000000100101;
  assign mem[743] = 62'b11111111010011001001000001111110110110001110001011101010101111;
  assign mem[744] = 62'b11111111010010000000111000010110000011110101110010011110111110;
  assign mem[745] = 62'b11111111101110101101001100111101010001010110111000100000010001;
  assign mem[746] = 62'b11111111101100000101001101100111011100010001100101111001010111;
  assign mem[747] = 62'b11111111011110101100000000011010010101111100100101011000100000;
  assign mem[748] = 62'b11111111100100000100100111001001100110001111010001000010001100;
  assign mem[749] = 62'b11111111101000111011000001000010011011010010000110110001001001;
  assign mem[750] = 62'b11111111101111110100001101000101011000110110000110000010000111;
  assign mem[751] = 62'b11111110111011011011111010011011101100001110001111011001001100;
  assign mem[752] = 62'b11111111000111110100001010011110111011110100101100101100011100;
  assign mem[753] = 62'b11111111101111011100001111011001000011010010110111111010110111;
  assign mem[754] = 62'b11111111101010011100010011100011011110100111010110000011110101;
  assign mem[755] = 62'b11111111100010000001011011101010100001011101010110000011010110;
  assign mem[756] = 62'b11111111100001100010000101100100011111001110100100011011100101;
  assign mem[757] = 62'b11111111101010110001001111111110111101001111101111101011001000;
  assign mem[758] = 62'b11111111101111010100111000101100011111101011110010110100000111;
  assign mem[759] = 62'b11111111001010001000000011111000011011000110000011000111011010;
  assign mem[760] = 62'b11111111010111111100100100110111010011011100110100000111100100;
  assign mem[761] = 62'b11111111101101101011001111010000101100111001101000101010111001;
  assign mem[762] = 62'b11111111101101011100110011111101010000100011000000110111111111;
  assign mem[763] = 62'b11111111011001000010001110111110000001111011110111101111010001;
  assign mem[764] = 62'b11111111100110011010110000111100111111010100101011001110000110;
  assign mem[765] = 62'b11111111100110110101011010111111101111010010101010111111001101;
  assign mem[766] = 62'b11111111101111111111111010011100101100100101111000110001001111;
  assign mem[767] = 62'b11111110000010110110010110101100001110010100001001011100000011;
  assign mem[768] = 62'b11111110000010110110010110101100001110010100001001011100000011;
  assign mem[769] = 62'b11111111101111111111111010011100101100100101111000110001001111;
  assign mem[770] = 62'b11111111100110110101011010111111101111010010101010111111001101;
  assign mem[771] = 62'b11111111100110011010110000111100111111010100101011001110000110;
  assign mem[772] = 62'b11111111011001000010001110111110000001111011110111101111010001;
  assign mem[773] = 62'b11111111101101011100110011111101010000100011000000110111111111;
  assign mem[774] = 62'b11111111101101101011001111010000101100111001101000101010111001;
  assign mem[775] = 62'b11111111010111111100100100110111010011011100110100000111100100;
  assign mem[776] = 62'b11111111001010001000000011111000011011000110000011000111011010;
  assign mem[777] = 62'b11111111101111010100111000101100011111101011110010110100000111;
  assign mem[778] = 62'b11111111101010110001001111111110111101001111101111101011001000;
  assign mem[779] = 62'b11111111100001100010000101100100011111001110100100011011100101;
  assign mem[780] = 62'b11111111100010000001011011101010100001011101010110000011010110;
  assign mem[781] = 62'b11111111101010011100010011100011011110100111010110000011110101;
  assign mem[782] = 62'b11111111101111011100001111011001000011010010110111111010110111;
  assign mem[783] = 62'b11111111000111110100001010011110111011110100101100101100011100;
  assign mem[784] = 62'b11111110111011011011111010011011101100001110001111011001001100;
  assign mem[785] = 62'b11111111101111110100001101000101011000110110000110000010000111;
  assign mem[786] = 62'b11111111101000111011000001000010011011010010000110110001001001;
  assign mem[787] = 62'b11111111100100000100100111001001100110001111010001000010001100;
  assign mem[788] = 62'b11111111011110101100000000011010010101111100100101011000100000;
  assign mem[789] = 62'b11111111101100000101001101100111011100010001100101111001010111;
  assign mem[790] = 62'b11111111101110101101001100111101010001010110111000100000010001;
  assign mem[791] = 62'b11111111010010000000111000010110000011110101110010011110111110;
  assign mem[792] = 62'b11111111010011001001000001111110110110001110001011101010101111;
  assign mem[793] = 62'b11111111101110100010010000100101011011101011010110000000100101;
  assign mem[794] = 62'b11111111101100010110111110111101011001111111101111100001011010;
  assign mem[795] = 62'b11111111011101101001100000110001011100111110100001000011011001;
  assign mem[796] = 62'b11111111100100100001110000001100110000011000001001000111111111;
  assign mem[797] = 62'b11111111101000100011000110011011100111010010000001101110100001;
  assign mem[798] = 62'b11111111101111110111111001100100100010111101110011001100000111;
  assign mem[799] = 62'b11111110110110101111110001101100111110011110011011000100101001;
  assign mem[800] = 62'b11111110101101110101000000011011111001100000001000111011001001;
  assign mem[801] = 62'b11111111101111111100100001011000010100111000010011000111101101;
  assign mem[802] = 62'b11111111100111111010000011111110000111101100000011011010000110;
  assign mem[803] = 62'b11111111100101010001010100111111110101000101011001110111111100;
  assign mem[804] = 62'b11111111011011111001010001010100010111111111111100000011011001;
  assign mem[805] = 62'b11111111101100110011001110111000100000110000101101111010100000;
  assign mem[806] = 62'b11111111101110001110100011001111101100011101011100111010000101;
  assign mem[807] = 62'b11111111010101000000010110001111011100000110010111000001001000;
  assign mem[808] = 62'b11111111010000000111110001100000000110101110011111110111010010;
  assign mem[809] = 62'b11111111101110111101111101011011100101000111001010001111000000;
  assign mem[810] = 62'b11111111101011100110001111101000011111110110010001010101011110;
  assign mem[811] = 62'b11111111100000001100101010111001010101111011011011110110010110;
  assign mem[812] = 62'b11111111100011010011000101001001010010110000010100110111100001;
  assign mem[813] = 62'b11111111101001100001101010111011110001010001010111010110010100;
  assign mem[814] = 62'b11111111101111101100100000110111000110100000011101010101001101;
  assign mem[815] = 62'b11111111000001100111011000100101000000101111100010010011100111;
  assign mem[816] = 62'b11111111000011111100100010111101010111110110110100100010010011;
  assign mem[817] = 62'b11111111101111100110111110110101111100111110111101111000101001;
  assign mem[818] = 62'b11111111101001111000001000001011101101101101000010010001110010;
  assign mem[819] = 62'b11111111100010110100110011001111010011010011101001101110111000;
  assign mem[820] = 62'b11111111100000101101000000010110000111100011111000010111101100;
  assign mem[821] = 62'b11111111101011010010110111010000001001110111100111100100100101;
  assign mem[822] = 62'b11111111101111000111000111101010111110001010000100011100001000;
  assign mem[823] = 62'b11111111001101111101010001011000111111000000010000100110011010;
  assign mem[824] = 62'b11111111010110000111010101100101011100100010001100001000000010;
  assign mem[825] = 62'b11111111101110000001110110011011011001001010000000111101010100;
  assign mem[826] = 62'b11111111101101000011010110011100101111010110011101001010111001;
  assign mem[827] = 62'b11111111011010110101000111001100010010010111001101110000001001;
  assign mem[828] = 62'b11111111100101101101010000101100100110010011110111010001001000;
  assign mem[829] = 62'b11111111100111100000101111101100011011100100001011001101011011;
  assign mem[830] = 62'b11111111101111111110010111110001000010000010001100000000010100;
  assign mem[831] = 62'b11111110100100011010100011100101101111111110000110000101111001;
  assign mem[832] = 62'b11111110100001010001101000010111011011010000101100000101111111;
  assign mem[833] = 62'b11111111101111111110110101010111100100001001011111110110101110;
  assign mem[834] = 62'b11111111100111011000001100010100101100001100000100011101100100;
  assign mem[835] = 62'b11111111100101110110011101111011100111001111100011010001011100;
  assign mem[836] = 62'b11111111011010011110010000110011010011110110111111001100011011;
  assign mem[837] = 62'b11111111101101001000100101010111000110111001011010010011100001;
  assign mem[838] = 62'b11111111101101111101011110001101101010100110111010010110011100;
  assign mem[839] = 62'b11111111010110011110111001010010011100101011010110001111001011;
  assign mem[840] = 62'b11111111001101001100010111011101001101001011001011110111101110;
  assign mem[841] = 62'b11111111101111001010000001011111111100010001100000100111001110;
  assign mem[842] = 62'b11111111101011001100010001010110100101111100110111101111110011;
  assign mem[843] = 62'b11111111100000110111101101000010111000010010111100010010110110;
  assign mem[844] = 62'b11111111100010101010100111011011101000011110101110101101011000;
  assign mem[845] = 62'b11111111101001111111011111010011110001001100010100100111011110;
  assign mem[846] = 62'b11111111101111100100111111000101001111100001011010110000001000;
  assign mem[847] = 62'b11111111000100101110001011000101111111011110011111101010001000;
  assign mem[848] = 62'b11111111000000110101100100110110111100101100100110011110000110;
  assign mem[849] = 62'b11111111101111101110001101000110001101011001101010110110110111;
  assign mem[850] = 62'b11111111101001011010000011111101000010101111010111111111100001;
  assign mem[851] = 62'b11111111100011011101000101001100011011100000010111111110001101;
  assign mem[852] = 62'b11111111100000000001110100000011001000001010111000001011100001;
  assign mem[853] = 62'b11111111101011101100100100100110100000101101101100010000001101;
  assign mem[854] = 62'b11111111101110111010110000011101001100010100001010010101000100;
  assign mem[855] = 62'b11111111010000100000000100111000000101111010110110011000011110;
  assign mem[856] = 62'b11111111010100101000100101001111010001000110111000001011110011;
  assign mem[857] = 62'b11111111101110010010101000110111111111100000011100111001011110;
  assign mem[858] = 62'b11111111101100101101101110001000001010000000001101101010011001;
  assign mem[859] = 62'b11111111011100001111110110110101000111001001100011000100101001;
  assign mem[860] = 62'b11111111100101000111111010100000011100110110011001101010100110;
  assign mem[861] = 62'b11111111101000000010011000101101110101011011100101001011111010;
  assign mem[862] = 62'b11111111101111111011110000000100000010100000100110000110010001;
  assign mem[863] = 62'b11111110110000011110110110000101001110010001100011000001100100;
  assign mem[864] = 62'b11111110110101001011100111011101001010010011010100110100001010;
  assign mem[865] = 62'b11111111101111111000111110100100101011111010011101100010000110;
  assign mem[866] = 62'b11111111101000011011000000101000011101100110101010000110010101;
  assign mem[867] = 62'b11111111100100101011010111100101010001011001110010001011110001;
  assign mem[868] = 62'b11111111011101010011001101000000101011101010000110000010011101;
  assign mem[869] = 62'b11111111101100011100110001010110001001100111101010101011010111;
  assign mem[870] = 62'b11111111101110011110011101101100101001101001010001011001011010;
  assign mem[871] = 62'b11111111010011100000111111010111100011010100111011011010101011;
  assign mem[872] = 62'b11111111010001101000101111011111111011111010001111001001000011;
  assign mem[873] = 62'b11111111101110110000101100111101001011000110101111011010110010;
  assign mem[874] = 62'b11111111101011111111001001110100100101101000011011000101000111;
  assign mem[875] = 62'b11111111011111000010000001100100000110101111111111011111111110;
  assign mem[876] = 62'b11111111100011111010110011001111101010101111100000011010000000;
  assign mem[877] = 62'b11111111101001000010110111100101000011010101110101111011111110;
  assign mem[878] = 62'b11111111101111110010110100011100000011100100010100001101010100;
  assign mem[879] = 62'b11111110111100111111110101001100111011001100000111110111000001;
  assign mem[880] = 62'b11111111000111000010101111110110001101000010001100010011111111;
  assign mem[881] = 62'b11111111101111011110100010100110011100000110100011001000101010;
  assign mem[882] = 62'b11111111101010010101001100100100010000100100001111010100100011;
  assign mem[883] = 62'b11111111100010001011110010110101100110001011000001001111100010;
  assign mem[884] = 62'b11111111100001010111100011011011100100110110111110001010111100;
  assign mem[885] = 62'b11111111101010111000000110100011110011010001011110110011101111;
  assign mem[886] = 62'b11111111101111010010010010001000000110101111001010101110110100;
  assign mem[887] = 62'b11111111001010111001001111000111010101111100111011100110101011;
  assign mem[888] = 62'b11111111010111100101001111010111100110000100111101111110101110;
  assign mem[889] = 62'b11111111101101101111111001111001000011100101010111010110011010;
  assign mem[890] = 62'b11111111101101010111110111000101110010100010001000101001111111;
  assign mem[891] = 62'b11111111011001011001010101010110110111101010111001010010001111;
  assign mem[892] = 62'b11111111100110010001110001010101000011011111110101001101011011;
  assign mem[893] = 62'b11111111100110111110001100101010011001110010010101101101110101;
  assign mem[894] = 62'b11111111101111111111110000100101000011110001010011101111010001;
  assign mem[895] = 62'b11111110001111011010100010100101101010101110011001011111001011;
  assign mem[896] = 62'b11111110010101111111010100110100100001111110101011001000100110;
  assign mem[897] = 62'b11111111101111111111100001110001101000011100001100101101110111;
  assign mem[898] = 62'b11111111100111000110111010110010010110000011100100000110111111;
  assign mem[899] = 62'b11111111100110001000101110010001001111111011000010001011111111;
  assign mem[900] = 62'b11111111011001110000010111110101000100000011011111100111110010;
  assign mem[901] = 62'b11111111101101010010110101101100011011000110000111010100100100;
  assign mem[902] = 62'b11111111101101110100011111111011110011100010101001000101011010;
  assign mem[903] = 62'b11111111010111001101110110001111001001001001100001000010010010;
  assign mem[904] = 62'b11111111001011101010010110001100110100111100010101110110101101;
  assign mem[905] = 62'b11111111101111001111100110101110111100000110111011110001100101;
  assign mem[906] = 62'b11111111101010111110111000111111011000100111110101011110110110;
  assign mem[907] = 62'b11111111100001001100111110100111001111111011100010010101001111;
  assign mem[908] = 62'b11111111100010010110000111001101001100101110110111000100010000;
  assign mem[909] = 62'b11111111101010001110000001100001001010010110010011101111000110;
  assign mem[910] = 62'b11111111101111100000110000111101001010010000001100011000001100;
  assign mem[911] = 62'b11111111000110010001010001101010000011000111011000001100001101;
  assign mem[912] = 62'b11111110111110100011101011011111111101111001001010101000111111;
  assign mem[913] = 62'b11111111101111110001010110111000111011011111011001101011110110;
  assign mem[914] = 62'b11111111101001001010101010010000011111110001011010100000010101;
  assign mem[915] = 62'b11111111100011110000111100010001001001100000011100010100011000;
  assign mem[916] = 62'b11111111011111010111111101111011100110010101101100110110100011;
  assign mem[917] = 62'b11111111101011111001000001101101100001000100010101010011000001;
  assign mem[918] = 62'b11111111101110110100001000001101011110100110011001000000001001;
  assign mem[919] = 62'b11111111010001010000100011111011101111110001101001001101111000;
  assign mem[920] = 62'b11111111010011111000111001101111101001011011101100001001110001;
  assign mem[921] = 62'b11111111101110011010100110000111000101010111010101001110100111;
  assign mem[922] = 62'b11111111101100100010011111010110000111000000101001110000010011;
  assign mem[923] = 62'b11111111011100111100110100101110101110111000011100110100100001;
  assign mem[924] = 62'b11111111100100110100111011110001101101010110001001111101111111;
  assign mem[925] = 62'b11111111101000010010110111000100010001101011111000001111111010;
  assign mem[926] = 62'b11111111101111111001111110101010000101010010000010110101100000;
  assign mem[927] = 62'b11111110110011100111011001111100010010110001011010001010011001;
  assign mem[928] = 62'b11111110110010000011001001011001110100111011010100010001001101;
  assign mem[929] = 62'b11111111101111111010111001110100100101001100000100000100001111;
  assign mem[930] = 62'b11111111101000001010101001110000010011111101010100010111111111;
  assign mem[931] = 62'b11111111100100111110011100110000100101110011001010010010000110;
  assign mem[932] = 62'b11111111011100100110010111111111000011100001100101001110001001;
  assign mem[933] = 62'b11111111101100101000001000111100011001101110011100010001001001;
  assign mem[934] = 62'b11111111101110010110101001110101010101000001000110011111010011;
  assign mem[935] = 62'b11111111010100010000110001000011011100100010010011011011110000;
  assign mem[936] = 62'b11111111010000111000010101101101001110000101110100100111001110;
  assign mem[937] = 62'b11111111101110110111011110101101101010000001111000011001010001;
  assign mem[938] = 62'b11111111101011110010110101010011001011000011010010001100100111;
  assign mem[939] = 62'b11111111011111101101110101011101011100001001001101001011011110;
  assign mem[940] = 62'b11111111100011100111000010001111100011110101100011000000101001;
  assign mem[941] = 62'b11111111101001010010011001000011100011101011000100101001101100;
  assign mem[942] = 62'b11111111101111101111110100011100001111000010101000110110001000;
  assign mem[943] = 62'b11111111000000000011101110100010101101011011111011100001011011;
  assign mem[944] = 62'b11111111000101011111110000000010000110010101001100101111011110;
  assign mem[945] = 62'b11111111101111100010111010011100110111110010110100101101111000;
  assign mem[946] = 62'b11111111101010000110110010011011010010110000001010011101011110;
  assign mem[947] = 62'b11111111100010100000011000101111101111010011010011110010111010;
  assign mem[948] = 62'b11111111100001000010010111001001001000110100001010100101010111;
  assign mem[949] = 62'b11111111101011000101100111010000101010010011001010001011110101;
  assign mem[950] = 62'b11111111101111001100110110100001011010001110101010111011110000;
  assign mem[951] = 62'b11111111001100011011011001000001010011010111010111010011011101;
  assign mem[952] = 62'b11111111010110110110011001100001100011100010100000110010110110;
  assign mem[953] = 62'b11111111101101111001000001011000001111011011011000110110000001;
  assign mem[954] = 62'b11111111101101001101101111110001111011110010111111101111011100;
  assign mem[955] = 62'b11111111011010000111010110010101000011101101010000101011000000;
  assign mem[956] = 62'b11111111100101111111100111110010111101111001010110101000010000;
  assign mem[957] = 62'b11111111100111001111100101010110001110000001111001100101000010;
  assign mem[958] = 62'b11111111101111111111001110000010011100111000101010011001111001;
  assign mem[959] = 62'b11111110011100010001010100111101001100111001010011101100011101;
  assign mem[960] = 62'b11111110100111100011011011101010100101100001110100011010000110;
  assign mem[961] = 62'b11111111101111111101110101001110111011000110111001000101100100;
  assign mem[962] = 62'b11111111100111101001001111011100000111101111111001011111010010;
  assign mem[963] = 62'b11111111100101100100000000000111010101111101110010001111011111;
  assign mem[964] = 62'b11111111011011001011111001011100011101101100110001100101110010;
  assign mem[965] = 62'b11111111101100111110000011000011101000110011100100011001111011;
  assign mem[966] = 62'b11111111101110000110001010000000101111110111000110011011011001;
  assign mem[967] = 62'b11111111010101101111101110011110001011100111011011001110110110;
  assign mem[968] = 62'b11111111001110101110000110101101000110001011011110001101001000;
  assign mem[969] = 62'b11111111101111000100001001000010111100100010011000111101011111;
  assign mem[970] = 62'b11111111101011011001011000111100010100111111011011110001000111;
  assign mem[971] = 62'b11111111100000100010010001000100100000001100101011000010001100;
  assign mem[972] = 62'b11111111100010111110111100001001001011010001000001000000010101;
  assign mem[973] = 62'b11111111101001110000101101000100010000111100000111010111000010;
  assign mem[974] = 62'b11111111101111101000111001101110101100011110100001011110010001;
  assign mem[975] = 62'b11111111000011001010110111101111111001010001010001011010100111;
  assign mem[976] = 62'b11111111000010011001001001100101001101111111010011010000001001;
  assign mem[977] = 62'b11111111101111101010101111101111001011000011001111110111011100;
  assign mem[978] = 62'b11111111101001101001001101111110100100001010110000011010110010;
  assign mem[979] = 62'b11111111100011001001000010000111101100010010011010011000011111;
  assign mem[980] = 62'b11111111100000010111011111001111101100001100011011100010110111;
  assign mem[981] = 62'b11111111101011011111110110011010000110111001111001001011101001;
  assign mem[982] = 62'b11111111101111000001000101101000010100110011110111001110001100;
  assign mem[983] = 62'b11111111001111011110110111010010000000101111010011100000000010;
  assign mem[984] = 62'b11111111010101011000000100000000010010111101000110011110110100;
  assign mem[985] = 62'b11111111101110001010011000111101000100001110010001100101111010;
  assign mem[986] = 62'b11111111101100111000101011001100100111100110011010000001100000;
  assign mem[987] = 62'b11111111011011100010100111100000010100111111010101011010010011;
  assign mem[988] = 62'b11111111100101011010101100001101010001100101110110010010011111;
  assign mem[989] = 62'b11111111100111110001101011100010011100111000101101001100110011;
  assign mem[990] = 62'b11111111101111111101001101110001010100101100011011111011010011;
  assign mem[991] = 62'b11111110101010101100010000000110111101010111111000001100010111;
  assign mem[992] = 62'b11111110111000010011111000011100010010110000010011000010100001;
  assign mem[993] = 62'b11111111101111110110101111101001110101000101000101001110001100;
  assign mem[994] = 62'b11111111101000101011001000011100011110110111100001110110001000;
  assign mem[995] = 62'b11111111100100011000000101101001101001001010110011001010100010;
  assign mem[996] = 62'b11111111011101111111101111111101100110101010010100000111011110;
  assign mem[997] = 62'b11111111101100010001001000001100110001010000011100000000000100;
  assign mem[998] = 62'b11111111101110100101111110110000110110000000010110101100110000;
  assign mem[999] = 62'b11111111010010110001000001101001001110100101010100010100100000;
  assign mem[1000] = 62'b11111111010010011000111110011010011001010101010101010010111010;
  assign mem[1001] = 62'b11111111101110101001101000001110010011111001100101100000000000;
  assign mem[1002] = 62'b11111111101100001011001101000101001001001100011110001111110001;
  assign mem[1003] = 62'b11111111011110010101111010100001101101001111001101100000100101;
  assign mem[1004] = 62'b11111111100100001110010111111101011011001010100100001110000000;
  assign mem[1005] = 62'b11111111101000110011000110101001110101000110000100011001010101;
  assign mem[1006] = 62'b11111111101111110101100000110100101101101001110101110010011110;
  assign mem[1007] = 62'b11111110111001110111111011011011101011001001001010100001011100;
  assign mem[1008] = 62'b11111111001000100101100001011100100111110001000001100000000100;
  assign mem[1009] = 62'b11111111101111011001110111010101010110100010000011110011101110;
  assign mem[1010] = 62'b11111111101010100011010110011101101110010101000101101011010010;
  assign mem[1011] = 62'b11111111100001110111000001101101100100110111000100100001110010;
  assign mem[1012] = 62'b11111111100001101100100101000000010111000100110111001110111111;
  assign mem[1013] = 62'b11111111101010101010010101010001111010001011001011100110001110;
  assign mem[1014] = 62'b11111111101111010111011010011011101101010000110110100001011101;
  assign mem[1015] = 62'b11111111001001010110110100100111101001101101100010101011111010;
  assign mem[1016] = 62'b11111111011000010011110110101010101010111100111001000000111111;
  assign mem[1017] = 62'b11111111101101100110100000000011011101100010110011110101000110;
  assign mem[1018] = 62'b11111111101101100001101100010010000100010001011010010001001111;
  assign mem[1019] = 62'b11111111011000101011000100101110000110110101011110110101000100;
  assign mem[1020] = 62'b11111111100110100011101101000111101010101000011001110001110001;
  assign mem[1021] = 62'b11111111100110101100100101110011101101001011111110001010011100;
  assign mem[1022] = 62'b11111111101111111111111111011000100001011000100001110100000010;
  assign mem[1023] = 62'b11111101101001001000011111100010111110110011001010010010111010;
  always@(*)
  begin
    data_out_t <= mem[addr_f];
  end
  wire [61:0] data_out_reg [n_outreg:0];
  generate if (n_outreg > 0)
  begin
    for( i=n_outreg-1; i >= 1; i=i-1)
    begin: data_out_reg_stage
      mgc_generic_reg #(
        .width(62),
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_data_out_reg (
        .d(data_out_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(data_out_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(62),
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_data_out_reg_init (
      .d(data_out_t),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(data_out_reg[0])
    );
    assign data_out = data_out_reg[n_outreg-1];
  end
  else
  begin
    assign data_out = data_out_t;
  end
  endgenerate
endmodule
module stagemgc_rom_sync_regout_9_1024_64_1_0_0_1_0_1_0_0_0_1_60 (addr, data_out,
    clk, s_rst, a_rst, en
);
  input [9:0]addr ;
  output [63:0]data_out ;
  input clk ;
  input s_rst ;
  input a_rst ;
  input en ;
  parameter n_width = 64;
  parameter n_size = 1024;
  parameter n_numports = 1;
  parameter n_addr_w = 10;
  parameter n_inreg = 0;
  parameter n_outreg = 1;
  wire [9:0] addr_f;
  wire [9:0] addr_reg [n_inreg:0];
  genvar i;
  generate if (n_inreg > 0)
  begin
    for( i=n_inreg-1; i >= 1; i=i-1)
    begin: addr_reg_stage
      mgc_generic_reg #(
        .width(10),
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_addr_reg (
        .d(addr_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(addr_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(10),
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_addr_reg_init (
      .d(addr),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(addr_reg[0])
    );
    assign addr_f = addr_reg[n_inreg-1];
  end
  else
  begin
    assign addr_f = addr;
  end
  endgenerate
  wire [63:0] mem [1023:0];
  reg [63:0] data_out_t;
  assign mem[0] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  assign mem[1] = 64'b1000000000000000000000000000000000000000000000000000000000000000;
  assign mem[2] = 64'b0011111111100110101000001001111001100110011111110011101111001101;
  assign mem[3] = 64'b1011111111100110101000001001111001100110011111110011101111001101;
  assign mem[4] = 64'b0011111111101101100100000110101111001111001100101000110101000110;
  assign mem[5] = 64'b1011111111011000011111011110001010100110101011101010100101100011;
  assign mem[6] = 64'b0011111111011000011111011110001010100110101011101010100101100011;
  assign mem[7] = 64'b1011111111101101100100000110101111001111001100101000110101000110;
  assign mem[8] = 64'b0011111111101111011000101001011111001111111101110101110010110000;
  assign mem[9] = 64'b1011111111001000111110001011100000111100011010011010011000001011;
  assign mem[10] = 64'b0011111111100001110001110011101100111001101011100110100011001000;
  assign mem[11] = 64'b1011111111101010100110110110011000101001000011101010000110100011;
  assign mem[12] = 64'b0011111111101010100110110110011000101001000011101010000110100011;
  assign mem[13] = 64'b1011111111100001110001110011101100111001101011100110100011001000;
  assign mem[14] = 64'b0011111111001000111110001011100000111100011010011010011000001011;
  assign mem[15] = 64'b1011111111101111011000101001011111001111111101110101110010110000;
  assign mem[16] = 64'b0011111111101111110110001000110110100011110100010010010100100110;
  assign mem[17] = 64'b1011111110111001000101111010011010111100001010011011010000101100;
  assign mem[18] = 64'b0011111111100100010011001111001100100101000010010001110111010110;
  assign mem[19] = 64'b1011111111101000101111001000000001101011000101010001011101000001;
  assign mem[20] = 64'b0011111111101100001110001011001011110001100000001011110110110001;
  assign mem[21] = 64'b1011111111011110001010110101110100111000000001101111011000111011;
  assign mem[22] = 64'b0011111111010010100101000000011000101110110101011001111100000110;
  assign mem[23] = 64'b1011111111101110100111110100000101010110110001100010110111011010;
  assign mem[24] = 64'b0011111111101110100111110100000101010110110001100010110111011010;
  assign mem[25] = 64'b1011111111010010100101000000011000101110110101011001111100000110;
  assign mem[26] = 64'b0011111111011110001010110101110100111000000001101111011000111011;
  assign mem[27] = 64'b1011111111101100001110001011001011110001100000001011110110110001;
  assign mem[28] = 64'b0011111111101000101111001000000001101011000101010001011101000001;
  assign mem[29] = 64'b1011111111100100010011001111001100100101000010010001110111010110;
  assign mem[30] = 64'b0011111110111001000101111010011010111100001010011011010000101100;
  assign mem[31] = 64'b1011111111101111110110001000110110100011110100010010010100100110;
  assign mem[32] = 64'b0011111111101111111101100010000111100011011110010110110101111110;
  assign mem[33] = 64'b1011111110101001000111110110010111110001000011011101100000010100;
  assign mem[34] = 64'b0011111111100101011111010110100100110100100011001110110010100000;
  assign mem[35] = 64'b1011111111100111101101011101111100100010011010101010111110101111;
  assign mem[36] = 64'b0011111111101100111011010111101011110100001111001100011101110011;
  assign mem[37] = 64'b1011111111011011010111010001000000001001111000010101110011000000;
  assign mem[38] = 64'b0011111111010101100011111001101001110101101010110001111111011101;
  assign mem[39] = 64'b1011111111101110001000010010000100000100111101101000011011100101;
  assign mem[40] = 64'b0011111111101111000010100111111011111011100100100011000011010111;
  assign mem[41] = 64'b1011111111001111000110011111100101111011001000010101111100011011;
  assign mem[42] = 64'b0011111111100000011100111000011110011001001000101111111111101110;
  assign mem[43] = 64'b1011111111101011011100101000001101000101000110010110111000111110;
  assign mem[44] = 64'b0011111111101001101100111110000001000111111100111000011101000001;
  assign mem[45] = 64'b1011111111100011000011111111011111111100111000010111000000110101;
  assign mem[46] = 64'b0011111111000010110010000001000001101110100011100110000100111010;
  assign mem[47] = 64'b1011111111101111101001110101010101111111000010001010010100010111;
  assign mem[48] = 64'b0011111111101111101001110101010101111111000010001010010100010111;
  assign mem[49] = 64'b1011111111000010110010000001000001101110100011100110000100111010;
  assign mem[50] = 64'b0011111111100011000011111111011111111100111000010111000000110101;
  assign mem[51] = 64'b1011111111101001101100111110000001000111111100111000011101000001;
  assign mem[52] = 64'b0011111111101011011100101000001101000101000110010110111000111110;
  assign mem[53] = 64'b1011111111100000011100111000011110011001001000101111111111101110;
  assign mem[54] = 64'b0011111111001111000110011111100101111011001000010101111100011011;
  assign mem[55] = 64'b1011111111101111000010100111111011111011100100100011000011010111;
  assign mem[56] = 64'b0011111111101110001000010010000100000100111101101000011011100101;
  assign mem[57] = 64'b1011111111010101100011111001101001110101101010110001111111011101;
  assign mem[58] = 64'b0011111111011011010111010001000000001001111000010101110011000000;
  assign mem[59] = 64'b1011111111101100111011010111101011110100001111001100011101110011;
  assign mem[60] = 64'b0011111111100111101101011101111100100010011010101010111110101111;
  assign mem[61] = 64'b1011111111100101011111010110100100110100100011001110110010100000;
  assign mem[62] = 64'b0011111110101001000111110110010111110001000011011101100000010100;
  assign mem[63] = 64'b1011111111101111111101100010000111100011011110010110110101111110;
  assign mem[64] = 64'b0011111111101111111111011000100001100000100001001100110100001101;
  assign mem[65] = 64'b1011111110011001001000010101010111110111101000110110011001111110;
  assign mem[66] = 64'b0011111111100110000100001011011101010101000111010010110011011111;
  assign mem[67] = 64'b1011111111100111001011010000100000110111111011111111111110010110;
  assign mem[68] = 64'b0011111111101101010000010011010011010001010011011100100100111010;
  assign mem[69] = 64'b1011111111011001111011110111100101000011101010001110110110001010;
  assign mem[70] = 64'b0011111111010111000010001000010100110000111110100100010110011111;
  assign mem[71] = 64'b1011111111101101110110110001001110110110110011001100001000111100;
  assign mem[72] = 64'b0011111111101111001110001111001110101100011001001110010110001001;
  assign mem[73] = 64'b1011111111001100000010111000001001101010011111100100111101100011;
  assign mem[74] = 64'b0011111111100001000111101011001101010100000110110100101100100011;
  assign mem[75] = 64'b1011111111101011000010010000101001011000000101010000001000000000;
  assign mem[76] = 64'b0011111111101010001010011010011110100000010001100010011110000010;
  assign mem[77] = 64'b1011111111100010011011010000010101001100110111010001001011011111;
  assign mem[78] = 64'b0011111111000101111000100001010001000100100010110011111111000110;
  assign mem[79] = 64'b1011111111101111100001110110010011111010011100010100101110101001;
  assign mem[80] = 64'b0011111111101111110000100110010001110000111000011001111111010011;
  assign mem[81] = 64'b1011111110111111010101100100111001010110101010010111001100001110;
  assign mem[82] = 64'b0011111111100011101011111111101000101001001000000101000010111001;
  assign mem[83] = 64'b1011111111101001001110100010001001001001100100100110001111111011;
  assign mem[84] = 64'b0011111111101011110101111100000010101100011011111001010100101010;
  assign mem[85] = 64'b1011111111011111100010111010010011011011111110001001101010111010;
  assign mem[86] = 64'b0011111111010001000100011101001001100010101100011111011001110111;
  assign mem[87] = 64'b1011111111101110110101110100000011100111011010000100100101100011;
  assign mem[88] = 64'b0011111111101110011000101000100011101100010010001110000100010010;
  assign mem[89] = 64'b1011111111010100000100110101110010010100000101110110011000000001;
  assign mem[90] = 64'b0011111111011100110001100110111010011001001100011100010001011110;
  assign mem[91] = 64'b1011111111101100100101010100101100100001001101000001000111110101;
  assign mem[92] = 64'b0011111111101000001110110000111000001011111111111001011101101110;
  assign mem[93] = 64'b1011111111100100111001101100101010111011111000111110010111101001;
  assign mem[94] = 64'b0011111110110010110101010010000010010010110011100001100111110110;
  assign mem[95] = 64'b1011111111101111111010011100110110101101000000011000100000111010;
  assign mem[96] = 64'b0011111111101111111010011100110110101101000000011000100000111010;
  assign mem[97] = 64'b1011111110110010110101010010000010010010110011100001100111110110;
  assign mem[98] = 64'b0011111111100100111001101100101010111011111000111110010111101001;
  assign mem[99] = 64'b1011111111101000001110110000111000001011111111111001011101101110;
  assign mem[100] = 64'b0011111111101100100101010100101100100001001101000001000111110101;
  assign mem[101] = 64'b1011111111011100110001100110111010011001001100011100010001011110;
  assign mem[102] = 64'b0011111111010100000100110101110010010100000101110110011000000001;
  assign mem[103] = 64'b1011111111101110011000101000100011101100010010001110000100010010;
  assign mem[104] = 64'b0011111111101110110101110100000011100111011010000100100101100011;
  assign mem[105] = 64'b1011111111010001000100011101001001100010101100011111011001110111;
  assign mem[106] = 64'b0011111111011111100010111010010011011011111110001001101010111010;
  assign mem[107] = 64'b1011111111101011110101111100000010101100011011111001010100101010;
  assign mem[108] = 64'b0011111111101001001110100010001001001001100100100110001111111011;
  assign mem[109] = 64'b1011111111100011101011111111101000101001001000000101000010111001;
  assign mem[110] = 64'b0011111110111111010101100100111001010110101010010111001100001110;
  assign mem[111] = 64'b1011111111101111110000100110010001110000111000011001111111010011;
  assign mem[112] = 64'b0011111111101111100001110110010011111010011100010100101110101001;
  assign mem[113] = 64'b1011111111000101111000100001010001000100100010110011111111000110;
  assign mem[114] = 64'b0011111111100010011011010000010101001100110111010001001011011111;
  assign mem[115] = 64'b1011111111101010001010011010011110100000010001100010011110000010;
  assign mem[116] = 64'b0011111111101011000010010000101001011000000101010000001000000000;
  assign mem[117] = 64'b1011111111100001000111101011001101010100000110110100101100100011;
  assign mem[118] = 64'b0011111111001100000010111000001001101010011111100100111101100011;
  assign mem[119] = 64'b1011111111101111001110001111001110101100011001001110010110001001;
  assign mem[120] = 64'b0011111111101101110110110001001110110110110011001100001000111100;
  assign mem[121] = 64'b1011111111010111000010001000010100110000111110100100010110011111;
  assign mem[122] = 64'b0011111111011001111011110111100101000011101010001110110110001010;
  assign mem[123] = 64'b1011111111101101010000010011010011010001010011011100100100111010;
  assign mem[124] = 64'b0011111111100111001011010000100000110111111011111111111110010110;
  assign mem[125] = 64'b1011111111100110000100001011011101010101000111010010110011011111;
  assign mem[126] = 64'b0011111110011001001000010101010111110111101000110110011001111110;
  assign mem[127] = 64'b1011111111101111111111011000100001100000100001001100110100001101;
  assign mem[128] = 64'b0011111111101111111111110110001000010110100110111001001011011011;
  assign mem[129] = 64'b1011111110001001001000011101000111111100110111101100011110000100;
  assign mem[130] = 64'b0011111111100110010110010001100100100101111100000111100000111101;
  assign mem[131] = 64'b1011111111100110111001110100010001010100111010101010100010101111;
  assign mem[132] = 64'b0011111111101101011010010110000101110011110010011110011010001011;
  assign mem[133] = 64'b1011111111011001001101110010101001100011101111001001001111010111;
  assign mem[134] = 64'b0011111111010111110000111010100100110001000111011100110011100111;
  assign mem[135] = 64'b1011111111101101101101100101001001100010001110001010000010011011;
  assign mem[136] = 64'b0011111111101111010011100110000000111011000010110010111100101101;
  assign mem[137] = 64'b1011111111001010100000101010000000100101101100000000010001010001;
  assign mem[138] = 64'b0011111111100001011100110100110101100011110111101101101101001001;
  assign mem[139] = 64'b1011111111101010110100101011110010011110001000011101010100010001;
  assign mem[140] = 64'b0011111111101010011000110000100100011011000000101111101011100010;
  assign mem[141] = 64'b1011111111100010000110100111100110011001001100111110101101011001;
  assign mem[142] = 64'b0011111111000111011011011101100111011110010100001011111100110001;
  assign mem[143] = 64'b1011111111101111011101011001100110100011101000010010000001110111;
  assign mem[144] = 64'b0011111111101111110011100001010111111101011011011010011001111011;
  assign mem[145] = 64'b1011111110111100001101111000010111000111100111101100001011010101;
  assign mem[146] = 64'b0011111111100011111111101101100101010011010001010101011011010100;
  assign mem[147] = 64'b1011111111101000111110111100110010100011111011111001010000001101;
  assign mem[148] = 64'b0011111111101100000010001100010000100110011100100101010101001001;
  assign mem[149] = 64'b1011111111011110110111000001100101010010111011110111100011010110;
  assign mem[150] = 64'b0011111111010001110100110100010000111111010011001101101100111110;
  assign mem[151] = 64'b1011111111101110101110111101100011001000110111110000101101110100;
  assign mem[152] = 64'b0011111111101110100000010111101110101011010011001101000100001101;
  assign mem[153] = 64'b1011111111010011010101000001000011000010111000011000000101010010;
  assign mem[154] = 64'b0011111111011101011110010111011101011011100001101110001110001001;
  assign mem[155] = 64'b1011111111101100011001111000101100110100100010000111001110011011;
  assign mem[156] = 64'b0011111111101000011111000100000000001111101110100010111010111111;
  assign mem[157] = 64'b1011111111100100100110100100010010011011100110110000100100111001;
  assign mem[158] = 64'b0011111110110101111101101101000000001010100110101010010000011001;
  assign mem[159] = 64'b1011111111101111111000011100101011111100101111010101101100001001;
  assign mem[160] = 64'b0011111111101111111100001001010101100101100011100111000110101101;
  assign mem[161] = 64'b1011111110101111011001010110111001111001111110000010000011100000;
  assign mem[162] = 64'b0011111111100101001100101000001010010010101000110101010110010110;
  assign mem[163] = 64'b1011111111100111111110001110110011100011010101110001011101110001;
  assign mem[164] = 64'b0011111111101100110000011111000011110011111111001111110001011100;
  assign mem[165] = 64'b1011111111011100000100100100100111011000000000010001111011100111;
  assign mem[166] = 64'b0011111111010100110100011110001001000010011110001110011101101010;
  assign mem[167] = 64'b1011111111101110010000100110101001001011001010111100000101111110;
  assign mem[168] = 64'b0011111111101110111100010111100010100011111001000111001111000010;
  assign mem[169] = 64'b1011111111010000010011111011100000001110001101111111110110101110;
  assign mem[170] = 64'b0011111111100000000111001111110010000111010011000011111010110111;
  assign mem[171] = 64'b1011111111101011101001011010101001100111001101011001000011010010;
  assign mem[172] = 64'b0011111111101001011101110111111011110100110001111101011101000010;
  assign mem[173] = 64'b1011111111100011011000000101100010110001000001100101100111110011;
  assign mem[174] = 64'b0011111111000001001110011111000011001110110110101111010101110111;
  assign mem[175] = 64'b1011111111101111101101010111100101110001100101011101011101000001;
  assign mem[176] = 64'b0011111111101111100101111111100100100100110010010000100110011011;
  assign mem[177] = 64'b1011111111000100010101010111011010110001001010010011111001011010;
  assign mem[178] = 64'b0011111111100010101111101101101100100101111110101111001111101010;
  assign mem[179] = 64'b1011111111101001111011110100001111101111001010011010111110010100;
  assign mem[180] = 64'b0011111111101011001111100100110100111110111101010101011100010010;
  assign mem[181] = 64'b1011111111100000110010010111000001001101010111011000100110001111;
  assign mem[182] = 64'b0011111111001101100100110100111111100101010001010100001100010001;
  assign mem[183] = 64'b1011111111101111001000100101001011110111011101100011101011011010;
  assign mem[184] = 64'b0011111111101101111111101010111001100010001011011011111000101011;
  assign mem[185] = 64'b1011111111010110010011000111110111011101001111110010011111000110;
  assign mem[186] = 64'b0011111111011010101001101100100000101011011011010011111111001010;
  assign mem[187] = 64'b1011111111101101000101111110011101110100001111100011010111011100;
  assign mem[188] = 64'b0011111111100111011100011110011101011111000000110111001001100001;
  assign mem[189] = 64'b1011111111100101110001110111101110111110011001010000000110001100;
  assign mem[190] = 64'b0011111110100010110110000110010101110101100101000101010111001101;
  assign mem[191] = 64'b1011111111101111111110100111001011101111111111101111011101011101;
  assign mem[192] = 64'b0011111111101111111110100111001011101111111111101111011101011101;
  assign mem[193] = 64'b1011111110100010110110000110010101110101100101000101010111001101;
  assign mem[194] = 64'b0011111111100101110001110111101110111110011001010000000110001100;
  assign mem[195] = 64'b1011111111100111011100011110011101011111000000110111001001100001;
  assign mem[196] = 64'b0011111111101101000101111110011101110100001111100011010111011100;
  assign mem[197] = 64'b1011111111011010101001101100100000101011011011010011111111001010;
  assign mem[198] = 64'b0011111111010110010011000111110111011101001111110010011111000110;
  assign mem[199] = 64'b1011111111101101111111101010111001100010001011011011111000101011;
  assign mem[200] = 64'b0011111111101111001000100101001011110111011101100011101011011010;
  assign mem[201] = 64'b1011111111001101100100110100111111100101010001010100001100010001;
  assign mem[202] = 64'b0011111111100000110010010111000001001101010111011000100110001111;
  assign mem[203] = 64'b1011111111101011001111100100110100111110111101010101011100010010;
  assign mem[204] = 64'b0011111111101001111011110100001111101111001010011010111110010100;
  assign mem[205] = 64'b1011111111100010101111101101101100100101111110101111001111101010;
  assign mem[206] = 64'b0011111111000100010101010111011010110001001010010011111001011010;
  assign mem[207] = 64'b1011111111101111100101111111100100100100110010010000100110011011;
  assign mem[208] = 64'b0011111111101111101101010111100101110001100101011101011101000001;
  assign mem[209] = 64'b1011111111000001001110011111000011001110110110101111010101110111;
  assign mem[210] = 64'b0011111111100011011000000101100010110001000001100101100111110011;
  assign mem[211] = 64'b1011111111101001011101110111111011110100110001111101011101000010;
  assign mem[212] = 64'b0011111111101011101001011010101001100111001101011001000011010010;
  assign mem[213] = 64'b1011111111100000000111001111110010000111010011000011111010110111;
  assign mem[214] = 64'b0011111111010000010011111011100000001110001101111111110110101110;
  assign mem[215] = 64'b1011111111101110111100010111100010100011111001000111001111000010;
  assign mem[216] = 64'b0011111111101110010000100110101001001011001010111100000101111110;
  assign mem[217] = 64'b1011111111010100110100011110001001000010011110001110011101101010;
  assign mem[218] = 64'b0011111111011100000100100100100111011000000000010001111011100111;
  assign mem[219] = 64'b1011111111101100110000011111000011110011111111001111110001011100;
  assign mem[220] = 64'b0011111111100111111110001110110011100011010101110001011101110001;
  assign mem[221] = 64'b1011111111100101001100101000001010010010101000110101010110010110;
  assign mem[222] = 64'b0011111110101111011001010110111001111001111110000010000011100000;
  assign mem[223] = 64'b1011111111101111111100001001010101100101100011100111000110101101;
  assign mem[224] = 64'b0011111111101111111000011100101011111100101111010101101100001001;
  assign mem[225] = 64'b1011111110110101111101101101000000001010100110101010010000011001;
  assign mem[226] = 64'b0011111111100100100110100100010010011011100110110000100100111001;
  assign mem[227] = 64'b1011111111101000011111000100000000001111101110100010111010111111;
  assign mem[228] = 64'b0011111111101100011001111000101100110100100010000111001110011011;
  assign mem[229] = 64'b1011111111011101011110010111011101011011100001101110001110001001;
  assign mem[230] = 64'b0011111111010011010101000001000011000010111000011000000101010010;
  assign mem[231] = 64'b1011111111101110100000010111101110101011010011001101000100001101;
  assign mem[232] = 64'b0011111111101110101110111101100011001000110111110000101101110100;
  assign mem[233] = 64'b1011111111010001110100110100010000111111010011001101101100111110;
  assign mem[234] = 64'b0011111111011110110111000001100101010010111011110111100011010110;
  assign mem[235] = 64'b1011111111101100000010001100010000100110011100100101010101001001;
  assign mem[236] = 64'b0011111111101000111110111100110010100011111011111001010000001101;
  assign mem[237] = 64'b1011111111100011111111101101100101010011010001010101011011010100;
  assign mem[238] = 64'b0011111110111100001101111000010111000111100111101100001011010101;
  assign mem[239] = 64'b1011111111101111110011100001010111111101011011011010011001111011;
  assign mem[240] = 64'b0011111111101111011101011001100110100011101000010010000001110111;
  assign mem[241] = 64'b1011111111000111011011011101100111011110010100001011111100110001;
  assign mem[242] = 64'b0011111111100010000110100111100110011001001100111110101101011001;
  assign mem[243] = 64'b1011111111101010011000110000100100011011000000101111101011100010;
  assign mem[244] = 64'b0011111111101010110100101011110010011110001000011101010100010001;
  assign mem[245] = 64'b1011111111100001011100110100110101100011110111101101101101001001;
  assign mem[246] = 64'b0011111111001010100000101010000000100101101100000000010001010001;
  assign mem[247] = 64'b1011111111101111010011100110000000111011000010110010111100101101;
  assign mem[248] = 64'b0011111111101101101101100101001001100010001110001010000010011011;
  assign mem[249] = 64'b1011111111010111110000111010100100110001000111011100110011100111;
  assign mem[250] = 64'b0011111111011001001101110010101001100011101111001001001111010111;
  assign mem[251] = 64'b1011111111101101011010010110000101110011110010011110011010001011;
  assign mem[252] = 64'b0011111111100110111001110100010001010100111010101010100010101111;
  assign mem[253] = 64'b1011111111100110010110010001100100100101111100000111100000111101;
  assign mem[254] = 64'b0011111110001001001000011101000111111100110111101100011110000100;
  assign mem[255] = 64'b1011111111101111111111110110001000010110100110111001001011011011;
  assign mem[256] = 64'b0011111111101111111111111101100010000101100011101000101010010010;
  assign mem[257] = 64'b1011111101111001001000011111000011111110011001110000000001110001;
  assign mem[258] = 64'b0011111111100110011111001111011110000100100100011010111100010000;
  assign mem[259] = 64'b1011111111100110110001000000110101110011110000011000001001110101;
  assign mem[260] = 64'b0011111111101101011111010000101100000010101110001110110011111001;
  assign mem[261] = 64'b1011111111011000110110101010010100101110110010001010010010110000;
  assign mem[262] = 64'b0011111111011000001000001110001110110000010011101010101011000100;
  assign mem[263] = 64'b1011111111101101101000111000001110101001011001101000100110001000;
  assign mem[264] = 64'b0011111111101111010110001010001010110001011110001001111010000100;
  assign mem[265] = 64'b1011111111001001101111011100101111110010110111000100001101100110;
  assign mem[266] = 64'b0011111111100001100111010101101000001001111100101011100110111000;
  assign mem[267] = 64'b1011111111101010101101110011001001011001000101101100000011010100;
  assign mem[268] = 64'b0011111111101010011111110101100001010010100111111110011010011101;
  assign mem[269] = 64'b1011111111100001111100001111000010001011101111001000011000011011;
  assign mem[270] = 64'b0011111111001000001100110110011011101000100111000110010011000110;
  assign mem[271] = 64'b1011111111101111011011000011111101111101111101011011101110110111;
  assign mem[272] = 64'b0011111111101111110100110111100100010100001000100000101110000100;
  assign mem[273] = 64'b1011111110111010101001111011011100100100010010010101110000000011;
  assign mem[274] = 64'b0011111111100100001001011111111100010111100011100110101110110001;
  assign mem[275] = 64'b1011111111101000110111000100010100110011000101101001100011001100;
  assign mem[276] = 64'b0011111111101100001000001101111000111111101010010111000110110000;
  assign mem[277] = 64'b1011111111011110100000111110000011101010111110000101000100010100;
  assign mem[278] = 64'b0011111111010010001100111011101110101011110000111011101101110001;
  assign mem[279] = 64'b1011111111101110101011011011001011101000111001111010100010001110;
  assign mem[280] = 64'b0011111111101110100100001000010000110110000111011111011111110010;
  assign mem[281] = 64'b1011111111010010111101000010001011011010111011000000001110000111;
  assign mem[282] = 64'b0011111111011101110100101000111100010100100000011100110001011000;
  assign mem[283] = 64'b1011111111101100010100000100001000000001001010110110100100000111;
  assign mem[284] = 64'b0011111111101000100111000111111010011010010011011101010010101010;
  assign mem[285] = 64'b1011111111100100011100111011010100011011100110000111001101000111;
  assign mem[286] = 64'b0011111110110111100001110101100001101010010111010101101100100001;
  assign mem[287] = 64'b1011111111101111110111010101001110011111111100011111010001010110;
  assign mem[288] = 64'b0011111111101111111100111000001100001111100011010101011101011100;
  assign mem[289] = 64'b1011111110101100010000101000110100010010110000001101011111100011;
  assign mem[290] = 64'b0011111111100101010110000001000000111000100101110101000100110111;
  assign mem[291] = 64'b1011111111100111110101111000001101101100110000110011110110110010;
  assign mem[292] = 64'b0011111111101100110101111101100110001001100010110011001011110110;
  assign mem[293] = 64'b1011111111011011101101111100111100100011000001001011110100000001;
  assign mem[294] = 64'b0011111111010101001100001101100010000000101011110011110000100100;
  assign mem[295] = 64'b1011111111101110001100011110101011101000011100001100111000100101;
  assign mem[296] = 64'b0011111111101110111111100010001000001100000010111001010111101100;
  assign mem[297] = 64'b1011111111001111110111001101110000011010110111111110110111111001;
  assign mem[298] = 64'b0011111111100000010010000101011000100110101011100010001000011010;
  assign mem[299] = 64'b1011111111101011100011000011100011010010011101010000010011101001;
  assign mem[300] = 64'b0011111111101001100101011100111100101110110110000000110100100010;
  assign mem[301] = 64'b1011111111100011001110000100000000001101000011001000111001010111;
  assign mem[302] = 64'b0011111111000010000000010001011011010100111011000111101111001111;
  assign mem[303] = 64'b1011111111101111101011101000111010001110010001101100111110111011;
  assign mem[304] = 64'b0011111111101111100111111100111001010101101011011011001011001000;
  assign mem[305] = 64'b1011111111000011100011101101101110110000110011011000110100010100;
  assign mem[306] = 64'b0011111111100010111001111000000011100011111010001110101000010111;
  assign mem[307] = 64'b1011111111101001110100011011000111110101111010101000000011010101;
  assign mem[308] = 64'b0011111111101011010110001000100111111110100100100001010000000101;
  assign mem[309] = 64'b1011111111100000100111101001000001110100000101111100010111100001;
  assign mem[310] = 64'b0011111111001110010101101100101000011110000100000001101000011011;
  assign mem[311] = 64'b1011111111101111000101101000111101010011111101110010000001011101;
  assign mem[312] = 64'b0011111111101110000100000000110011001010001010011000000010101100;
  assign mem[313] = 64'b1011111111010101111011100010011100110111100111101010011010010011;
  assign mem[314] = 64'b0011111111011011000000100000110101101100011111110100000000001001;
  assign mem[315] = 64'b1011111111101101000000101101010011111110101100101011110110010010;
  assign mem[316] = 64'b0011111111100111100101000000000001010111010011110101010111100101;
  assign mem[317] = 64'b1011111111100101101000101000110100101010010111010111001001010000;
  assign mem[318] = 64'b0011111110100101111111000000000011010010100100001100110101000011;
  assign mem[319] = 64'b1011111111101111111110000111000111011010110110111000000111011111;
  assign mem[320] = 64'b0011111111101111111111000010010100011101111100011101001111111000;
  assign mem[321] = 64'b1011111110011111011010010011011100110001110100011100111100000001;
  assign mem[322] = 64'b0011111111100101111011000011010010010101100000110111000001110100;
  assign mem[323] = 64'b1011111111100111010011111001010010001101101010001101001010001101;
  assign mem[324] = 64'b0011111111101101001011001011001000100000111000001110111110011111;
  assign mem[325] = 64'b1011111111011010010010110100000100100111110111101010000111100101;
  assign mem[326] = 64'b0011111111010110101010101001110101111101110001110111111000010111;
  assign mem[327] = 64'b1011111111101101111011010000010111110111110111100100011111011010;
  assign mem[328] = 64'b0011111111101111001011011100100111001001000010001001101010011101;
  assign mem[329] = 64'b1011111111001100110011111000110010110011000100101011001010000110;
  assign mem[330] = 64'b0011111111100000111101000010011010111011001010101000111001111110;
  assign mem[331] = 64'b1011111111101011001000111100110101000111000000000001001110110100;
  assign mem[332] = 64'b0011111111101010000011001001010111101010101110101111100100110111;
  assign mem[333] = 64'b1011111111100010100101100000011100100111011000101001110010101000;
  assign mem[334] = 64'b0011111111000101000110111101111110000101100101111100010111110010;
  assign mem[335] = 64'b1011111111101111100011111101010111111111101011100100000111011011;
  assign mem[336] = 64'b0011111111101111101111000001011000010111111001000100000110000110;
  assign mem[337] = 64'b1011111111000000011100101010000001000111101110101000001100011101;
  assign mem[338] = 64'b0011111111100011100010000100000110000101110111111110101100100010;
  assign mem[339] = 64'b1011111111101001010110001110111111100100100011100110110111010111;
  assign mem[340] = 64'b0011111111101011101111101101011111000100100100111000000011101010;
  assign mem[341] = 64'b1011111111011111111000101111011001001011111001110001001000010000;
  assign mem[342] = 64'b0011111111010000101100001101100111001111110110111101101110010000;
  assign mem[343] = 64'b1011111111101110111001001000001011100010010110101001110110111100;
  assign mem[344] = 64'b0011111111101110010100101001111100000100011100101001111111111100;
  assign mem[345] = 64'b1011111111010100011100101011100010100101010101110001000001010100;
  assign mem[346] = 64'b0011111111011100011011000111111101001001100101110000000000001011;
  assign mem[347] = 64'b1011111111101100101010111100000101101001101000001011100100000000;
  assign mem[348] = 64'b0011111111101000000110100001101100110011101101010111101011001100;
  assign mem[349] = 64'b1011111111100101000011001100000010011111010110011010000010011011;
  assign mem[350] = 64'b0011111110110001010001000000000100110100110101110000100110110011;
  assign mem[351] = 64'b1011111111101111111011010101100011101100101101100111001111000100;
  assign mem[352] = 64'b0011111111101111111001011111001110101111001011100011100101000000;
  assign mem[353] = 64'b1011111110110100011001100001000101111001001001110010000010010110;
  assign mem[354] = 64'b0011111111100100110000001010000101000101111011000000000000000100;
  assign mem[355] = 64'b1011111111101000010110111100010100011010111010010101100011001100;
  assign mem[356] = 64'b0011111111101100011111101000111001010010001000110011110011110011;
  assign mem[357] = 64'b1011111111011101001000000001011011101000111010011101101101011011;
  assign mem[358] = 64'b0011111111010011101100111100111011111010000001000001010010110111;
  assign mem[359] = 64'b1011111111101110011100100010011111011011011010101001011101000100;
  assign mem[360] = 64'b0011111111101110110010011011001011010011110000111011111110000100;
  assign mem[361] = 64'b1011111111010001011100101010000011010111011101100101000101110111;
  assign mem[362] = 64'b0011111111011111001101000000010110010110001111111101000001100111;
  assign mem[363] = 64'b1011111111101011111100000110010011100001010100110111011111011101;
  assign mem[364] = 64'b0011111111101001000110110001011001101111110101001001110110100010;
  assign mem[365] = 64'b1011111111100011110101111000001000111000110001011000001101000100;
  assign mem[366] = 64'b0011111110111101110001110000111011001011101011101001111111001001;
  assign mem[367] = 64'b1011111111101111110010000110010001101100111111101011011100100001;
  assign mem[368] = 64'b0011111111101111011111101010011000101001111001100011110101101110;
  assign mem[369] = 64'b1011111111000110101010000001001100000100111101100100101010110010;
  assign mem[370] = 64'b0011111111100010010000111101010111111011100110001010110000011111;
  assign mem[371] = 64'b1011111111101010010001100111100011001000000100011001101011001000;
  assign mem[372] = 64'b0011111111101010111011100000010010110100001111000001010001110100;
  assign mem[373] = 64'b1011111111100001010010010001010110101111001100110110110011101011;
  assign mem[374] = 64'b0011111111001011010001110011001011101111001111010110011100100010;
  assign mem[375] = 64'b1011111111101111010000111101000010000101111111111001001011011101;
  assign mem[376] = 64'b0011111111101101110010001101011111001011010000010000001001100000;
  assign mem[377] = 64'b1011111111010111011001100011010000001111001001000001100011110110;
  assign mem[378] = 64'b0011111111011001100100110111000101100001010000011011110111111111;
  assign mem[379] = 64'b1011111111101101010101010110111101010010111010010011111010110001;
  assign mem[380] = 64'b0011111111100111000010100100001010110011000101110110110101111010;
  assign mem[381] = 64'b1011111111100110001101010000001110100011000111000001101111101001;
  assign mem[382] = 64'b0011111110010010110110010011011010111011111000110000111011111101;
  assign mem[383] = 64'b1011111111101111111111101001110010110100010010110101000110100001;
  assign mem[384] = 64'b0011111111101111111111101001110010110100010010110101000110100001;
  assign mem[385] = 64'b1011111110010010110110010011011010111011111000110000111011111101;
  assign mem[386] = 64'b0011111111100110001101010000001110100011000111000001101111101001;
  assign mem[387] = 64'b1011111111100111000010100100001010110011000101110110110101111010;
  assign mem[388] = 64'b0011111111101101010101010110111101010010111010010011111010110001;
  assign mem[389] = 64'b1011111111011001100100110111000101100001010000011011110111111111;
  assign mem[390] = 64'b0011111111010111011001100011010000001111001001000001100011110110;
  assign mem[391] = 64'b1011111111101101110010001101011111001011010000010000001001100000;
  assign mem[392] = 64'b0011111111101111010000111101000010000101111111111001001011011101;
  assign mem[393] = 64'b1011111111001011010001110011001011101111001111010110011100100010;
  assign mem[394] = 64'b0011111111100001010010010001010110101111001100110110110011101011;
  assign mem[395] = 64'b1011111111101010111011100000010010110100001111000001010001110100;
  assign mem[396] = 64'b0011111111101010010001100111100011001000000100011001101011001000;
  assign mem[397] = 64'b1011111111100010010000111101010111111011100110001010110000011111;
  assign mem[398] = 64'b0011111111000110101010000001001100000100111101100100101010110010;
  assign mem[399] = 64'b1011111111101111011111101010011000101001111001100011110101101110;
  assign mem[400] = 64'b0011111111101111110010000110010001101100111111101011011100100001;
  assign mem[401] = 64'b1011111110111101110001110000111011001011101011101001111111001001;
  assign mem[402] = 64'b0011111111100011110101111000001000111000110001011000001101000100;
  assign mem[403] = 64'b1011111111101001000110110001011001101111110101001001110110100010;
  assign mem[404] = 64'b0011111111101011111100000110010011100001010100110111011111011101;
  assign mem[405] = 64'b1011111111011111001101000000010110010110001111111101000001100111;
  assign mem[406] = 64'b0011111111010001011100101010000011010111011101100101000101110111;
  assign mem[407] = 64'b1011111111101110110010011011001011010011110000111011111110000100;
  assign mem[408] = 64'b0011111111101110011100100010011111011011011010101001011101000100;
  assign mem[409] = 64'b1011111111010011101100111100111011111010000001000001010010110111;
  assign mem[410] = 64'b0011111111011101001000000001011011101000111010011101101101011011;
  assign mem[411] = 64'b1011111111101100011111101000111001010010001000110011110011110011;
  assign mem[412] = 64'b0011111111101000010110111100010100011010111010010101100011001100;
  assign mem[413] = 64'b1011111111100100110000001010000101000101111011000000000000000100;
  assign mem[414] = 64'b0011111110110100011001100001000101111001001001110010000010010110;
  assign mem[415] = 64'b1011111111101111111001011111001110101111001011100011100101000000;
  assign mem[416] = 64'b0011111111101111111011010101100011101100101101100111001111000100;
  assign mem[417] = 64'b1011111110110001010001000000000100110100110101110000100110110011;
  assign mem[418] = 64'b0011111111100101000011001100000010011111010110011010000010011011;
  assign mem[419] = 64'b1011111111101000000110100001101100110011101101010111101011001100;
  assign mem[420] = 64'b0011111111101100101010111100000101101001101000001011100100000000;
  assign mem[421] = 64'b1011111111011100011011000111111101001001100101110000000000001011;
  assign mem[422] = 64'b0011111111010100011100101011100010100101010101110001000001010100;
  assign mem[423] = 64'b1011111111101110010100101001111100000100011100101001111111111100;
  assign mem[424] = 64'b0011111111101110111001001000001011100010010110101001110110111100;
  assign mem[425] = 64'b1011111111010000101100001101100111001111110110111101101110010000;
  assign mem[426] = 64'b0011111111011111111000101111011001001011111001110001001000010000;
  assign mem[427] = 64'b1011111111101011101111101101011111000100100100111000000011101010;
  assign mem[428] = 64'b0011111111101001010110001110111111100100100011100110110111010111;
  assign mem[429] = 64'b1011111111100011100010000100000110000101110111111110101100100010;
  assign mem[430] = 64'b0011111111000000011100101010000001000111101110101000001100011101;
  assign mem[431] = 64'b1011111111101111101111000001011000010111111001000100000110000110;
  assign mem[432] = 64'b0011111111101111100011111101010111111111101011100100000111011011;
  assign mem[433] = 64'b1011111111000101000110111101111110000101100101111100010111110010;
  assign mem[434] = 64'b0011111111100010100101100000011100100111011000101001110010101000;
  assign mem[435] = 64'b1011111111101010000011001001010111101010101110101111100100110111;
  assign mem[436] = 64'b0011111111101011001000111100110101000111000000000001001110110100;
  assign mem[437] = 64'b1011111111100000111101000010011010111011001010101000111001111110;
  assign mem[438] = 64'b0011111111001100110011111000110010110011000100101011001010000110;
  assign mem[439] = 64'b1011111111101111001011011100100111001001000010001001101010011101;
  assign mem[440] = 64'b0011111111101101111011010000010111110111110111100100011111011010;
  assign mem[441] = 64'b1011111111010110101010101001110101111101110001110111111000010111;
  assign mem[442] = 64'b0011111111011010010010110100000100100111110111101010000111100101;
  assign mem[443] = 64'b1011111111101101001011001011001000100000111000001110111110011111;
  assign mem[444] = 64'b0011111111100111010011111001010010001101101010001101001010001101;
  assign mem[445] = 64'b1011111111100101111011000011010010010101100000110111000001110100;
  assign mem[446] = 64'b0011111110011111011010010011011100110001110100011100111100000001;
  assign mem[447] = 64'b1011111111101111111111000010010100011101111100011101001111111000;
  assign mem[448] = 64'b0011111111101111111110000111000111011010110110111000000111011111;
  assign mem[449] = 64'b1011111110100101111111000000000011010010100100001100110101000011;
  assign mem[450] = 64'b0011111111100101101000101000110100101010010111010111001001010000;
  assign mem[451] = 64'b1011111111100111100101000000000001010111010011110101010111100101;
  assign mem[452] = 64'b0011111111101101000000101101010011111110101100101011110110010010;
  assign mem[453] = 64'b1011111111011011000000100000110101101100011111110100000000001001;
  assign mem[454] = 64'b0011111111010101111011100010011100110111100111101010011010010011;
  assign mem[455] = 64'b1011111111101110000100000000110011001010001010011000000010101100;
  assign mem[456] = 64'b0011111111101111000101101000111101010011111101110010000001011101;
  assign mem[457] = 64'b1011111111001110010101101100101000011110000100000001101000011011;
  assign mem[458] = 64'b0011111111100000100111101001000001110100000101111100010111100001;
  assign mem[459] = 64'b1011111111101011010110001000100111111110100100100001010000000101;
  assign mem[460] = 64'b0011111111101001110100011011000111110101111010101000000011010101;
  assign mem[461] = 64'b1011111111100010111001111000000011100011111010001110101000010111;
  assign mem[462] = 64'b0011111111000011100011101101101110110000110011011000110100010100;
  assign mem[463] = 64'b1011111111101111100111111100111001010101101011011011001011001000;
  assign mem[464] = 64'b0011111111101111101011101000111010001110010001101100111110111011;
  assign mem[465] = 64'b1011111111000010000000010001011011010100111011000111101111001111;
  assign mem[466] = 64'b0011111111100011001110000100000000001101000011001000111001010111;
  assign mem[467] = 64'b1011111111101001100101011100111100101110110110000000110100100010;
  assign mem[468] = 64'b0011111111101011100011000011100011010010011101010000010011101001;
  assign mem[469] = 64'b1011111111100000010010000101011000100110101011100010001000011010;
  assign mem[470] = 64'b0011111111001111110111001101110000011010110111111110110111111001;
  assign mem[471] = 64'b1011111111101110111111100010001000001100000010111001010111101100;
  assign mem[472] = 64'b0011111111101110001100011110101011101000011100001100111000100101;
  assign mem[473] = 64'b1011111111010101001100001101100010000000101011110011110000100100;
  assign mem[474] = 64'b0011111111011011101101111100111100100011000001001011110100000001;
  assign mem[475] = 64'b1011111111101100110101111101100110001001100010110011001011110110;
  assign mem[476] = 64'b0011111111100111110101111000001101101100110000110011110110110010;
  assign mem[477] = 64'b1011111111100101010110000001000000111000100101110101000100110111;
  assign mem[478] = 64'b0011111110101100010000101000110100010010110000001101011111100011;
  assign mem[479] = 64'b1011111111101111111100111000001100001111100011010101011101011100;
  assign mem[480] = 64'b0011111111101111110111010101001110011111111100011111010001010110;
  assign mem[481] = 64'b1011111110110111100001110101100001101010010111010101101100100001;
  assign mem[482] = 64'b0011111111100100011100111011010100011011100110000111001101000111;
  assign mem[483] = 64'b1011111111101000100111000111111010011010010011011101010010101010;
  assign mem[484] = 64'b0011111111101100010100000100001000000001001010110110100100000111;
  assign mem[485] = 64'b1011111111011101110100101000111100010100100000011100110001011000;
  assign mem[486] = 64'b0011111111010010111101000010001011011010111011000000001110000111;
  assign mem[487] = 64'b1011111111101110100100001000010000110110000111011111011111110010;
  assign mem[488] = 64'b0011111111101110101011011011001011101000111001111010100010001110;
  assign mem[489] = 64'b1011111111010010001100111011101110101011110000111011101101110001;
  assign mem[490] = 64'b0011111111011110100000111110000011101010111110000101000100010100;
  assign mem[491] = 64'b1011111111101100001000001101111000111111101010010111000110110000;
  assign mem[492] = 64'b0011111111101000110111000100010100110011000101101001100011001100;
  assign mem[493] = 64'b1011111111100100001001011111111100010111100011100110101110110001;
  assign mem[494] = 64'b0011111110111010101001111011011100100100010010010101110000000011;
  assign mem[495] = 64'b1011111111101111110100110111100100010100001000100000101110000100;
  assign mem[496] = 64'b0011111111101111011011000011111101111101111101011011101110110111;
  assign mem[497] = 64'b1011111111001000001100110110011011101000100111000110010011000110;
  assign mem[498] = 64'b0011111111100001111100001111000010001011101111001000011000011011;
  assign mem[499] = 64'b1011111111101010011111110101100001010010100111111110011010011101;
  assign mem[500] = 64'b0011111111101010101101110011001001011001000101101100000011010100;
  assign mem[501] = 64'b1011111111100001100111010101101000001001111100101011100110111000;
  assign mem[502] = 64'b0011111111001001101111011100101111110010110111000100001101100110;
  assign mem[503] = 64'b1011111111101111010110001010001010110001011110001001111010000100;
  assign mem[504] = 64'b0011111111101101101000111000001110101001011001101000100110001000;
  assign mem[505] = 64'b1011111111011000001000001110001110110000010011101010101011000100;
  assign mem[506] = 64'b0011111111011000110110101010010100101110110010001010010010110000;
  assign mem[507] = 64'b1011111111101101011111010000101100000010101110001110110011111001;
  assign mem[508] = 64'b0011111111100110110001000000110101110011110000011000001001110101;
  assign mem[509] = 64'b1011111111100110011111001111011110000100100100011010111100010000;
  assign mem[510] = 64'b0011111101111001001000011111000011111110011001110000000001110001;
  assign mem[511] = 64'b1011111111101111111111111101100010000101100011101000101010010010;
  assign mem[512] = 64'b0011111111101111111111111111011000100001011000100001110100000010;
  assign mem[513] = 64'b1011111101101001001000011111100010111110110011001010010010111010;
  assign mem[514] = 64'b0011111111100110100011101101000111101010101000011001110001110001;
  assign mem[515] = 64'b1011111111100110101100100101110011101101001011111110001010011100;
  assign mem[516] = 64'b0011111111101101100001101100010010000100010001011010010001001111;
  assign mem[517] = 64'b1011111111011000101011000100101110000110110101011110110101000100;
  assign mem[518] = 64'b0011111111011000010011110110101010101010111100111001000000111111;
  assign mem[519] = 64'b1011111111101101100110100000000011011101100010110011110101000110;
  assign mem[520] = 64'b0011111111101111010111011010011011101101010000110110100001011101;
  assign mem[521] = 64'b1011111111001001010110110100100111101001101101100010101011111010;
  assign mem[522] = 64'b0011111111100001101100100101000000010111000100110111001110111111;
  assign mem[523] = 64'b1011111111101010101010010101010001111010001011001011100110001110;
  assign mem[524] = 64'b0011111111101010100011010110011101101110010101000101101011010010;
  assign mem[525] = 64'b1011111111100001110111000001101101100100110111000100100001110010;
  assign mem[526] = 64'b0011111111001000100101100001011100100111110001000001100000000100;
  assign mem[527] = 64'b1011111111101111011001110111010101010110100010000011110011101110;
  assign mem[528] = 64'b0011111111101111110101100000110100101101101001110101110010011110;
  assign mem[529] = 64'b1011111110111001110111111011011011101011001001001010100001011100;
  assign mem[530] = 64'b0011111111100100001110010111111101011011001010100100001110000000;
  assign mem[531] = 64'b1011111111101000110011000110101001110101000110000100011001010101;
  assign mem[532] = 64'b0011111111101100001011001101000101001001001100011110001111110001;
  assign mem[533] = 64'b1011111111011110010101111010100001101101001111001101100000100101;
  assign mem[534] = 64'b0011111111010010011000111110011010011001010101010101010010111010;
  assign mem[535] = 64'b1011111111101110101001101000001110010011111001100101100000000000;
  assign mem[536] = 64'b0011111111101110100101111110110000110110000000010110101100110000;
  assign mem[537] = 64'b1011111111010010110001000001101001001110100101010100010100100000;
  assign mem[538] = 64'b0011111111011101111111101111111101100110101010010100000111011110;
  assign mem[539] = 64'b1011111111101100010001001000001100110001010000011100000000000100;
  assign mem[540] = 64'b0011111111101000101011001000011100011110110111100001110110001000;
  assign mem[541] = 64'b1011111111100100011000000101101001101001001010110011001010100010;
  assign mem[542] = 64'b0011111110111000010011111000011100010010110000010011000010100001;
  assign mem[543] = 64'b1011111111101111110110101111101001110101000101000101001110001100;
  assign mem[544] = 64'b0011111111101111111101001101110001010100101100011011111011010011;
  assign mem[545] = 64'b1011111110101010101100010000000110111101010111111000001100010111;
  assign mem[546] = 64'b0011111111100101011010101100001101010001100101110110010010011111;
  assign mem[547] = 64'b1011111111100111110001101011100010011100111000101101001100110011;
  assign mem[548] = 64'b0011111111101100111000101011001100100111100110011010000001100000;
  assign mem[549] = 64'b1011111111011011100010100111100000010100111111010101011010010011;
  assign mem[550] = 64'b0011111111010101011000000100000000010010111101000110011110110100;
  assign mem[551] = 64'b1011111111101110001010011000111101000100001110010001100101111010;
  assign mem[552] = 64'b0011111111101111000001000101101000010100110011110111001110001100;
  assign mem[553] = 64'b1011111111001111011110110111010010000000101111010011100000000010;
  assign mem[554] = 64'b0011111111100000010111011111001111101100001100011011100010110111;
  assign mem[555] = 64'b1011111111101011011111110110011010000110111001111001001011101001;
  assign mem[556] = 64'b0011111111101001101001001101111110100100001010110000011010110010;
  assign mem[557] = 64'b1011111111100011001001000010000111101100010010011010011000011111;
  assign mem[558] = 64'b0011111111000010011001001001100101001101111111010011010000001001;
  assign mem[559] = 64'b1011111111101111101010101111101111001011000011001111110111011100;
  assign mem[560] = 64'b0011111111101111101000111001101110101100011110100001011110010001;
  assign mem[561] = 64'b1011111111000011001010110111101111111001010001010001011010100111;
  assign mem[562] = 64'b0011111111100010111110111100001001001011010001000001000000010101;
  assign mem[563] = 64'b1011111111101001110000101101000100010000111100000111010111000010;
  assign mem[564] = 64'b0011111111101011011001011000111100010100111111011011110001000111;
  assign mem[565] = 64'b1011111111100000100010010001000100100000001100101011000010001100;
  assign mem[566] = 64'b0011111111001110101110000110101101000110001011011110001101001000;
  assign mem[567] = 64'b1011111111101111000100001001000010111100100010011000111101011111;
  assign mem[568] = 64'b0011111111101110000110001010000000101111110111000110011011011001;
  assign mem[569] = 64'b1011111111010101101111101110011110001011100111011011001110110110;
  assign mem[570] = 64'b0011111111011011001011111001011100011101101100110001100101110010;
  assign mem[571] = 64'b1011111111101100111110000011000011101000110011100100011001111011;
  assign mem[572] = 64'b0011111111100111101001001111011100000111101111111001011111010010;
  assign mem[573] = 64'b1011111111100101100100000000000111010101111101110010001111011111;
  assign mem[574] = 64'b0011111110100111100011011011101010100101100001110100011010000110;
  assign mem[575] = 64'b1011111111101111111101110101001110111011000110111001000101100100;
  assign mem[576] = 64'b0011111111101111111111001110000010011100111000101010011001111001;
  assign mem[577] = 64'b1011111110011100010001010100111101001100111001010011101100011101;
  assign mem[578] = 64'b0011111111100101111111100111110010111101111001010110101000010000;
  assign mem[579] = 64'b1011111111100111001111100101010110001110000001111001100101000010;
  assign mem[580] = 64'b0011111111101101001101101111110001111011110010111111101111011100;
  assign mem[581] = 64'b1011111111011010000111010110010101000011101101010000101011000000;
  assign mem[582] = 64'b0011111111010110110110011001100001100011100010100000110010110110;
  assign mem[583] = 64'b1011111111101101111001000001011000001111011011011000110110000001;
  assign mem[584] = 64'b0011111111101111001100110110100001011010001110101010111011110000;
  assign mem[585] = 64'b1011111111001100011011011001000001010011010111010111010011011101;
  assign mem[586] = 64'b0011111111100001000010010111001001001000110100001010100101010111;
  assign mem[587] = 64'b1011111111101011000101100111010000101010010011001010001011110101;
  assign mem[588] = 64'b0011111111101010000110110010011011010010110000001010011101011110;
  assign mem[589] = 64'b1011111111100010100000011000101111101111010011010011110010111010;
  assign mem[590] = 64'b0011111111000101011111110000000010000110010101001100101111011110;
  assign mem[591] = 64'b1011111111101111100010111010011100110111110010110100101101111000;
  assign mem[592] = 64'b0011111111101111101111110100011100001111000010101000110110001000;
  assign mem[593] = 64'b1011111111000000000011101110100010101101011011111011100001011011;
  assign mem[594] = 64'b0011111111100011100111000010001111100011110101100011000000101001;
  assign mem[595] = 64'b1011111111101001010010011001000011100011101011000100101001101100;
  assign mem[596] = 64'b0011111111101011110010110101010011001011000011010010001100100111;
  assign mem[597] = 64'b1011111111011111101101110101011101011100001001001101001011011110;
  assign mem[598] = 64'b0011111111010000111000010101101101001110000101110100100111001110;
  assign mem[599] = 64'b1011111111101110110111011110101101101010000001111000011001010001;
  assign mem[600] = 64'b0011111111101110010110101001110101010101000001000110011111010011;
  assign mem[601] = 64'b1011111111010100010000110001000011011100100010010011011011110000;
  assign mem[602] = 64'b0011111111011100100110010111111111000011100001100101001110001001;
  assign mem[603] = 64'b1011111111101100101000001000111100011001101110011100010001001001;
  assign mem[604] = 64'b0011111111101000001010101001110000010011111101010100010111111111;
  assign mem[605] = 64'b1011111111100100111110011100110000100101110011001010010010000110;
  assign mem[606] = 64'b0011111110110010000011001001011001110100111011010100010001001101;
  assign mem[607] = 64'b1011111111101111111010111001110100100101001100000100000100001111;
  assign mem[608] = 64'b0011111111101111111001111110101010000101010010000010110101100000;
  assign mem[609] = 64'b1011111110110011100111011001111100010010110001011010001010011001;
  assign mem[610] = 64'b0011111111100100110100111011110001101101010110001001111101111111;
  assign mem[611] = 64'b1011111111101000010010110111000100010001101011111000001111111010;
  assign mem[612] = 64'b0011111111101100100010011111010110000111000000101001110000010011;
  assign mem[613] = 64'b1011111111011100111100110100101110101110111000011100110100100001;
  assign mem[614] = 64'b0011111111010011111000111001101111101001011011101100001001110001;
  assign mem[615] = 64'b1011111111101110011010100110000111000101010111010101001110100111;
  assign mem[616] = 64'b0011111111101110110100001000001101011110100110011001000000001001;
  assign mem[617] = 64'b1011111111010001010000100011111011101111110001101001001101111000;
  assign mem[618] = 64'b0011111111011111010111111101111011100110010101101100110110100011;
  assign mem[619] = 64'b1011111111101011111001000001101101100001000100010101010011000001;
  assign mem[620] = 64'b0011111111101001001010101010010000011111110001011010100000010101;
  assign mem[621] = 64'b1011111111100011110000111100010001001001100000011100010100011000;
  assign mem[622] = 64'b0011111110111110100011101011011111111101111001001010101000111111;
  assign mem[623] = 64'b1011111111101111110001010110111000111011011111011001101011110110;
  assign mem[624] = 64'b0011111111101111100000110000111101001010010000001100011000001100;
  assign mem[625] = 64'b1011111111000110010001010001101010000011000111011000001100001101;
  assign mem[626] = 64'b0011111111100010010110000111001101001100101110110111000100010000;
  assign mem[627] = 64'b1011111111101010001110000001100001001010010110010011101111000110;
  assign mem[628] = 64'b0011111111101010111110111000111111011000100111110101011110110110;
  assign mem[629] = 64'b1011111111100001001100111110100111001111111011100010010101001111;
  assign mem[630] = 64'b0011111111001011101010010110001100110100111100010101110110101101;
  assign mem[631] = 64'b1011111111101111001111100110101110111100000110111011110001100101;
  assign mem[632] = 64'b0011111111101101110100011111111011110011100010101001000101011010;
  assign mem[633] = 64'b1011111111010111001101110110001111001001001001100001000010010010;
  assign mem[634] = 64'b0011111111011001110000010111110101000100000011011111100111110010;
  assign mem[635] = 64'b1011111111101101010010110101101100011011000110000111010100100100;
  assign mem[636] = 64'b0011111111100111000110111010110010010110000011100100000110111111;
  assign mem[637] = 64'b1011111111100110001000101110010001001111111011000010001011111111;
  assign mem[638] = 64'b0011111110010101111111010100110100100001111110101011001000100110;
  assign mem[639] = 64'b1011111111101111111111100001110001101000011100001100101101110111;
  assign mem[640] = 64'b0011111111101111111111110000100101000011110001010011101111010001;
  assign mem[641] = 64'b1011111110001111011010100010100101101010101110011001011111001011;
  assign mem[642] = 64'b0011111111100110010001110001010101000011011111110101001101011011;
  assign mem[643] = 64'b1011111111100110111110001100101010011001110010010101101101110101;
  assign mem[644] = 64'b0011111111101101010111110111000101110010100010001000101001111111;
  assign mem[645] = 64'b1011111111011001011001010101010110110111101010111001010010001111;
  assign mem[646] = 64'b0011111111010111100101001111010111100110000100111101111110101110;
  assign mem[647] = 64'b1011111111101101101111111001111001000011100101010111010110011010;
  assign mem[648] = 64'b0011111111101111010010010010001000000110101111001010101110110100;
  assign mem[649] = 64'b1011111111001010111001001111000111010101111100111011100110101011;
  assign mem[650] = 64'b0011111111100001010111100011011011100100110110111110001010111100;
  assign mem[651] = 64'b1011111111101010111000000110100011110011010001011110110011101111;
  assign mem[652] = 64'b0011111111101010010101001100100100010000100100001111010100100011;
  assign mem[653] = 64'b1011111111100010001011110010110101100110001011000001001111100010;
  assign mem[654] = 64'b0011111111000111000010101111110110001101000010001100010011111111;
  assign mem[655] = 64'b1011111111101111011110100010100110011100000110100011001000101010;
  assign mem[656] = 64'b0011111111101111110010110100011100000011100100010100001101010100;
  assign mem[657] = 64'b1011111110111100111111110101001100111011001100000111110111000001;
  assign mem[658] = 64'b0011111111100011111010110011001111101010101111100000011010000000;
  assign mem[659] = 64'b1011111111101001000010110111100101000011010101110101111011111110;
  assign mem[660] = 64'b0011111111101011111111001001110100100101101000011011000101000111;
  assign mem[661] = 64'b1011111111011111000010000001100100000110101111111111011111111110;
  assign mem[662] = 64'b0011111111010001101000101111011111111011111010001111001001000011;
  assign mem[663] = 64'b1011111111101110110000101100111101001011000110101111011010110010;
  assign mem[664] = 64'b0011111111101110011110011101101100101001101001010001011001011010;
  assign mem[665] = 64'b1011111111010011100000111111010111100011010100111011011010101011;
  assign mem[666] = 64'b0011111111011101010011001101000000101011101010000110000010011101;
  assign mem[667] = 64'b1011111111101100011100110001010110001001100111101010101011010111;
  assign mem[668] = 64'b0011111111101000011011000000101000011101100110101010000110010101;
  assign mem[669] = 64'b1011111111100100101011010111100101010001011001110010001011110001;
  assign mem[670] = 64'b0011111110110101001011100111011101001010010011010100110100001010;
  assign mem[671] = 64'b1011111111101111111000111110100100101011111010011101100010000110;
  assign mem[672] = 64'b0011111111101111111011110000000100000010100000100110000110010001;
  assign mem[673] = 64'b1011111110110000011110110110000101001110010001100011000001100100;
  assign mem[674] = 64'b0011111111100101000111111010100000011100110110011001101010100110;
  assign mem[675] = 64'b1011111111101000000010011000101101110101011011100101001011111010;
  assign mem[676] = 64'b0011111111101100101101101110001000001010000000001101101010011001;
  assign mem[677] = 64'b1011111111011100001111110110110101000111001001100011000100101001;
  assign mem[678] = 64'b0011111111010100101000100101001111010001000110111000001011110011;
  assign mem[679] = 64'b1011111111101110010010101000110111111111100000011100111001011110;
  assign mem[680] = 64'b0011111111101110111010110000011101001100010100001010010101000100;
  assign mem[681] = 64'b1011111111010000100000000100111000000101111010110110011000011110;
  assign mem[682] = 64'b0011111111100000000001110100000011001000001010111000001011100001;
  assign mem[683] = 64'b1011111111101011101100100100100110100000101101101100010000001101;
  assign mem[684] = 64'b0011111111101001011010000011111101000010101111010111111111100001;
  assign mem[685] = 64'b1011111111100011011101000101001100011011100000010111111110001101;
  assign mem[686] = 64'b0011111111000000110101100100110110111100101100100110011110000110;
  assign mem[687] = 64'b1011111111101111101110001101000110001101011001101010110110110111;
  assign mem[688] = 64'b0011111111101111100100111111000101001111100001011010110000001000;
  assign mem[689] = 64'b1011111111000100101110001011000101111111011110011111101010001000;
  assign mem[690] = 64'b0011111111100010101010100111011011101000011110101110101101011000;
  assign mem[691] = 64'b1011111111101001111111011111010011110001001100010100100111011110;
  assign mem[692] = 64'b0011111111101011001100010001010110100101111100110111101111110011;
  assign mem[693] = 64'b1011111111100000110111101101000010111000010010111100010010110110;
  assign mem[694] = 64'b0011111111001101001100010111011101001101001011001011110111101110;
  assign mem[695] = 64'b1011111111101111001010000001011111111100010001100000100111001110;
  assign mem[696] = 64'b0011111111101101111101011110001101101010100110111010010110011100;
  assign mem[697] = 64'b1011111111010110011110111001010010011100101011010110001111001011;
  assign mem[698] = 64'b0011111111011010011110010000110011010011110110111111001100011011;
  assign mem[699] = 64'b1011111111101101001000100101010111000110111001011010010011100001;
  assign mem[700] = 64'b0011111111100111011000001100010100101100001100000100011101100100;
  assign mem[701] = 64'b1011111111100101110110011101111011100111001111100011010001011100;
  assign mem[702] = 64'b0011111110100001010001101000010111011011010000101100000101111111;
  assign mem[703] = 64'b1011111111101111111110110101010111100100001001011111110110101110;
  assign mem[704] = 64'b0011111111101111111110010111110001000010000010001100000000010100;
  assign mem[705] = 64'b1011111110100100011010100011100101101111111110000110000101111001;
  assign mem[706] = 64'b0011111111100101101101010000101100100110010011110111010001001000;
  assign mem[707] = 64'b1011111111100111100000101111101100011011100100001011001101011011;
  assign mem[708] = 64'b0011111111101101000011010110011100101111010110011101001010111001;
  assign mem[709] = 64'b1011111111011010110101000111001100010010010111001101110000001001;
  assign mem[710] = 64'b0011111111010110000111010101100101011100100010001100001000000010;
  assign mem[711] = 64'b1011111111101110000001110110011011011001001010000000111101010100;
  assign mem[712] = 64'b0011111111101111000111000111101010111110001010000100011100001000;
  assign mem[713] = 64'b1011111111001101111101010001011000111111000000010000100110011010;
  assign mem[714] = 64'b0011111111100000101101000000010110000111100011111000010111101100;
  assign mem[715] = 64'b1011111111101011010010110111010000001001110111100111100100100101;
  assign mem[716] = 64'b0011111111101001111000001000001011101101101101000010010001110010;
  assign mem[717] = 64'b1011111111100010110100110011001111010011010011101001101110111000;
  assign mem[718] = 64'b0011111111000011111100100010111101010111110110110100100010010011;
  assign mem[719] = 64'b1011111111101111100110111110110101111100111110111101111000101001;
  assign mem[720] = 64'b0011111111101111101100100000110111000110100000011101010101001101;
  assign mem[721] = 64'b1011111111000001100111011000100101000000101111100010010011100111;
  assign mem[722] = 64'b0011111111100011010011000101001001010010110000010100110111100001;
  assign mem[723] = 64'b1011111111101001100001101010111011110001010001010111010110010100;
  assign mem[724] = 64'b0011111111101011100110001111101000011111110110010001010101011110;
  assign mem[725] = 64'b1011111111100000001100101010111001010101111011011011110110010110;
  assign mem[726] = 64'b0011111111010000000111110001100000000110101110011111110111010010;
  assign mem[727] = 64'b1011111111101110111101111101011011100101000111001010001111000000;
  assign mem[728] = 64'b0011111111101110001110100011001111101100011101011100111010000101;
  assign mem[729] = 64'b1011111111010101000000010110001111011100000110010111000001001000;
  assign mem[730] = 64'b0011111111011011111001010001010100010111111111111100000011011001;
  assign mem[731] = 64'b1011111111101100110011001110111000100000110000101101111010100000;
  assign mem[732] = 64'b0011111111100111111010000011111110000111101100000011011010000110;
  assign mem[733] = 64'b1011111111100101010001010100111111110101000101011001110111111100;
  assign mem[734] = 64'b0011111110101101110101000000011011111001100000001000111011001001;
  assign mem[735] = 64'b1011111111101111111100100001011000010100111000010011000111101101;
  assign mem[736] = 64'b0011111111101111110111111001100100100010111101110011001100000111;
  assign mem[737] = 64'b1011111110110110101111110001101100111110011110011011000100101001;
  assign mem[738] = 64'b0011111111100100100001110000001100110000011000001001000111111111;
  assign mem[739] = 64'b1011111111101000100011000110011011100111010010000001101110100001;
  assign mem[740] = 64'b0011111111101100010110111110111101011001111111101111100001011010;
  assign mem[741] = 64'b1011111111011101101001100000110001011100111110100001000011011001;
  assign mem[742] = 64'b0011111111010011001001000001111110110110001110001011101010101111;
  assign mem[743] = 64'b1011111111101110100010010000100101011011101011010110000000100101;
  assign mem[744] = 64'b0011111111101110101101001100111101010001010110111000100000010001;
  assign mem[745] = 64'b1011111111010010000000111000010110000011110101110010011110111110;
  assign mem[746] = 64'b0011111111011110101100000000011010010101111100100101011000100000;
  assign mem[747] = 64'b1011111111101100000101001101100111011100010001100101111001010111;
  assign mem[748] = 64'b0011111111101000111011000001000010011011010010000110110001001001;
  assign mem[749] = 64'b1011111111100100000100100111001001100110001111010001000010001100;
  assign mem[750] = 64'b0011111110111011011011111010011011101100001110001111011001001100;
  assign mem[751] = 64'b1011111111101111110100001101000101011000110110000110000010000111;
  assign mem[752] = 64'b0011111111101111011100001111011001000011010010110111111010110111;
  assign mem[753] = 64'b1011111111000111110100001010011110111011110100101100101100011100;
  assign mem[754] = 64'b0011111111100010000001011011101010100001011101010110000011010110;
  assign mem[755] = 64'b1011111111101010011100010011100011011110100111010110000011110101;
  assign mem[756] = 64'b0011111111101010110001001111111110111101001111101111101011001000;
  assign mem[757] = 64'b1011111111100001100010000101100100011111001110100100011011100101;
  assign mem[758] = 64'b0011111111001010001000000011111000011011000110000011000111011010;
  assign mem[759] = 64'b1011111111101111010100111000101100011111101011110010110100000111;
  assign mem[760] = 64'b0011111111101101101011001111010000101100111001101000101010111001;
  assign mem[761] = 64'b1011111111010111111100100100110111010011011100110100000111100100;
  assign mem[762] = 64'b0011111111011001000010001110111110000001111011110111101111010001;
  assign mem[763] = 64'b1011111111101101011100110011111101010000100011000000110111111111;
  assign mem[764] = 64'b0011111111100110110101011010111111101111010010101010111111001101;
  assign mem[765] = 64'b1011111111100110011010110000111100111111010100101011001110000110;
  assign mem[766] = 64'b0011111110000010110110010110101100001110010100001001011100000011;
  assign mem[767] = 64'b1011111111101111111111111010011100101100100101111000110001001111;
  assign mem[768] = 64'b0011111111101111111111111010011100101100100101111000110001001111;
  assign mem[769] = 64'b1011111110000010110110010110101100001110010100001001011100000011;
  assign mem[770] = 64'b0011111111100110011010110000111100111111010100101011001110000110;
  assign mem[771] = 64'b1011111111100110110101011010111111101111010010101010111111001101;
  assign mem[772] = 64'b0011111111101101011100110011111101010000100011000000110111111111;
  assign mem[773] = 64'b1011111111011001000010001110111110000001111011110111101111010001;
  assign mem[774] = 64'b0011111111010111111100100100110111010011011100110100000111100100;
  assign mem[775] = 64'b1011111111101101101011001111010000101100111001101000101010111001;
  assign mem[776] = 64'b0011111111101111010100111000101100011111101011110010110100000111;
  assign mem[777] = 64'b1011111111001010001000000011111000011011000110000011000111011010;
  assign mem[778] = 64'b0011111111100001100010000101100100011111001110100100011011100101;
  assign mem[779] = 64'b1011111111101010110001001111111110111101001111101111101011001000;
  assign mem[780] = 64'b0011111111101010011100010011100011011110100111010110000011110101;
  assign mem[781] = 64'b1011111111100010000001011011101010100001011101010110000011010110;
  assign mem[782] = 64'b0011111111000111110100001010011110111011110100101100101100011100;
  assign mem[783] = 64'b1011111111101111011100001111011001000011010010110111111010110111;
  assign mem[784] = 64'b0011111111101111110100001101000101011000110110000110000010000111;
  assign mem[785] = 64'b1011111110111011011011111010011011101100001110001111011001001100;
  assign mem[786] = 64'b0011111111100100000100100111001001100110001111010001000010001100;
  assign mem[787] = 64'b1011111111101000111011000001000010011011010010000110110001001001;
  assign mem[788] = 64'b0011111111101100000101001101100111011100010001100101111001010111;
  assign mem[789] = 64'b1011111111011110101100000000011010010101111100100101011000100000;
  assign mem[790] = 64'b0011111111010010000000111000010110000011110101110010011110111110;
  assign mem[791] = 64'b1011111111101110101101001100111101010001010110111000100000010001;
  assign mem[792] = 64'b0011111111101110100010010000100101011011101011010110000000100101;
  assign mem[793] = 64'b1011111111010011001001000001111110110110001110001011101010101111;
  assign mem[794] = 64'b0011111111011101101001100000110001011100111110100001000011011001;
  assign mem[795] = 64'b1011111111101100010110111110111101011001111111101111100001011010;
  assign mem[796] = 64'b0011111111101000100011000110011011100111010010000001101110100001;
  assign mem[797] = 64'b1011111111100100100001110000001100110000011000001001000111111111;
  assign mem[798] = 64'b0011111110110110101111110001101100111110011110011011000100101001;
  assign mem[799] = 64'b1011111111101111110111111001100100100010111101110011001100000111;
  assign mem[800] = 64'b0011111111101111111100100001011000010100111000010011000111101101;
  assign mem[801] = 64'b1011111110101101110101000000011011111001100000001000111011001001;
  assign mem[802] = 64'b0011111111100101010001010100111111110101000101011001110111111100;
  assign mem[803] = 64'b1011111111100111111010000011111110000111101100000011011010000110;
  assign mem[804] = 64'b0011111111101100110011001110111000100000110000101101111010100000;
  assign mem[805] = 64'b1011111111011011111001010001010100010111111111111100000011011001;
  assign mem[806] = 64'b0011111111010101000000010110001111011100000110010111000001001000;
  assign mem[807] = 64'b1011111111101110001110100011001111101100011101011100111010000101;
  assign mem[808] = 64'b0011111111101110111101111101011011100101000111001010001111000000;
  assign mem[809] = 64'b1011111111010000000111110001100000000110101110011111110111010010;
  assign mem[810] = 64'b0011111111100000001100101010111001010101111011011011110110010110;
  assign mem[811] = 64'b1011111111101011100110001111101000011111110110010001010101011110;
  assign mem[812] = 64'b0011111111101001100001101010111011110001010001010111010110010100;
  assign mem[813] = 64'b1011111111100011010011000101001001010010110000010100110111100001;
  assign mem[814] = 64'b0011111111000001100111011000100101000000101111100010010011100111;
  assign mem[815] = 64'b1011111111101111101100100000110111000110100000011101010101001101;
  assign mem[816] = 64'b0011111111101111100110111110110101111100111110111101111000101001;
  assign mem[817] = 64'b1011111111000011111100100010111101010111110110110100100010010011;
  assign mem[818] = 64'b0011111111100010110100110011001111010011010011101001101110111000;
  assign mem[819] = 64'b1011111111101001111000001000001011101101101101000010010001110010;
  assign mem[820] = 64'b0011111111101011010010110111010000001001110111100111100100100101;
  assign mem[821] = 64'b1011111111100000101101000000010110000111100011111000010111101100;
  assign mem[822] = 64'b0011111111001101111101010001011000111111000000010000100110011010;
  assign mem[823] = 64'b1011111111101111000111000111101010111110001010000100011100001000;
  assign mem[824] = 64'b0011111111101110000001110110011011011001001010000000111101010100;
  assign mem[825] = 64'b1011111111010110000111010101100101011100100010001100001000000010;
  assign mem[826] = 64'b0011111111011010110101000111001100010010010111001101110000001001;
  assign mem[827] = 64'b1011111111101101000011010110011100101111010110011101001010111001;
  assign mem[828] = 64'b0011111111100111100000101111101100011011100100001011001101011011;
  assign mem[829] = 64'b1011111111100101101101010000101100100110010011110111010001001000;
  assign mem[830] = 64'b0011111110100100011010100011100101101111111110000110000101111001;
  assign mem[831] = 64'b1011111111101111111110010111110001000010000010001100000000010100;
  assign mem[832] = 64'b0011111111101111111110110101010111100100001001011111110110101110;
  assign mem[833] = 64'b1011111110100001010001101000010111011011010000101100000101111111;
  assign mem[834] = 64'b0011111111100101110110011101111011100111001111100011010001011100;
  assign mem[835] = 64'b1011111111100111011000001100010100101100001100000100011101100100;
  assign mem[836] = 64'b0011111111101101001000100101010111000110111001011010010011100001;
  assign mem[837] = 64'b1011111111011010011110010000110011010011110110111111001100011011;
  assign mem[838] = 64'b0011111111010110011110111001010010011100101011010110001111001011;
  assign mem[839] = 64'b1011111111101101111101011110001101101010100110111010010110011100;
  assign mem[840] = 64'b0011111111101111001010000001011111111100010001100000100111001110;
  assign mem[841] = 64'b1011111111001101001100010111011101001101001011001011110111101110;
  assign mem[842] = 64'b0011111111100000110111101101000010111000010010111100010010110110;
  assign mem[843] = 64'b1011111111101011001100010001010110100101111100110111101111110011;
  assign mem[844] = 64'b0011111111101001111111011111010011110001001100010100100111011110;
  assign mem[845] = 64'b1011111111100010101010100111011011101000011110101110101101011000;
  assign mem[846] = 64'b0011111111000100101110001011000101111111011110011111101010001000;
  assign mem[847] = 64'b1011111111101111100100111111000101001111100001011010110000001000;
  assign mem[848] = 64'b0011111111101111101110001101000110001101011001101010110110110111;
  assign mem[849] = 64'b1011111111000000110101100100110110111100101100100110011110000110;
  assign mem[850] = 64'b0011111111100011011101000101001100011011100000010111111110001101;
  assign mem[851] = 64'b1011111111101001011010000011111101000010101111010111111111100001;
  assign mem[852] = 64'b0011111111101011101100100100100110100000101101101100010000001101;
  assign mem[853] = 64'b1011111111100000000001110100000011001000001010111000001011100001;
  assign mem[854] = 64'b0011111111010000100000000100111000000101111010110110011000011110;
  assign mem[855] = 64'b1011111111101110111010110000011101001100010100001010010101000100;
  assign mem[856] = 64'b0011111111101110010010101000110111111111100000011100111001011110;
  assign mem[857] = 64'b1011111111010100101000100101001111010001000110111000001011110011;
  assign mem[858] = 64'b0011111111011100001111110110110101000111001001100011000100101001;
  assign mem[859] = 64'b1011111111101100101101101110001000001010000000001101101010011001;
  assign mem[860] = 64'b0011111111101000000010011000101101110101011011100101001011111010;
  assign mem[861] = 64'b1011111111100101000111111010100000011100110110011001101010100110;
  assign mem[862] = 64'b0011111110110000011110110110000101001110010001100011000001100100;
  assign mem[863] = 64'b1011111111101111111011110000000100000010100000100110000110010001;
  assign mem[864] = 64'b0011111111101111111000111110100100101011111010011101100010000110;
  assign mem[865] = 64'b1011111110110101001011100111011101001010010011010100110100001010;
  assign mem[866] = 64'b0011111111100100101011010111100101010001011001110010001011110001;
  assign mem[867] = 64'b1011111111101000011011000000101000011101100110101010000110010101;
  assign mem[868] = 64'b0011111111101100011100110001010110001001100111101010101011010111;
  assign mem[869] = 64'b1011111111011101010011001101000000101011101010000110000010011101;
  assign mem[870] = 64'b0011111111010011100000111111010111100011010100111011011010101011;
  assign mem[871] = 64'b1011111111101110011110011101101100101001101001010001011001011010;
  assign mem[872] = 64'b0011111111101110110000101100111101001011000110101111011010110010;
  assign mem[873] = 64'b1011111111010001101000101111011111111011111010001111001001000011;
  assign mem[874] = 64'b0011111111011111000010000001100100000110101111111111011111111110;
  assign mem[875] = 64'b1011111111101011111111001001110100100101101000011011000101000111;
  assign mem[876] = 64'b0011111111101001000010110111100101000011010101110101111011111110;
  assign mem[877] = 64'b1011111111100011111010110011001111101010101111100000011010000000;
  assign mem[878] = 64'b0011111110111100111111110101001100111011001100000111110111000001;
  assign mem[879] = 64'b1011111111101111110010110100011100000011100100010100001101010100;
  assign mem[880] = 64'b0011111111101111011110100010100110011100000110100011001000101010;
  assign mem[881] = 64'b1011111111000111000010101111110110001101000010001100010011111111;
  assign mem[882] = 64'b0011111111100010001011110010110101100110001011000001001111100010;
  assign mem[883] = 64'b1011111111101010010101001100100100010000100100001111010100100011;
  assign mem[884] = 64'b0011111111101010111000000110100011110011010001011110110011101111;
  assign mem[885] = 64'b1011111111100001010111100011011011100100110110111110001010111100;
  assign mem[886] = 64'b0011111111001010111001001111000111010101111100111011100110101011;
  assign mem[887] = 64'b1011111111101111010010010010001000000110101111001010101110110100;
  assign mem[888] = 64'b0011111111101101101111111001111001000011100101010111010110011010;
  assign mem[889] = 64'b1011111111010111100101001111010111100110000100111101111110101110;
  assign mem[890] = 64'b0011111111011001011001010101010110110111101010111001010010001111;
  assign mem[891] = 64'b1011111111101101010111110111000101110010100010001000101001111111;
  assign mem[892] = 64'b0011111111100110111110001100101010011001110010010101101101110101;
  assign mem[893] = 64'b1011111111100110010001110001010101000011011111110101001101011011;
  assign mem[894] = 64'b0011111110001111011010100010100101101010101110011001011111001011;
  assign mem[895] = 64'b1011111111101111111111110000100101000011110001010011101111010001;
  assign mem[896] = 64'b0011111111101111111111100001110001101000011100001100101101110111;
  assign mem[897] = 64'b1011111110010101111111010100110100100001111110101011001000100110;
  assign mem[898] = 64'b0011111111100110001000101110010001001111111011000010001011111111;
  assign mem[899] = 64'b1011111111100111000110111010110010010110000011100100000110111111;
  assign mem[900] = 64'b0011111111101101010010110101101100011011000110000111010100100100;
  assign mem[901] = 64'b1011111111011001110000010111110101000100000011011111100111110010;
  assign mem[902] = 64'b0011111111010111001101110110001111001001001001100001000010010010;
  assign mem[903] = 64'b1011111111101101110100011111111011110011100010101001000101011010;
  assign mem[904] = 64'b0011111111101111001111100110101110111100000110111011110001100101;
  assign mem[905] = 64'b1011111111001011101010010110001100110100111100010101110110101101;
  assign mem[906] = 64'b0011111111100001001100111110100111001111111011100010010101001111;
  assign mem[907] = 64'b1011111111101010111110111000111111011000100111110101011110110110;
  assign mem[908] = 64'b0011111111101010001110000001100001001010010110010011101111000110;
  assign mem[909] = 64'b1011111111100010010110000111001101001100101110110111000100010000;
  assign mem[910] = 64'b0011111111000110010001010001101010000011000111011000001100001101;
  assign mem[911] = 64'b1011111111101111100000110000111101001010010000001100011000001100;
  assign mem[912] = 64'b0011111111101111110001010110111000111011011111011001101011110110;
  assign mem[913] = 64'b1011111110111110100011101011011111111101111001001010101000111111;
  assign mem[914] = 64'b0011111111100011110000111100010001001001100000011100010100011000;
  assign mem[915] = 64'b1011111111101001001010101010010000011111110001011010100000010101;
  assign mem[916] = 64'b0011111111101011111001000001101101100001000100010101010011000001;
  assign mem[917] = 64'b1011111111011111010111111101111011100110010101101100110110100011;
  assign mem[918] = 64'b0011111111010001010000100011111011101111110001101001001101111000;
  assign mem[919] = 64'b1011111111101110110100001000001101011110100110011001000000001001;
  assign mem[920] = 64'b0011111111101110011010100110000111000101010111010101001110100111;
  assign mem[921] = 64'b1011111111010011111000111001101111101001011011101100001001110001;
  assign mem[922] = 64'b0011111111011100111100110100101110101110111000011100110100100001;
  assign mem[923] = 64'b1011111111101100100010011111010110000111000000101001110000010011;
  assign mem[924] = 64'b0011111111101000010010110111000100010001101011111000001111111010;
  assign mem[925] = 64'b1011111111100100110100111011110001101101010110001001111101111111;
  assign mem[926] = 64'b0011111110110011100111011001111100010010110001011010001010011001;
  assign mem[927] = 64'b1011111111101111111001111110101010000101010010000010110101100000;
  assign mem[928] = 64'b0011111111101111111010111001110100100101001100000100000100001111;
  assign mem[929] = 64'b1011111110110010000011001001011001110100111011010100010001001101;
  assign mem[930] = 64'b0011111111100100111110011100110000100101110011001010010010000110;
  assign mem[931] = 64'b1011111111101000001010101001110000010011111101010100010111111111;
  assign mem[932] = 64'b0011111111101100101000001000111100011001101110011100010001001001;
  assign mem[933] = 64'b1011111111011100100110010111111111000011100001100101001110001001;
  assign mem[934] = 64'b0011111111010100010000110001000011011100100010010011011011110000;
  assign mem[935] = 64'b1011111111101110010110101001110101010101000001000110011111010011;
  assign mem[936] = 64'b0011111111101110110111011110101101101010000001111000011001010001;
  assign mem[937] = 64'b1011111111010000111000010101101101001110000101110100100111001110;
  assign mem[938] = 64'b0011111111011111101101110101011101011100001001001101001011011110;
  assign mem[939] = 64'b1011111111101011110010110101010011001011000011010010001100100111;
  assign mem[940] = 64'b0011111111101001010010011001000011100011101011000100101001101100;
  assign mem[941] = 64'b1011111111100011100111000010001111100011110101100011000000101001;
  assign mem[942] = 64'b0011111111000000000011101110100010101101011011111011100001011011;
  assign mem[943] = 64'b1011111111101111101111110100011100001111000010101000110110001000;
  assign mem[944] = 64'b0011111111101111100010111010011100110111110010110100101101111000;
  assign mem[945] = 64'b1011111111000101011111110000000010000110010101001100101111011110;
  assign mem[946] = 64'b0011111111100010100000011000101111101111010011010011110010111010;
  assign mem[947] = 64'b1011111111101010000110110010011011010010110000001010011101011110;
  assign mem[948] = 64'b0011111111101011000101100111010000101010010011001010001011110101;
  assign mem[949] = 64'b1011111111100001000010010111001001001000110100001010100101010111;
  assign mem[950] = 64'b0011111111001100011011011001000001010011010111010111010011011101;
  assign mem[951] = 64'b1011111111101111001100110110100001011010001110101010111011110000;
  assign mem[952] = 64'b0011111111101101111001000001011000001111011011011000110110000001;
  assign mem[953] = 64'b1011111111010110110110011001100001100011100010100000110010110110;
  assign mem[954] = 64'b0011111111011010000111010110010101000011101101010000101011000000;
  assign mem[955] = 64'b1011111111101101001101101111110001111011110010111111101111011100;
  assign mem[956] = 64'b0011111111100111001111100101010110001110000001111001100101000010;
  assign mem[957] = 64'b1011111111100101111111100111110010111101111001010110101000010000;
  assign mem[958] = 64'b0011111110011100010001010100111101001100111001010011101100011101;
  assign mem[959] = 64'b1011111111101111111111001110000010011100111000101010011001111001;
  assign mem[960] = 64'b0011111111101111111101110101001110111011000110111001000101100100;
  assign mem[961] = 64'b1011111110100111100011011011101010100101100001110100011010000110;
  assign mem[962] = 64'b0011111111100101100100000000000111010101111101110010001111011111;
  assign mem[963] = 64'b1011111111100111101001001111011100000111101111111001011111010010;
  assign mem[964] = 64'b0011111111101100111110000011000011101000110011100100011001111011;
  assign mem[965] = 64'b1011111111011011001011111001011100011101101100110001100101110010;
  assign mem[966] = 64'b0011111111010101101111101110011110001011100111011011001110110110;
  assign mem[967] = 64'b1011111111101110000110001010000000101111110111000110011011011001;
  assign mem[968] = 64'b0011111111101111000100001001000010111100100010011000111101011111;
  assign mem[969] = 64'b1011111111001110101110000110101101000110001011011110001101001000;
  assign mem[970] = 64'b0011111111100000100010010001000100100000001100101011000010001100;
  assign mem[971] = 64'b1011111111101011011001011000111100010100111111011011110001000111;
  assign mem[972] = 64'b0011111111101001110000101101000100010000111100000111010111000010;
  assign mem[973] = 64'b1011111111100010111110111100001001001011010001000001000000010101;
  assign mem[974] = 64'b0011111111000011001010110111101111111001010001010001011010100111;
  assign mem[975] = 64'b1011111111101111101000111001101110101100011110100001011110010001;
  assign mem[976] = 64'b0011111111101111101010101111101111001011000011001111110111011100;
  assign mem[977] = 64'b1011111111000010011001001001100101001101111111010011010000001001;
  assign mem[978] = 64'b0011111111100011001001000010000111101100010010011010011000011111;
  assign mem[979] = 64'b1011111111101001101001001101111110100100001010110000011010110010;
  assign mem[980] = 64'b0011111111101011011111110110011010000110111001111001001011101001;
  assign mem[981] = 64'b1011111111100000010111011111001111101100001100011011100010110111;
  assign mem[982] = 64'b0011111111001111011110110111010010000000101111010011100000000010;
  assign mem[983] = 64'b1011111111101111000001000101101000010100110011110111001110001100;
  assign mem[984] = 64'b0011111111101110001010011000111101000100001110010001100101111010;
  assign mem[985] = 64'b1011111111010101011000000100000000010010111101000110011110110100;
  assign mem[986] = 64'b0011111111011011100010100111100000010100111111010101011010010011;
  assign mem[987] = 64'b1011111111101100111000101011001100100111100110011010000001100000;
  assign mem[988] = 64'b0011111111100111110001101011100010011100111000101101001100110011;
  assign mem[989] = 64'b1011111111100101011010101100001101010001100101110110010010011111;
  assign mem[990] = 64'b0011111110101010101100010000000110111101010111111000001100010111;
  assign mem[991] = 64'b1011111111101111111101001101110001010100101100011011111011010011;
  assign mem[992] = 64'b0011111111101111110110101111101001110101000101000101001110001100;
  assign mem[993] = 64'b1011111110111000010011111000011100010010110000010011000010100001;
  assign mem[994] = 64'b0011111111100100011000000101101001101001001010110011001010100010;
  assign mem[995] = 64'b1011111111101000101011001000011100011110110111100001110110001000;
  assign mem[996] = 64'b0011111111101100010001001000001100110001010000011100000000000100;
  assign mem[997] = 64'b1011111111011101111111101111111101100110101010010100000111011110;
  assign mem[998] = 64'b0011111111010010110001000001101001001110100101010100010100100000;
  assign mem[999] = 64'b1011111111101110100101111110110000110110000000010110101100110000;
  assign mem[1000] = 64'b0011111111101110101001101000001110010011111001100101100000000000;
  assign mem[1001] = 64'b1011111111010010011000111110011010011001010101010101010010111010;
  assign mem[1002] = 64'b0011111111011110010101111010100001101101001111001101100000100101;
  assign mem[1003] = 64'b1011111111101100001011001101000101001001001100011110001111110001;
  assign mem[1004] = 64'b0011111111101000110011000110101001110101000110000100011001010101;
  assign mem[1005] = 64'b1011111111100100001110010111111101011011001010100100001110000000;
  assign mem[1006] = 64'b0011111110111001110111111011011011101011001001001010100001011100;
  assign mem[1007] = 64'b1011111111101111110101100000110100101101101001110101110010011110;
  assign mem[1008] = 64'b0011111111101111011001110111010101010110100010000011110011101110;
  assign mem[1009] = 64'b1011111111001000100101100001011100100111110001000001100000000100;
  assign mem[1010] = 64'b0011111111100001110111000001101101100100110111000100100001110010;
  assign mem[1011] = 64'b1011111111101010100011010110011101101110010101000101101011010010;
  assign mem[1012] = 64'b0011111111101010101010010101010001111010001011001011100110001110;
  assign mem[1013] = 64'b1011111111100001101100100101000000010111000100110111001110111111;
  assign mem[1014] = 64'b0011111111001001010110110100100111101001101101100010101011111010;
  assign mem[1015] = 64'b1011111111101111010111011010011011101101010000110110100001011101;
  assign mem[1016] = 64'b0011111111101101100110100000000011011101100010110011110101000110;
  assign mem[1017] = 64'b1011111111011000010011110110101010101010111100111001000000111111;
  assign mem[1018] = 64'b0011111111011000101011000100101110000110110101011110110101000100;
  assign mem[1019] = 64'b1011111111101101100001101100010010000100010001011010010001001111;
  assign mem[1020] = 64'b0011111111100110101100100101110011101101001011111110001010011100;
  assign mem[1021] = 64'b1011111111100110100011101101000111101010101000011001110001110001;
  assign mem[1022] = 64'b0011111101101001001000011111100010111110110011001010010010111010;
  assign mem[1023] = 64'b1011111111101111111111111111011000100001011000100001110100000010;
  always@(*)
  begin
    data_out_t <= mem[addr_f];
  end
  wire [63:0] data_out_reg [n_outreg:0];
  generate if (n_outreg > 0)
  begin
    for( i=n_outreg-1; i >= 1; i=i-1)
    begin: data_out_reg_stage
      mgc_generic_reg #(
        .width(64),
        .ph_clk(1),
        .ph_en(0),
        .ph_a_rst(0),
        .ph_s_rst(0),
        .a_rst_used(0),
        .s_rst_used(0),
        .en_used(0)
      ) i_data_out_reg (
        .d(data_out_reg[i-1]),
        .clk(clk),
        .en(en),
        .a_rst(1'b1),
        .s_rst(1'b1),
        .q(data_out_reg[i])
      );
    end
    mgc_generic_reg #(
      .width(64),
      .ph_clk(1),
      .ph_en(0),
      .ph_a_rst(0),
      .ph_s_rst(0),
      .a_rst_used(0),
      .s_rst_used(0),
      .en_used(0)
    ) i_data_out_reg_init (
      .d(data_out_t),
      .clk(clk),
      .en(en),
      .a_rst(1'b1),
      .s_rst(1'b1),
      .q(data_out_reg[0])
    );
    assign data_out = data_out_reg[n_outreg-1];
  end
  else
  begin
    assign data_out = data_out_t;
  end
  endgenerate
endmodule
module stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_7_16_10_1024_1024_16_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [15:0] q;
  output we;
  output [15:0] d;
  output [9:0] adr;
  input [9:0] adr_d;
  input [15:0] d_d;
  input en_d;
  input we_d;
  output [15:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule
module stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_6_64_10_1024_1024_64_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [9:0] adr;
  input [9:0] adr_d;
  input [63:0] d_d;
  input en_d;
  input we_d;
  output [63:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule
module stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_5_16_10_1024_1024_16_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [15:0] q;
  output we;
  output [15:0] d;
  output [9:0] adr;
  input [9:0] adr_d;
  input [15:0] d_d;
  input en_d;
  input we_d;
  output [15:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule
module stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_4_64_10_1024_1024_64_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [9:0] adr;
  input [9:0] adr_d;
  input [63:0] d_d;
  input en_d;
  input we_d;
  output [63:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule
module stage_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output, for_C_0_tr0, BUTTERFLY_C_24_tr0, BUTTERFLY_C_24_tr1,
      BUTTERFLY_1_C_24_tr0, BUTTERFLY_1_C_24_tr1, for_1_C_2_tr0
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [56:0] fsm_output;
  reg [56:0] fsm_output;
  input for_C_0_tr0;
  input BUTTERFLY_C_24_tr0;
  input BUTTERFLY_C_24_tr1;
  input BUTTERFLY_1_C_24_tr0;
  input BUTTERFLY_1_C_24_tr1;
  input for_1_C_2_tr0;
  parameter
    run_rlp_C_0 = 6'd0,
    main_C_0 = 6'd1,
    for_C_0 = 6'd2,
    BUTTERFLY_C_0 = 6'd3,
    BUTTERFLY_C_1 = 6'd4,
    BUTTERFLY_C_2 = 6'd5,
    BUTTERFLY_C_3 = 6'd6,
    BUTTERFLY_C_4 = 6'd7,
    BUTTERFLY_C_5 = 6'd8,
    BUTTERFLY_C_6 = 6'd9,
    BUTTERFLY_C_7 = 6'd10,
    BUTTERFLY_C_8 = 6'd11,
    BUTTERFLY_C_9 = 6'd12,
    BUTTERFLY_C_10 = 6'd13,
    BUTTERFLY_C_11 = 6'd14,
    BUTTERFLY_C_12 = 6'd15,
    BUTTERFLY_C_13 = 6'd16,
    BUTTERFLY_C_14 = 6'd17,
    BUTTERFLY_C_15 = 6'd18,
    BUTTERFLY_C_16 = 6'd19,
    BUTTERFLY_C_17 = 6'd20,
    BUTTERFLY_C_18 = 6'd21,
    BUTTERFLY_C_19 = 6'd22,
    BUTTERFLY_C_20 = 6'd23,
    BUTTERFLY_C_21 = 6'd24,
    BUTTERFLY_C_22 = 6'd25,
    BUTTERFLY_C_23 = 6'd26,
    BUTTERFLY_C_24 = 6'd27,
    BUTTERFLY_1_C_0 = 6'd28,
    BUTTERFLY_1_C_1 = 6'd29,
    BUTTERFLY_1_C_2 = 6'd30,
    BUTTERFLY_1_C_3 = 6'd31,
    BUTTERFLY_1_C_4 = 6'd32,
    BUTTERFLY_1_C_5 = 6'd33,
    BUTTERFLY_1_C_6 = 6'd34,
    BUTTERFLY_1_C_7 = 6'd35,
    BUTTERFLY_1_C_8 = 6'd36,
    BUTTERFLY_1_C_9 = 6'd37,
    BUTTERFLY_1_C_10 = 6'd38,
    BUTTERFLY_1_C_11 = 6'd39,
    BUTTERFLY_1_C_12 = 6'd40,
    BUTTERFLY_1_C_13 = 6'd41,
    BUTTERFLY_1_C_14 = 6'd42,
    BUTTERFLY_1_C_15 = 6'd43,
    BUTTERFLY_1_C_16 = 6'd44,
    BUTTERFLY_1_C_17 = 6'd45,
    BUTTERFLY_1_C_18 = 6'd46,
    BUTTERFLY_1_C_19 = 6'd47,
    BUTTERFLY_1_C_20 = 6'd48,
    BUTTERFLY_1_C_21 = 6'd49,
    BUTTERFLY_1_C_22 = 6'd50,
    BUTTERFLY_1_C_23 = 6'd51,
    BUTTERFLY_1_C_24 = 6'd52,
    for_1_C_0 = 6'd53,
    for_1_C_1 = 6'd54,
    for_1_C_2 = 6'd55,
    main_C_1 = 6'd56;
  reg [5:0] state_var;
  reg [5:0] state_var_NS;
  always @(*)
  begin : stage_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000000000010;
        state_var_NS = for_C_0;
      end
      for_C_0 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000000000100;
        if ( for_C_0_tr0 ) begin
          state_var_NS = BUTTERFLY_C_0;
        end
        else begin
          state_var_NS = BUTTERFLY_1_C_0;
        end
      end
      BUTTERFLY_C_0 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000000001000;
        state_var_NS = BUTTERFLY_C_1;
      end
      BUTTERFLY_C_1 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000000010000;
        state_var_NS = BUTTERFLY_C_2;
      end
      BUTTERFLY_C_2 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000000100000;
        state_var_NS = BUTTERFLY_C_3;
      end
      BUTTERFLY_C_3 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000001000000;
        state_var_NS = BUTTERFLY_C_4;
      end
      BUTTERFLY_C_4 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000010000000;
        state_var_NS = BUTTERFLY_C_5;
      end
      BUTTERFLY_C_5 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000100000000;
        state_var_NS = BUTTERFLY_C_6;
      end
      BUTTERFLY_C_6 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000001000000000;
        state_var_NS = BUTTERFLY_C_7;
      end
      BUTTERFLY_C_7 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000010000000000;
        state_var_NS = BUTTERFLY_C_8;
      end
      BUTTERFLY_C_8 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000100000000000;
        state_var_NS = BUTTERFLY_C_9;
      end
      BUTTERFLY_C_9 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000001000000000000;
        state_var_NS = BUTTERFLY_C_10;
      end
      BUTTERFLY_C_10 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000010000000000000;
        state_var_NS = BUTTERFLY_C_11;
      end
      BUTTERFLY_C_11 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000100000000000000;
        state_var_NS = BUTTERFLY_C_12;
      end
      BUTTERFLY_C_12 : begin
        fsm_output = 57'b000000000000000000000000000000000000000001000000000000000;
        state_var_NS = BUTTERFLY_C_13;
      end
      BUTTERFLY_C_13 : begin
        fsm_output = 57'b000000000000000000000000000000000000000010000000000000000;
        state_var_NS = BUTTERFLY_C_14;
      end
      BUTTERFLY_C_14 : begin
        fsm_output = 57'b000000000000000000000000000000000000000100000000000000000;
        state_var_NS = BUTTERFLY_C_15;
      end
      BUTTERFLY_C_15 : begin
        fsm_output = 57'b000000000000000000000000000000000000001000000000000000000;
        state_var_NS = BUTTERFLY_C_16;
      end
      BUTTERFLY_C_16 : begin
        fsm_output = 57'b000000000000000000000000000000000000010000000000000000000;
        state_var_NS = BUTTERFLY_C_17;
      end
      BUTTERFLY_C_17 : begin
        fsm_output = 57'b000000000000000000000000000000000000100000000000000000000;
        state_var_NS = BUTTERFLY_C_18;
      end
      BUTTERFLY_C_18 : begin
        fsm_output = 57'b000000000000000000000000000000000001000000000000000000000;
        state_var_NS = BUTTERFLY_C_19;
      end
      BUTTERFLY_C_19 : begin
        fsm_output = 57'b000000000000000000000000000000000010000000000000000000000;
        state_var_NS = BUTTERFLY_C_20;
      end
      BUTTERFLY_C_20 : begin
        fsm_output = 57'b000000000000000000000000000000000100000000000000000000000;
        state_var_NS = BUTTERFLY_C_21;
      end
      BUTTERFLY_C_21 : begin
        fsm_output = 57'b000000000000000000000000000000001000000000000000000000000;
        state_var_NS = BUTTERFLY_C_22;
      end
      BUTTERFLY_C_22 : begin
        fsm_output = 57'b000000000000000000000000000000010000000000000000000000000;
        state_var_NS = BUTTERFLY_C_23;
      end
      BUTTERFLY_C_23 : begin
        fsm_output = 57'b000000000000000000000000000000100000000000000000000000000;
        state_var_NS = BUTTERFLY_C_24;
      end
      BUTTERFLY_C_24 : begin
        fsm_output = 57'b000000000000000000000000000001000000000000000000000000000;
        if ( BUTTERFLY_C_24_tr0 ) begin
          state_var_NS = for_1_C_0;
        end
        else if ( BUTTERFLY_C_24_tr1 ) begin
          state_var_NS = BUTTERFLY_C_0;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      BUTTERFLY_1_C_0 : begin
        fsm_output = 57'b000000000000000000000000000010000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_1;
      end
      BUTTERFLY_1_C_1 : begin
        fsm_output = 57'b000000000000000000000000000100000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_2;
      end
      BUTTERFLY_1_C_2 : begin
        fsm_output = 57'b000000000000000000000000001000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_3;
      end
      BUTTERFLY_1_C_3 : begin
        fsm_output = 57'b000000000000000000000000010000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_4;
      end
      BUTTERFLY_1_C_4 : begin
        fsm_output = 57'b000000000000000000000000100000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_5;
      end
      BUTTERFLY_1_C_5 : begin
        fsm_output = 57'b000000000000000000000001000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_6;
      end
      BUTTERFLY_1_C_6 : begin
        fsm_output = 57'b000000000000000000000010000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_7;
      end
      BUTTERFLY_1_C_7 : begin
        fsm_output = 57'b000000000000000000000100000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_8;
      end
      BUTTERFLY_1_C_8 : begin
        fsm_output = 57'b000000000000000000001000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_9;
      end
      BUTTERFLY_1_C_9 : begin
        fsm_output = 57'b000000000000000000010000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_10;
      end
      BUTTERFLY_1_C_10 : begin
        fsm_output = 57'b000000000000000000100000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_11;
      end
      BUTTERFLY_1_C_11 : begin
        fsm_output = 57'b000000000000000001000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_12;
      end
      BUTTERFLY_1_C_12 : begin
        fsm_output = 57'b000000000000000010000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_13;
      end
      BUTTERFLY_1_C_13 : begin
        fsm_output = 57'b000000000000000100000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_14;
      end
      BUTTERFLY_1_C_14 : begin
        fsm_output = 57'b000000000000001000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_15;
      end
      BUTTERFLY_1_C_15 : begin
        fsm_output = 57'b000000000000010000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_16;
      end
      BUTTERFLY_1_C_16 : begin
        fsm_output = 57'b000000000000100000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_17;
      end
      BUTTERFLY_1_C_17 : begin
        fsm_output = 57'b000000000001000000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_18;
      end
      BUTTERFLY_1_C_18 : begin
        fsm_output = 57'b000000000010000000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_19;
      end
      BUTTERFLY_1_C_19 : begin
        fsm_output = 57'b000000000100000000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_20;
      end
      BUTTERFLY_1_C_20 : begin
        fsm_output = 57'b000000001000000000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_21;
      end
      BUTTERFLY_1_C_21 : begin
        fsm_output = 57'b000000010000000000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_22;
      end
      BUTTERFLY_1_C_22 : begin
        fsm_output = 57'b000000100000000000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_23;
      end
      BUTTERFLY_1_C_23 : begin
        fsm_output = 57'b000001000000000000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_24;
      end
      BUTTERFLY_1_C_24 : begin
        fsm_output = 57'b000010000000000000000000000000000000000000000000000000000;
        if ( BUTTERFLY_1_C_24_tr0 ) begin
          state_var_NS = for_1_C_0;
        end
        else if ( BUTTERFLY_1_C_24_tr1 ) begin
          state_var_NS = BUTTERFLY_1_C_0;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      for_1_C_0 : begin
        fsm_output = 57'b000100000000000000000000000000000000000000000000000000000;
        state_var_NS = for_1_C_1;
      end
      for_1_C_1 : begin
        fsm_output = 57'b001000000000000000000000000000000000000000000000000000000;
        state_var_NS = for_1_C_2;
      end
      for_1_C_2 : begin
        fsm_output = 57'b010000000000000000000000000000000000000000000000000000000;
        if ( for_1_C_2_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_1_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 57'b100000000000000000000000000000000000000000000000000000000;
        state_var_NS = main_C_0;
      end
      default : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end
endmodule
module stage_run_staller (
  clk, rst, arst_n, run_wen, run_wten, ap_start_rsci_wen_comp, ap_done_rsci_wen_comp,
      out1_rsci_wen_comp
);
  input clk;
  input rst;
  input arst_n;
  output run_wen;
  output run_wten;
  reg run_wten;
  input ap_start_rsci_wen_comp;
  input ap_done_rsci_wen_comp;
  input out1_rsci_wen_comp;
  assign run_wen = ap_start_rsci_wen_comp & ap_done_rsci_wen_comp & out1_rsci_wen_comp;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten <= 1'b0;
    end
    else if ( rst ) begin
      run_wten <= 1'b0;
    end
    else begin
      run_wten <= ~ run_wen;
    end
  end
endmodule
module stage_run_out_u_triosy_obj_out_u_triosy_wait_ctrl (
  run_wten, out_u_triosy_obj_iswt0, out_u_triosy_obj_biwt
);
  input run_wten;
  input out_u_triosy_obj_iswt0;
  output out_u_triosy_obj_biwt;
  assign out_u_triosy_obj_biwt = (~ run_wten) & out_u_triosy_obj_iswt0;
endmodule
module stage_run_out_f_d_triosy_obj_out_f_d_triosy_wait_ctrl (
  run_wten, out_f_d_triosy_obj_iswt0, out_f_d_triosy_obj_biwt
);
  input run_wten;
  input out_f_d_triosy_obj_iswt0;
  output out_f_d_triosy_obj_biwt;
  assign out_f_d_triosy_obj_biwt = (~ run_wten) & out_f_d_triosy_obj_iswt0;
endmodule
module stage_run_in_u_triosy_obj_in_u_triosy_wait_ctrl (
  run_wten, in_u_triosy_obj_iswt0, in_u_triosy_obj_biwt
);
  input run_wten;
  input in_u_triosy_obj_iswt0;
  output in_u_triosy_obj_biwt;
  assign in_u_triosy_obj_biwt = (~ run_wten) & in_u_triosy_obj_iswt0;
endmodule
module stage_run_in_f_d_triosy_obj_in_f_d_triosy_wait_ctrl (
  run_wten, in_f_d_triosy_obj_iswt0, in_f_d_triosy_obj_biwt
);
  input run_wten;
  input in_f_d_triosy_obj_iswt0;
  output in_f_d_triosy_obj_biwt;
  assign in_f_d_triosy_obj_biwt = (~ run_wten) & in_f_d_triosy_obj_iswt0;
endmodule
module stage_run_mode1_triosy_obj_mode1_triosy_wait_ctrl (
  run_wten, mode1_triosy_obj_iswt0, mode1_triosy_obj_biwt
);
  input run_wten;
  input mode1_triosy_obj_iswt0;
  output mode1_triosy_obj_biwt;
  assign mode1_triosy_obj_biwt = (~ run_wten) & mode1_triosy_obj_iswt0;
endmodule
module stage_run_out1_rsci_out1_wait_ctrl (
  out1_rsci_iswt0, out1_rsci_biwt, out1_rsci_irdy
);
  input out1_rsci_iswt0;
  output out1_rsci_biwt;
  input out1_rsci_irdy;
  assign out1_rsci_biwt = out1_rsci_iswt0 & out1_rsci_irdy;
endmodule
module stage_run_wait_dp (
  in_f_d_rsci_en_d, in_u_rsci_en_d, out_f_d_rsci_en_d, out_u_rsci_en_d, BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en,
      BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en, BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en,
      BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en, r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en,
      run_wen, in_f_d_rsci_cgo, in_f_d_rsci_cgo_ir_unreg, in_u_rsci_cgo, in_u_rsci_cgo_ir_unreg,
      out_f_d_rsci_cgo, out_f_d_rsci_cgo_ir_unreg, out_u_rsci_cgo, out_u_rsci_cgo_ir_unreg,
      BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo, BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo,
      BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo, BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo,
      r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_cgo
);
  output in_f_d_rsci_en_d;
  output in_u_rsci_en_d;
  output out_f_d_rsci_en_d;
  output out_u_rsci_en_d;
  output BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en;
  output BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en;
  output BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en;
  output BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en;
  output r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en;
  input run_wen;
  input in_f_d_rsci_cgo;
  input in_f_d_rsci_cgo_ir_unreg;
  input in_u_rsci_cgo;
  input in_u_rsci_cgo_ir_unreg;
  input out_f_d_rsci_cgo;
  input out_f_d_rsci_cgo_ir_unreg;
  input out_u_rsci_cgo;
  input out_u_rsci_cgo_ir_unreg;
  input BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo;
  input BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo;
  input BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo;
  input BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo;
  input r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_cgo;
  assign in_f_d_rsci_en_d = run_wen & (in_f_d_rsci_cgo | in_f_d_rsci_cgo_ir_unreg);
  assign in_u_rsci_en_d = run_wen & (in_u_rsci_cgo | in_u_rsci_cgo_ir_unreg);
  assign out_f_d_rsci_en_d = run_wen & (out_f_d_rsci_cgo | out_f_d_rsci_cgo_ir_unreg);
  assign out_u_rsci_en_d = run_wen & (out_u_rsci_cgo | out_u_rsci_cgo_ir_unreg);
  assign BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en = ~(run_wen & BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo);
  assign BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en = ~(run_wen & BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo);
  assign BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en = ~(run_wen & BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo);
  assign BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en = ~(run_wen & BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo);
  assign r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en = ~(run_wen &
      r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_cgo);
endmodule
module stage_run_ap_done_rsci_ap_done_wait_ctrl (
  ap_done_rsci_iswt0, ap_done_rsci_biwt, ap_done_rsci_irdy
);
  input ap_done_rsci_iswt0;
  output ap_done_rsci_biwt;
  input ap_done_rsci_irdy;
  assign ap_done_rsci_biwt = ap_done_rsci_iswt0 & ap_done_rsci_irdy;
endmodule
module stage_run_ap_start_rsci_ap_start_wait_ctrl (
  ap_start_rsci_iswt0, ap_start_rsci_biwt, ap_start_rsci_ivld
);
  input ap_start_rsci_iswt0;
  output ap_start_rsci_biwt;
  input ap_start_rsci_ivld;
  assign ap_start_rsci_biwt = ap_start_rsci_iswt0 & ap_start_rsci_ivld;
endmodule
module stage_run_out_u_triosy_obj (
  out_u_triosy_lz, run_wten, out_u_triosy_obj_iswt0
);
  output out_u_triosy_lz;
  input run_wten;
  input out_u_triosy_obj_iswt0;
  wire out_u_triosy_obj_biwt;
  mgc_io_sync_v2 #(.valid(32'sd0)) out_u_triosy_obj (
      .ld(out_u_triosy_obj_biwt),
      .lz(out_u_triosy_lz)
    );
  stage_run_out_u_triosy_obj_out_u_triosy_wait_ctrl stage_run_out_u_triosy_obj_out_u_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .out_u_triosy_obj_iswt0(out_u_triosy_obj_iswt0),
      .out_u_triosy_obj_biwt(out_u_triosy_obj_biwt)
    );
endmodule
module stage_run_out_f_d_triosy_obj (
  out_f_d_triosy_lz, run_wten, out_f_d_triosy_obj_iswt0
);
  output out_f_d_triosy_lz;
  input run_wten;
  input out_f_d_triosy_obj_iswt0;
  wire out_f_d_triosy_obj_biwt;
  mgc_io_sync_v2 #(.valid(32'sd0)) out_f_d_triosy_obj (
      .ld(out_f_d_triosy_obj_biwt),
      .lz(out_f_d_triosy_lz)
    );
  stage_run_out_f_d_triosy_obj_out_f_d_triosy_wait_ctrl stage_run_out_f_d_triosy_obj_out_f_d_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .out_f_d_triosy_obj_iswt0(out_f_d_triosy_obj_iswt0),
      .out_f_d_triosy_obj_biwt(out_f_d_triosy_obj_biwt)
    );
endmodule
module stage_run_in_u_triosy_obj (
  in_u_triosy_lz, run_wten, in_u_triosy_obj_iswt0
);
  output in_u_triosy_lz;
  input run_wten;
  input in_u_triosy_obj_iswt0;
  wire in_u_triosy_obj_biwt;
  mgc_io_sync_v2 #(.valid(32'sd0)) in_u_triosy_obj (
      .ld(in_u_triosy_obj_biwt),
      .lz(in_u_triosy_lz)
    );
  stage_run_in_u_triosy_obj_in_u_triosy_wait_ctrl stage_run_in_u_triosy_obj_in_u_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .in_u_triosy_obj_iswt0(in_u_triosy_obj_iswt0),
      .in_u_triosy_obj_biwt(in_u_triosy_obj_biwt)
    );
endmodule
module stage_run_in_f_d_triosy_obj (
  in_f_d_triosy_lz, run_wten, in_f_d_triosy_obj_iswt0
);
  output in_f_d_triosy_lz;
  input run_wten;
  input in_f_d_triosy_obj_iswt0;
  wire in_f_d_triosy_obj_biwt;
  mgc_io_sync_v2 #(.valid(32'sd0)) in_f_d_triosy_obj (
      .ld(in_f_d_triosy_obj_biwt),
      .lz(in_f_d_triosy_lz)
    );
  stage_run_in_f_d_triosy_obj_in_f_d_triosy_wait_ctrl stage_run_in_f_d_triosy_obj_in_f_d_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .in_f_d_triosy_obj_iswt0(in_f_d_triosy_obj_iswt0),
      .in_f_d_triosy_obj_biwt(in_f_d_triosy_obj_biwt)
    );
endmodule
module stage_run_mode1_triosy_obj (
  mode1_triosy_lz, run_wten, mode1_triosy_obj_iswt0
);
  output mode1_triosy_lz;
  input run_wten;
  input mode1_triosy_obj_iswt0;
  wire mode1_triosy_obj_biwt;
  mgc_io_sync_v2 #(.valid(32'sd0)) mode1_triosy_obj (
      .ld(mode1_triosy_obj_biwt),
      .lz(mode1_triosy_lz)
    );
  stage_run_mode1_triosy_obj_mode1_triosy_wait_ctrl stage_run_mode1_triosy_obj_mode1_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .mode1_triosy_obj_iswt0(mode1_triosy_obj_iswt0),
      .mode1_triosy_obj_biwt(mode1_triosy_obj_biwt)
    );
endmodule
module stage_run_out1_rsci (
  out1_rsc_dat, out1_rsc_vld, out1_rsc_rdy, out1_rsci_oswt, out1_rsci_wen_comp, out1_rsci_idat
);
  output [79:0] out1_rsc_dat;
  output out1_rsc_vld;
  input out1_rsc_rdy;
  input out1_rsci_oswt;
  output out1_rsci_wen_comp;
  input [79:0] out1_rsci_idat;
  wire out1_rsci_biwt;
  wire out1_rsci_irdy;
  ccs_out_wait_v1 #(.rscid(32'sd8),
  .width(32'sd80)) out1_rsci (
      .irdy(out1_rsci_irdy),
      .ivld(out1_rsci_oswt),
      .idat(out1_rsci_idat),
      .rdy(out1_rsc_rdy),
      .vld(out1_rsc_vld),
      .dat(out1_rsc_dat)
    );
  stage_run_out1_rsci_out1_wait_ctrl stage_run_out1_rsci_out1_wait_ctrl_inst (
      .out1_rsci_iswt0(out1_rsci_oswt),
      .out1_rsci_biwt(out1_rsci_biwt),
      .out1_rsci_irdy(out1_rsci_irdy)
    );
  assign out1_rsci_wen_comp = (~ out1_rsci_oswt) | out1_rsci_biwt;
endmodule
module stage_run_ap_done_rsci (
  ap_done_rsc_dat, ap_done_rsc_vld, ap_done_rsc_rdy, ap_done_rsci_oswt, ap_done_rsci_wen_comp
);
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input ap_done_rsci_oswt;
  output ap_done_rsci_wen_comp;
  wire ap_done_rsci_biwt;
  wire ap_done_rsci_irdy;
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd1)) ap_done_rsci (
      .irdy(ap_done_rsci_irdy),
      .ivld(ap_done_rsci_oswt),
      .idat(1'b1),
      .rdy(ap_done_rsc_rdy),
      .vld(ap_done_rsc_vld),
      .dat(ap_done_rsc_dat)
    );
  stage_run_ap_done_rsci_ap_done_wait_ctrl stage_run_ap_done_rsci_ap_done_wait_ctrl_inst
      (
      .ap_done_rsci_iswt0(ap_done_rsci_oswt),
      .ap_done_rsci_biwt(ap_done_rsci_biwt),
      .ap_done_rsci_irdy(ap_done_rsci_irdy)
    );
  assign ap_done_rsci_wen_comp = (~ ap_done_rsci_oswt) | ap_done_rsci_biwt;
endmodule
module stage_run_ap_start_rsci (
  ap_start_rsc_dat, ap_start_rsc_vld, ap_start_rsc_rdy, ap_start_rsci_oswt, ap_start_rsci_wen_comp
);
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  input ap_start_rsci_oswt;
  output ap_start_rsci_wen_comp;
  wire ap_start_rsci_biwt;
  wire ap_start_rsci_ivld;
  wire ap_start_rsci_idat;
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd1)) ap_start_rsci (
      .rdy(ap_start_rsc_rdy),
      .vld(ap_start_rsc_vld),
      .dat(ap_start_rsc_dat),
      .irdy(ap_start_rsci_oswt),
      .ivld(ap_start_rsci_ivld),
      .idat(ap_start_rsci_idat)
    );
  stage_run_ap_start_rsci_ap_start_wait_ctrl stage_run_ap_start_rsci_ap_start_wait_ctrl_inst
      (
      .ap_start_rsci_iswt0(ap_start_rsci_oswt),
      .ap_start_rsci_biwt(ap_start_rsci_biwt),
      .ap_start_rsci_ivld(ap_start_rsci_ivld)
    );
  assign ap_start_rsci_wen_comp = (~ ap_start_rsci_oswt) | ap_start_rsci_biwt;
endmodule
module stage_run (
  clk, rst, arst_n, ap_start_rsc_dat, ap_start_rsc_vld, ap_start_rsc_rdy, ap_done_rsc_dat,
      ap_done_rsc_vld, ap_done_rsc_rdy, mode1_rsc_dat, mode1_triosy_lz, in_f_d_triosy_lz,
      in_u_triosy_lz, out_f_d_triosy_lz, out_u_triosy_lz, out1_rsc_dat, out1_rsc_vld,
      out1_rsc_rdy, in_f_d_rsci_adr_d, in_f_d_rsci_d_d, in_f_d_rsci_en_d, in_f_d_rsci_q_d,
      in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, in_u_rsci_adr_d, in_u_rsci_d_d,
      in_u_rsci_en_d, in_u_rsci_q_d, in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      out_f_d_rsci_adr_d, out_f_d_rsci_d_d, out_f_d_rsci_en_d, out_f_d_rsci_q_d,
      out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, out_u_rsci_adr_d, out_u_rsci_d_d,
      out_u_rsci_en_d, out_u_rsci_q_d, out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr, BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out,
      BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en, BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out,
      BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en, BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out,
      BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en, BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out,
      BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en, r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_addr,
      r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out, r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en,
      BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out, in_f_d_rsci_we_d_pff,
      in_u_rsci_we_d_pff, out_f_d_rsci_we_d_pff, out_u_rsci_we_d_pff
);
  input clk;
  input rst;
  input arst_n;
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input [15:0] mode1_rsc_dat;
  output mode1_triosy_lz;
  output in_f_d_triosy_lz;
  output in_u_triosy_lz;
  output out_f_d_triosy_lz;
  output out_u_triosy_lz;
  output [79:0] out1_rsc_dat;
  output out1_rsc_vld;
  input out1_rsc_rdy;
  output [9:0] in_f_d_rsci_adr_d;
  output [63:0] in_f_d_rsci_d_d;
  output in_f_d_rsci_en_d;
  input [63:0] in_f_d_rsci_q_d;
  output in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [9:0] in_u_rsci_adr_d;
  output [15:0] in_u_rsci_d_d;
  output in_u_rsci_en_d;
  input [15:0] in_u_rsci_q_d;
  output in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [9:0] out_f_d_rsci_adr_d;
  output [63:0] out_f_d_rsci_d_d;
  output out_f_d_rsci_en_d;
  input [63:0] out_f_d_rsci_q_d;
  output out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [9:0] out_u_rsci_adr_d;
  output [15:0] out_u_rsci_d_d;
  output out_u_rsci_en_d;
  input [15:0] out_u_rsci_q_d;
  output out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [9:0] BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr;
  input [13:0] BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out;
  output BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en;
  input [13:0] BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out;
  output BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en;
  input [13:0] BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out;
  output BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en;
  input [13:0] BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out;
  output BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en;
  output [9:0] r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_addr;
  input [61:0] r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out;
  output r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en;
  input [63:0] BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out;
  output in_f_d_rsci_we_d_pff;
  output in_u_rsci_we_d_pff;
  output out_f_d_rsci_we_d_pff;
  output out_u_rsci_we_d_pff;
  wire run_wen;
  wire run_wten;
  wire ap_start_rsci_wen_comp;
  wire ap_done_rsci_wen_comp;
  wire [15:0] mode1_rsci_idat;
  wire out1_rsci_wen_comp;
  reg BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo;
  reg BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo;
  reg BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo;
  reg BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo;
  reg [15:0] out1_rsci_idat_79_64;
  wire [56:0] fsm_output;
  wire [11:0] return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp;
  wire [12:0] nl_return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp;
  wire return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_9_e1_eq_e2_equal_tmp;
  wire return_extract_19_return_extract_19_nor_tmp;
  wire return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp;
  wire operator_11_true_19_operator_11_true_19_and_tmp;
  wire return_mult_generic_AC_RND_CONV_false_1_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_1_exp_ovf_oif_aelse_and_1_tmp;
  wire return_mult_generic_AC_RND_CONV_false_1_exp_ovf_return_mult_generic_AC_RND_CONV_false_1_exp_ovf_or_tmp;
  wire [11:0] return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_acc_tmp;
  wire [12:0] nl_return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_acc_tmp;
  wire return_extract_17_return_extract_17_nor_tmp;
  wire operator_11_true_17_operator_11_true_17_and_tmp;
  wire return_extract_15_return_extract_15_nor_tmp;
  wire operator_11_true_15_operator_11_true_15_and_tmp;
  wire [12:0] operator_33_true_12_acc_tmp;
  wire [13:0] nl_operator_33_true_12_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_6_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_3_if_5_return_add_generic_AC_RND_CONV_false_3_if_5_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_2_if_5_return_add_generic_AC_RND_CONV_false_2_if_5_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_if_5_return_add_generic_AC_RND_CONV_false_if_5_and_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_2_aif_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_tmp;
  wire return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_1_e1_eq_e2_equal_tmp;
  wire operator_11_true_3_operator_11_true_3_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_23_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_22_e1_eq_e2_equal_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp;
  wire [12:0] nl_return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp;
  wire return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp;
  wire [12:0] nl_return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp;
  wire return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp;
  wire return_extract_51_return_extract_51_nor_tmp;
  wire return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp;
  wire operator_11_true_51_operator_11_true_51_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp;
  wire return_extract_49_return_extract_49_nor_tmp;
  wire return_extract_49_m_zero_return_extract_49_m_zero_nor_tmp;
  wire operator_11_true_49_operator_11_true_49_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_18_if_5_return_add_generic_AC_RND_CONV_false_18_if_5_and_tmp;
  wire return_extract_47_return_extract_47_nor_tmp;
  wire return_extract_47_m_zero_return_extract_47_m_zero_nor_tmp;
  wire operator_11_true_47_operator_11_true_47_and_tmp;
  wire [12:0] operator_33_true_38_acc_tmp;
  wire [13:0] nl_operator_33_true_38_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_19_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_17_if_5_return_add_generic_AC_RND_CONV_false_17_if_5_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_16_if_5_return_add_generic_AC_RND_CONV_false_16_if_5_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_16_else_4_return_add_generic_AC_RND_CONV_false_16_else_4_nand_tmp;
  wire [12:0] operator_33_true_32_acc_tmp;
  wire [13:0] nl_operator_33_true_32_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_15_if_5_return_add_generic_AC_RND_CONV_false_15_if_5_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_15_aif_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_if_1_return_add_generic_AC_RND_CONV_false_17_op2_normal_return_extract_41_nor_tmp;
  wire [10:0] return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp;
  wire [11:0] nl_return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_17_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_14_e1_eq_e2_equal_tmp;
  wire operator_11_true_35_operator_11_true_35_and_tmp;
  wire stage_PE_1_and_1_tmp;
  wire operator_16_false_operator_16_false_nor_tmp;
  wire and_dcpl_18;
  wire or_tmp_21;
  wire or_tmp_26;
  wire or_tmp_30;
  wire mux_tmp_12;
  wire mux_tmp_15;
  wire mux_tmp_19;
  wire mux_tmp_22;
  wire and_tmp_1;
  wire and_dcpl_57;
  wire and_dcpl_64;
  wire or_dcpl_93;
  wire and_dcpl_75;
  wire and_dcpl_159;
  wire and_dcpl_160;
  wire and_dcpl_166;
  wire and_dcpl_172;
  wire and_dcpl_175;
  wire or_dcpl_179;
  wire or_dcpl_180;
  wire or_dcpl_184;
  wire or_dcpl_190;
  wire or_dcpl_192;
  wire and_dcpl_177;
  wire and_dcpl_183;
  wire or_dcpl_198;
  wire or_dcpl_200;
  wire or_dcpl_201;
  wire or_dcpl_204;
  wire or_dcpl_207;
  wire and_dcpl_185;
  wire or_dcpl_208;
  wire or_dcpl_209;
  wire or_dcpl_221;
  wire or_dcpl_223;
  wire or_dcpl_224;
  wire or_dcpl_227;
  wire or_dcpl_228;
  wire or_dcpl_230;
  wire or_dcpl_233;
  wire or_dcpl_235;
  wire or_dcpl_236;
  wire or_dcpl_239;
  wire or_dcpl_240;
  wire or_dcpl_245;
  wire or_dcpl_248;
  wire and_dcpl_202;
  wire or_dcpl_253;
  wire or_dcpl_269;
  wire or_dcpl_272;
  wire or_dcpl_273;
  wire or_dcpl_283;
  wire and_dcpl_203;
  wire and_dcpl_204;
  wire or_dcpl_284;
  wire or_dcpl_285;
  wire or_dcpl_289;
  wire and_dcpl_210;
  wire or_dcpl_296;
  wire and_dcpl_216;
  wire or_dcpl_301;
  wire and_dcpl_217;
  wire or_dcpl_308;
  wire or_dcpl_311;
  wire or_dcpl_312;
  wire and_dcpl_219;
  wire or_dcpl_320;
  wire and_dcpl_222;
  wire and_dcpl_223;
  wire and_dcpl_224;
  wire or_dcpl_324;
  wire and_dcpl_229;
  wire and_dcpl_231;
  wire and_dcpl_235;
  wire and_dcpl_237;
  wire or_dcpl_337;
  wire or_dcpl_342;
  wire and_dcpl_251;
  wire or_dcpl_359;
  wire and_dcpl_253;
  wire or_dcpl_367;
  wire or_dcpl_371;
  wire and_dcpl_259;
  wire and_dcpl_263;
  wire and_dcpl_266;
  wire and_dcpl_268;
  wire and_dcpl_274;
  wire and_dcpl_276;
  wire and_dcpl_285;
  wire or_dcpl_438;
  wire and_dcpl_323;
  wire and_dcpl_327;
  wire and_dcpl_329;
  wire and_dcpl_330;
  wire and_dcpl_333;
  wire or_dcpl_466;
  wire or_dcpl_470;
  wire or_dcpl_473;
  wire or_dcpl_476;
  wire and_dcpl_340;
  wire and_dcpl_341;
  wire and_dcpl_344;
  wire and_dcpl_354;
  wire and_dcpl_360;
  wire and_dcpl_369;
  wire and_dcpl_382;
  wire and_dcpl_389;
  wire and_dcpl_393;
  wire or_dcpl_484;
  wire and_dcpl_402;
  wire and_dcpl_403;
  wire and_dcpl_405;
  wire and_dcpl_420;
  wire and_dcpl_421;
  wire or_dcpl_485;
  wire or_dcpl_492;
  wire or_dcpl_493;
  wire or_dcpl_497;
  wire or_dcpl_502;
  wire or_dcpl_503;
  wire or_dcpl_504;
  wire or_dcpl_509;
  wire or_dcpl_511;
  wire or_dcpl_515;
  wire or_dcpl_516;
  wire or_dcpl_519;
  wire or_dcpl_520;
  wire or_dcpl_521;
  wire or_dcpl_522;
  wire and_dcpl_446;
  wire and_dcpl_447;
  wire or_dcpl_528;
  wire or_dcpl_529;
  wire or_dcpl_532;
  wire or_dcpl_534;
  wire or_dcpl_535;
  wire or_dcpl_545;
  wire or_dcpl_553;
  wire or_dcpl_554;
  wire or_dcpl_555;
  wire or_dcpl_559;
  wire or_dcpl_560;
  wire or_dcpl_562;
  wire and_dcpl_448;
  wire and_dcpl_452;
  wire or_dcpl_573;
  wire or_dcpl_575;
  wire or_dcpl_576;
  wire or_dcpl_579;
  wire or_dcpl_580;
  wire or_dcpl_584;
  wire or_dcpl_585;
  wire or_dcpl_586;
  wire or_dcpl_588;
  wire or_dcpl_590;
  wire and_dcpl_460;
  wire or_dcpl_596;
  wire or_dcpl_597;
  wire or_dcpl_598;
  wire or_dcpl_602;
  wire or_dcpl_604;
  wire or_dcpl_605;
  wire or_dcpl_606;
  wire or_dcpl_618;
  wire or_dcpl_619;
  wire or_dcpl_620;
  wire or_dcpl_621;
  wire or_dcpl_625;
  wire or_dcpl_626;
  wire or_dcpl_627;
  wire or_dcpl_628;
  wire and_dcpl_466;
  wire and_dcpl_467;
  wire and_dcpl_468;
  wire and_dcpl_469;
  wire or_dcpl_632;
  wire or_dcpl_633;
  wire or_dcpl_634;
  wire or_dcpl_635;
  wire or_dcpl_640;
  wire or_dcpl_645;
  wire or_dcpl_654;
  wire or_dcpl_664;
  wire and_dcpl_474;
  wire and_dcpl_475;
  wire and_dcpl_478;
  wire and_dcpl_479;
  wire or_dcpl_671;
  wire or_dcpl_673;
  wire or_dcpl_678;
  wire or_dcpl_679;
  wire or_dcpl_680;
  wire or_dcpl_684;
  wire or_dcpl_685;
  wire or_dcpl_686;
  wire or_dcpl_698;
  wire or_dcpl_699;
  wire or_dcpl_702;
  wire or_dcpl_708;
  wire or_dcpl_709;
  wire and_dcpl_501;
  wire or_dcpl_711;
  wire or_dcpl_719;
  wire or_dcpl_725;
  wire or_dcpl_726;
  wire or_dcpl_728;
  wire or_dcpl_740;
  wire or_dcpl_744;
  wire or_dcpl_750;
  wire or_dcpl_762;
  wire or_dcpl_763;
  wire or_dcpl_776;
  wire or_dcpl_788;
  wire or_dcpl_789;
  wire or_dcpl_800;
  wire or_dcpl_809;
  wire and_dcpl_503;
  wire or_dcpl_845;
  wire or_dcpl_848;
  wire or_dcpl_849;
  wire or_dcpl_854;
  wire or_dcpl_866;
  wire or_dcpl_870;
  wire or_dcpl_874;
  wire or_dcpl_876;
  wire or_dcpl_890;
  wire or_dcpl_906;
  wire or_dcpl_928;
  wire or_dcpl_933;
  wire or_dcpl_943;
  wire or_dcpl_967;
  wire or_dcpl_970;
  wire or_dcpl_980;
  wire or_dcpl_981;
  wire or_dcpl_982;
  wire and_dcpl_531;
  wire not_tmp_376;
  wire and_dcpl_534;
  wire and_dcpl_541;
  wire and_dcpl_543;
  wire not_tmp_395;
  wire or_tmp_64;
  wire or_tmp_231;
  wire or_tmp_334;
  wire or_tmp_450;
  wire or_tmp_759;
  wire or_tmp_762;
  wire or_tmp_946;
  wire and_660_cse;
  wire and_647_cse;
  wire and_680_cse;
  wire and_630_cse;
  wire and_662_cse;
  wire and_746_cse;
  wire and_741_cse;
  wire and_836_cse;
  wire and_840_cse;
  wire and_2185_cse;
  wire and_2184_cse;
  wire return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_6_lor_lpi_2_dfm_1;
  wire return_extract_3_m_zero_sva_mx1w0;
  wire return_mult_generic_AC_RND_CONV_false_6_op1_nan_sva_1;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3;
  wire return_mult_generic_AC_RND_CONV_false_6_e_incr_lpi_2_dfm_2;
  wire return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_or_2;
  wire return_add_generic_AC_RND_CONV_false_12_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_12_r_zero_1_sva;
  reg operator_11_true_return_22_sva;
  reg return_add_generic_AC_RND_CONV_false_10_op2_inf_sva;
  reg return_add_generic_AC_RND_CONV_false_10_op1_nan_sva;
  reg return_add_generic_AC_RND_CONV_false_10_op2_nan_sva;
  reg return_add_generic_AC_RND_CONV_false_12_else_4_unequal_tmp;
  reg return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  wire return_add_generic_AC_RND_CONV_false_11_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva;
  reg return_add_generic_AC_RND_CONV_false_22_op1_inf_sva;
  reg operator_11_true_return_26_sva;
  reg return_add_generic_AC_RND_CONV_false_14_op1_nan_sva;
  reg return_add_generic_AC_RND_CONV_false_10_unequal_tmp;
  reg return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_10_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  wire return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0;
  wire return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_mx2w0;
  reg return_add_generic_AC_RND_CONV_false_10_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_9_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0;
  wire return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0;
  reg return_add_generic_AC_RND_CONV_false_9_else_4_unequal_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_8_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_8_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_21_op1_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_21_op1_nan_sva_1;
  reg return_add_generic_AC_RND_CONV_false_8_else_4_unequal_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_9_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_7_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_7_else_4_unequal_tmp;
  reg operator_11_true_return_21_sva;
  reg return_extract_21_m_zero_sva;
  wire return_add_generic_AC_RND_CONV_false_17_mux_6_itm_mx2;
  wire return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1;
  reg return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm;
  reg return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm;
  wire return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_8_e_dif_qr_lpi_3_dfm_mx0;
  reg return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm;
  reg return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm;
  wire return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_7_e_dif_qr_lpi_3_dfm_mx0;
  wire return_mult_generic_AC_RND_CONV_false_2_m_r_51_lpi_3_dfm_mx1;
  wire [50:0] return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1;
  wire BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx2;
  reg return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_2_if_nor_ovfl_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_2_op2_inf_sva_1;
  reg return_add_generic_AC_RND_CONV_false_17_mux_6_itm;
  reg return_add_generic_AC_RND_CONV_false_10_do_sub_sva;
  reg [105:0] return_mult_generic_AC_RND_CONV_false_1_p_1_sva;
  wire return_add_generic_AC_RND_CONV_false_6_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm;
  reg return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp;
  wire drf_qr_lval_15_smx_0_lpi_3_dfm_mx2;
  wire [50:0] return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_1_op2_zero_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_1_op1_zero_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_1_op2_inf_sva_1;
  reg return_extract_12_m_zero_sva;
  wire return_add_generic_AC_RND_CONV_false_17_if_5_return_add_generic_AC_RND_CONV_false_17_if_5_nor_2;
  wire return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_op2_zero_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_op2_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_6_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx1;
  wire return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm_mx1;
  wire [49:0] return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_49_0_mx0;
  wire return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_6_e_dif_qr_lpi_3_dfm_mx0;
  reg stage_PE_1_tmp_re_d_1_lpi_3_dfm_63;
  wire stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0;
  reg operator_11_true_return_1_sva;
  wire return_add_generic_AC_RND_CONV_false_18_if_5_return_add_generic_AC_RND_CONV_false_18_if_5_nor_2;
  wire return_add_generic_AC_RND_CONV_false_3_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_2_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_2_r_inf_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_else_4_unequal_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_1_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_1_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_1_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_25_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_25_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_24_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_24_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_23_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1;
  reg return_add_generic_AC_RND_CONV_false_23_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_22_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1;
  reg return_add_generic_AC_RND_CONV_false_22_else_4_unequal_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_21_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1;
  reg return_extract_26_m_zero_sva;
  wire return_add_generic_AC_RND_CONV_false_21_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_21_else_4_unequal_tmp;
  reg return_extract_22_m_zero_sva;
  wire [11:0] return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1;
  reg operator_11_true_return_24_sva;
  reg return_add_generic_AC_RND_CONV_false_12_mux_itm;
  wire return_add_generic_AC_RND_CONV_false_20_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_20_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_17_mux_6_itm_mx4;
  wire return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2;
  wire return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1;
  reg drf_qr_lval_13_smx_0_lpi_3_dfm;
  wire return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_mx1;
  wire return_mult_generic_AC_RND_CONV_false_5_lor_lpi_3_dfm_1;
  reg return_add_generic_AC_RND_CONV_false_11_do_sub_sva;
  wire [50:0] return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_5_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_4_lor_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_19_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp;
  wire BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx5;
  wire return_mult_generic_AC_RND_CONV_false_4_op2_zero_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_4_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_3_lor_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_3_op2_zero_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_3_op2_inf_sva_1;
  wire drf_qr_lval_13_smx_0_lpi_3_dfm_mx3;
  wire return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm_mx3;
  wire [49:0] return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0_mx0;
  wire return_add_generic_AC_RND_CONV_false_19_op2_mu_0_lpi_3_dfm_1;
  wire stage_PE_1_tmp_im_d_1_lpi_3_dfm_63_mx0;
  wire stage_PE_1_tmp_im_d_1_lpi_3_dfm_51_mx1;
  wire return_add_generic_AC_RND_CONV_false_16_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_15_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_15_r_inf_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_13_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_13_else_4_unequal_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_13_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_14_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_14_else_4_unequal_tmp;
  reg inverse_lpi_1_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_14_e_dif_qr_lpi_3_dfm_mx0;
  wire [3:0] for_i_3_0_sva_2;
  wire [4:0] nl_for_i_3_0_sva_2;
  wire operator_16_false_1_operator_16_false_1_and_mdf_sva_1;
  reg operator_16_false_operator_16_false_nor_cse_sva;
  reg BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm;
  reg mode_lpi_1_dfm;
  reg [12:0] operator_33_true_12_acc_psp_sva;
  reg [3:0] for_i_3_0_sva;
  reg [15:0] operator_16_false_io_read_mode1_rsc_cse_sva;
  reg return_add_generic_AC_RND_CONV_false_16_do_sub_sva;
  reg return_add_generic_AC_RND_CONV_false_12_do_sub_sva;
  reg return_add_generic_AC_RND_CONV_false_20_do_sub_sva;
  reg return_add_generic_AC_RND_CONV_false_18_mux_itm;
  wire [11:0] operator_6_false_58_acc_psp_sva_1;
  wire [12:0] nl_operator_6_false_58_acc_psp_sva_1;
  reg return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva;
  wire return_add_generic_AC_RND_CONV_false_1_mux_28;
  wire [9:0] return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1;
  reg [63:0] stage_PE_1_tmp_re_d_sva;
  reg [63:0] stage_PE_1_x_re_d_sva;
  reg return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva;
  reg return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva;
  wire return_mult_generic_AC_RND_CONV_false_if_1_aelse_return_mult_generic_AC_RND_CONV_false_if_1_aelse_or_2;
  reg [5:0] return_add_generic_AC_RND_CONV_false_10_ls_sva;
  reg return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva;
  wire stage_d_mul_return_d_1_63_sva_1;
  wire stage_d_mul_return_d_2_63_sva_1;
  wire stage_d_mul_return_d_63_sva_1;
  wire stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50;
  wire [50:0] return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1;
  reg return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_1;
  wire return_mult_generic_AC_RND_CONV_false_1_zero_m_return_mult_generic_AC_RND_CONV_false_1_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_1_r_zero_return_mult_generic_AC_RND_CONV_false_1_r_zero_nor_mdf_sva_1;
  reg return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1;
  reg return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva;
  reg [11:0] operator_33_true_36_acc_psp_1_sva;
  wire stage_d_mul_return_d_4_63_sva_2;
  wire stage_d_mul_return_d_5_63_sva_1;
  wire stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50;
  wire [50:0] return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx2;
  wire return_add_generic_AC_RND_CONV_false_1_if_5_or_3;
  wire return_add_generic_AC_RND_CONV_false_4_unequal_tmp_1;
  wire for_1_if_and_ssc;
  reg out1_rsci_idat_63;
  reg [10:0] out1_rsci_idat_62_52;
  reg out1_rsci_idat_51;
  reg [50:0] out1_rsci_idat_50_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_12_e_dif_qr_lpi_3_dfm_mx0_10_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_2_e_dif_qr_lpi_3_dfm_mx0_10_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt;
  wire [11:0] nl_return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt;
  wire [9:0] return_add_generic_AC_RND_CONV_false_4_e_dif_qif_acc_pmx_lpi_3_dfm_mx0_9_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_3_e_dif_qr_lpi_3_dfm_mx0_10_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_24_e_dif_qr_lpi_3_dfm_mx0_10_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_15_e_dif_qr_lpi_3_dfm_mx0_10_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_16_e_dif_qr_lpi_3_dfm_mx0_10_0;
  wire [9:0] drf_qr_lval_10_smx_lpi_3_dfm_mx3_10_1;
  wire drf_qr_lval_10_smx_lpi_3_dfm_mx3_0;
  wire [9:0] drf_qr_lval_10_smx_lpi_3_dfm_mx7_10_1;
  wire drf_qr_lval_10_smx_lpi_3_dfm_mx7_0;
  wire return_add_generic_AC_RND_CONV_false_12_res_mant_and_ssc;
  reg reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_cgo_cse;
  reg reg_out_u_triosy_obj_iswt0_cse;
  reg reg_out1_rsci_iswt0_cse;
  reg reg_out_u_rsci_cgo_ir_cse;
  reg reg_out_f_d_rsci_cgo_ir_cse;
  reg reg_in_u_rsci_cgo_ir_cse;
  reg reg_in_f_d_rsci_cgo_ir_cse;
  reg reg_ap_start_rsci_iswt0_cse;
  reg [9:0] reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_addr_cse;
  reg [9:0] reg_BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_addr_cse;
  wire operator_16_false_and_cse;
  wire t_in_and_cse;
  wire mode_and_cse;
  wire stage_PE_1_and_2_cse;
  wire return_add_generic_AC_RND_CONV_false_10_and_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_cse;
  wire return_add_generic_AC_RND_CONV_false_12_op_bigger_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_cse;
  wire or_547_cse;
  wire return_add_generic_AC_RND_CONV_false_12_do_sub_mux1h_1_cse;
  wire return_add_generic_AC_RND_CONV_false_12_do_sub_mux1h_6_cse;
  wire or_1993_cse;
  wire return_extract_19_and_cse;
  wire return_add_generic_AC_RND_CONV_false_10_op2_nan_and_cse;
  wire or_673_cse;
  wire or_1102_cse;
  wire return_add_generic_AC_RND_CONV_false_23_op1_mu_and_cse;
  wire and_6_cse;
  wire return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse;
  wire [50:0] stage_PE_gm_re_d_mux_cse;
  wire stage_PE_gm_im_d_mux_cse;
  wire [50:0] stage_PE_gm_im_d_mux_2_cse;
  wire or_658_cse;
  wire and_276_cse;
  wire return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse;
  wire and_281_cse;
  wire or_1997_cse;
  wire and_293_cse;
  wire return_add_generic_AC_RND_CONV_false_7_mux_27_cse;
  wire [49:0] return_extract_21_mux_cse;
  wire and_300_cse;
  wire return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse;
  wire and_307_cse;
  wire and_340_cse;
  wire and_348_cse;
  wire and_356_cse;
  wire and_362_cse;
  wire [10:0] return_extract_32_mux_cse;
  wire return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse;
  wire and_311_cse;
  wire return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse;
  wire and_317_cse;
  wire and_324_cse;
  wire return_add_generic_AC_RND_CONV_false_20_mux_27_cse;
  wire and_328_cse;
  wire and_332_cse;
  wire and_368_cse;
  wire and_374_cse;
  wire and_382_cse;
  wire and_389_cse;
  wire or_87_cse;
  wire or_82_cse;
  wire or_81_cse;
  wire return_extract_51_and_cse;
  wire and_225_cse;
  wire or_32_cse;
  wire nor_34_cse;
  wire nor_35_cse;
  wire and_435_cse;
  wire and_528_cse;
  wire return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_and_cse;
  wire and_606_cse;
  wire and_526_cse;
  wire return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_and_cse;
  wire return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_and_cse;
  wire return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_and_cse;
  wire return_add_generic_AC_RND_CONV_false_19_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_19_op1_smaller_oelse_and_cse;
  reg t_in_10_0_lpi_1_dfm_1_10;
  reg t_in_10_0_lpi_1_dfm_1_9;
  reg BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm;
  reg [50:0] return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm;
  reg drf_qr_lval_15_smx_0_lpi_3_dfm;
  reg [50:0] return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm;
  reg stage_PE_1_tmp_im_d_1_lpi_3_dfm_51;
  reg drf_qr_lval_14_smx_0_lpi_3_dfm;
  reg [50:0] return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm;
  wire return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_10_op2_mu_1_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_10_op2_mu_1_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1;
  reg return_add_generic_AC_RND_CONV_false_23_op1_mu_52_lpi_3_dfm;
  reg [50:0] return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm;
  wire return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1;
  wire stage_PE_tmp_re_d_1_lpi_3_dfm_51_mx0;
  wire return_add_generic_AC_RND_CONV_false_4_op1_mu_52_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_4_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_4_op2_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1;
  reg [8:0] BUTTERFLY_1_n_9_0_sva_8_0;
  wire or_1146_ssc;
  wire or_1147_ssc;
  wire or_1148_ssc;
  wire or_1150_ssc;
  wire or_1174_ssc;
  wire or_1176_ssc;
  wire or_1177_ssc;
  wire or_1179_ssc;
  wire BUTTERFLY_1_i_and_ssc;
  reg reg_BUTTERFLY_1_i_9_0_ftd;
  reg [8:0] reg_BUTTERFLY_1_i_9_0_ftd_1;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_1;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_2;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_3;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_4;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_5;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_6;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_7;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_8;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_9;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_10;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_11;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_12;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_13;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_14;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_15;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_16;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_17;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_18;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_19;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_20;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_21;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_22;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_23;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_24;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_25;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_26;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_27;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_28;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_29;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_30;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_31;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_32;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_33;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_34;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_35;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_36;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_37;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_38;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_39;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_40;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_41;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_42;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_43;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_44;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_45;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_46;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_47;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_48;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_49;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_50;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_51;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_52;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_53;
  wire and_597_m1c;
  reg [2:0] operator_14_false_1_acc_psp_sva_12_10;
  reg [9:0] operator_14_false_1_acc_psp_sva_9_0;
  reg return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_50;
  reg [49:0] return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_49_0;
  wire return_add_generic_AC_RND_CONV_false_18_and_1_ssc;
  reg [5:0] return_add_generic_AC_RND_CONV_false_18_mux_1_itm_55_50;
  reg [49:0] return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0;
  reg [4:0] operator_32_false_1_acc_psp_sva_16_12;
  reg [11:0] operator_32_false_1_acc_psp_sva_11_0;
  wire t_in_or_3_cse;
  wire return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse;
  wire return_add_generic_AC_RND_CONV_false_r_nan_or_cse;
  wire return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_8_op1_smaller_return_add_generic_AC_RND_CONV_false_8_op1_smaller_or_cse;
  wire return_add_generic_AC_RND_CONV_false_21_op1_smaller_return_add_generic_AC_RND_CONV_false_21_op1_smaller_or_cse;
  reg m_in_0_lpi_1_dfm;
  wire [5:0] operator_6_false_17_mux1h_cse_1;
  wire BUTTERFLY_1_fiy_mux1h_4_cse;
  wire BUTTERFLY_1_fiy_mux1h_10_cse;
  wire return_add_generic_AC_RND_CONV_false_10_exp_mux1h_3_cse;
  wire return_add_generic_AC_RND_CONV_false_10_exp_mux1h_6_cse;
  wire return_add_generic_AC_RND_CONV_false_e_dif1_return_add_generic_AC_RND_CONV_false_e_dif1_and_cse;
  wire return_add_generic_AC_RND_CONV_false_13_e_dif1_return_add_generic_AC_RND_CONV_false_13_e_dif1_and_cse;
  wire operator_6_false_17_or_cse;
  wire return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse;
  wire and_1251_cse;
  wire and_1046_cse;
  wire and_1057_cse;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_or_5_cse;
  wire and_2393_rgt;
  wire and_2395_rgt;
  wire and_2407_rgt;
  wire and_2409_rgt;
  wire and_2325_rgt;
  wire and_2327_rgt;
  wire and_2339_rgt;
  wire and_2341_rgt;
  wire BUTTERFLY_if_1_if_or_cse;
  wire or_1302_cse;
  wire return_add_generic_AC_RND_CONV_false_13_or_2_cse;
  wire stage_PE_1_tmp_re_d_or_3_cse;
  wire and_2472_tmp;
  wire or_1122_rmff;
  wire or_1121_rmff;
  wire or_1120_rmff;
  wire or_1119_rmff;
  wire or_1159_ssc;
  wire or_1160_ssc;
  wire or_1132_ssc;
  wire or_1133_ssc;
  reg return_add_generic_AC_RND_CONV_false_11_mux_itm;
  reg return_add_generic_AC_RND_CONV_false_16_mux_itm;
  wire [9:0] return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_11;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1;
  reg [9:0] return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0;
  wire return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w1;
  wire return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_9;
  reg return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs;
  wire return_add_generic_AC_RND_CONV_false_13_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_22_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_23_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_24_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_25_or_1_svs_1;
  wire [9:0] BUTTERFLY_i_9_0_sva_1;
  wire [10:0] nl_BUTTERFLY_i_9_0_sva_1;
  reg [9:0] BUTTERFLY_1_fry_9_0_sva;
  wire [9:0] return_add_generic_AC_RND_CONV_false_1_e_r_qelse_qr_10_1_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_9_exp_plus_1_12_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_1_mux_30;
  reg return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs;
  wire return_add_generic_AC_RND_CONV_false_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_9_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_10_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_11_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_12_or_1_svs_1;
  wire [14:0] stage_monty_mul_acc_2_psp_sva_1;
  wire [15:0] nl_stage_monty_mul_acc_2_psp_sva_1;
  wire BUTTERFLY_1_else_nand_tmp;
  wire and_dcpl_564;
  wire or_tmp;
  wire or_tmp_954;
  wire or_tmp_955;
  wire or_tmp_956;
  wire or_tmp_958;
  wire or_tmp_959;
  wire or_tmp_960;
  wire or_tmp_963;
  wire or_tmp_964;
  wire or_tmp_965;
  wire [50:0] return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_mx1w0;
  reg [10:0] drf_qr_lval_19_smx_lpi_3_dfm;
  reg [9:0] drf_qr_lval_21_smx_9_0_lpi_3_dfm;
  reg [5:0] return_add_generic_AC_RND_CONV_false_11_ls_sva;
  reg [5:0] operator_6_false_17_acc_itm_6_1;
  wire return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_4_e_r_qelse_or_svs_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_5_e_r_qelse_or_svs_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_17_e_r_qelse_or_svs_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_svs_mx0w0;
  wire [11:0] return_add_generic_AC_RND_CONV_false_2_exp_plus_1_12_1_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_3_exp_plus_1_12_1_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_15_exp_plus_1_12_1_lpi_3_dfm_1;
  wire nor_174_m1c;
  wire nor_175_m1c;
  wire nor_177_m1c;
  wire BUTTERFLY_else_or_cse;
  wire BUTTERFLY_if_1_if_and_7_cse;
  wire BUTTERFLY_if_1_if_and_9_cse;
  wire BUTTERFLY_if_1_if_and_6_cse;
  wire BUTTERFLY_if_1_if_and_8_cse;
  wire BUTTERFLY_if_1_if_and_5_cse;
  wire BUTTERFLY_if_1_and_9_cse;
  wire BUTTERFLY_if_1_and_11_cse;
  wire BUTTERFLY_if_1_and_8_cse;
  wire BUTTERFLY_if_1_and_10_cse;
  wire BUTTERFLY_if_1_and_7_cse;
  wire BUTTERFLY_if_1_if_or_2_cse;
  wire BUTTERFLY_if_1_or_2_cse;
  wire [55:0] return_add_generic_AC_RND_CONV_false_12_res_mant_mux1h_1_itm;
  wire [5:0] return_add_generic_AC_RND_CONV_false_2_mux_4_itm;
  wire [5:0] return_add_generic_AC_RND_CONV_false_3_mux_15_itm;
  wire [53:0] return_mult_generic_AC_RND_CONV_false_6_else_1_rshift_itm;
  wire z_out_13;
  wire [17:0] z_out_58;
  wire [18:0] nl_z_out_58;
  wire [15:0] z_out_59;
  wire [16:0] nl_z_out_59;
  wire [15:0] z_out_60;
  wire [17:0] nl_z_out_60;
  wire [16:0] z_out_62;
  wire [5:0] rtn_out;
  wire [16:0] z_out_64;
  wire [17:0] nl_z_out_64;
  wire [53:0] z_out_65;
  wire [9:0] z_out_66;
  wire [10:0] nl_z_out_66;
  wire [9:0] z_out_67;
  wire [10:0] nl_z_out_67;
  wire [12:0] z_out_68;
  wire [11:0] z_out_69;
  wire [11:0] z_out_70;
  wire [56:0] z_out_73;
  wire [56:0] z_out_74;
  wire [56:0] z_out_75;
  wire [56:0] z_out_76;
  wire [56:0] z_out_77;
  wire [56:0] z_out_78;
  wire [56:0] z_out_79;
  wire [56:0] z_out_80;
  wire or_tmp_1400;
  wire [56:0] z_out_81;
  wire all_same_out;
  wire [5:0] rtn_out_1;
  wire all_same_out_1;
  wire [5:0] rtn_out_2;
  wire [17:0] z_out_82;
  wire [18:0] nl_z_out_82;
  wire [12:0] z_out_84;
  wire [13:0] nl_z_out_84;
  wire or_tmp_1439;
  wire or_tmp_1440;
  wire [12:0] z_out_85;
  wire [13:0] nl_z_out_85;
  wire [12:0] z_out_86;
  wire [51:0] z_out_87;
  wire [52:0] nl_z_out_87;
  wire [53:0] z_out_88;
  wire [54:0] nl_z_out_88;
  wire [53:0] z_out_89;
  wire [54:0] nl_z_out_89;
  wire [9:0] z_out_90;
  wire [9:0] z_out_91;
  wire or_tmp_1491;
  wire or_tmp_1492;
  wire [11:0] z_out_94;
  wire [11:0] z_out_95;
  wire [11:0] z_out_96;
  wire [17:0] z_out_98;
  wire [9:0] z_out_101;
  wire [10:0] nl_z_out_101;
  wire [11:0] z_out_102;
  wire [12:0] nl_z_out_102;
  wire [11:0] z_out_103;
  wire [12:0] nl_z_out_103;
  wire [105:0] z_out_104;
  wire [31:0] z_out_105;
  wire signed [32:0] nl_z_out_105;
  wire [105:0] z_out_106;
  wire [54:0] z_out_107;
  wire [54:0] z_out_108;
  wire [54:0] z_out_109;
  wire [54:0] z_out_110;
  wire [16:0] z_out_111;
  wire [10:0] z_out_112;
  wire [11:0] nl_z_out_112;
  wire [10:0] z_out_113;
  wire [11:0] nl_z_out_113;
  wire [11:0] z_out_114;
  wire [12:0] nl_z_out_114;
  reg return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs;
  reg stage_d_mul_return_d_2_63_sva;
  reg return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs;
  reg [5:0] return_add_generic_AC_RND_CONV_false_9_ls_sva;
  reg [56:0] return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva;
  reg return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm;
  reg return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm;
  reg [56:0] return_add_generic_AC_RND_CONV_false_11_res_mant_4_sva;
  reg stage_PE_1_index_const_15_lpi_2_dfm;
  reg stage_PE_1_index_const_10_lpi_2_dfm;
  reg stage_PE_1_index_const_0_lpi_2_dfm;
  reg stage_PE_1_qr_0_lpi_2_dfm;
  reg stage_PE_1_qr_1_0_lpi_2_dfm;
  reg [61:0] stage_PE_1_gm_im_d_61_0_lpi_3_dfm;
  reg return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs;
  reg return_extract_41_return_extract_41_or_1_cse_sva;
  reg return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs;
  reg stage_d_mul_return_d_4_63_sva;
  reg return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs;
  reg [55:0] return_add_generic_AC_RND_CONV_false_11_mux_1_itm;
  reg return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm;
  reg return_add_generic_AC_RND_CONV_false_12_mux_2_itm;
  reg return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_itm;
  reg return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm;
  reg return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_8;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_7;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_8;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_8;
  reg operator_6_false_17_acc_itm_0;
  reg [5:0] operator_6_false_21_acc_itm_6_1;
  reg operator_6_false_21_acc_itm_0;
  wire out1_rsci_idat_63_0_mx0c1;
  wire out1_rsci_idat_63_0_mx0c2;
  wire out1_rsci_idat_79_64_mx0c1;
  wire return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1;
  wire t_in_10_0_lpi_1_dfm_1_10_mx0w0;
  wire mode_lpi_1_dfm_mx0w0;
  wire return_extract_56_m_zero_sva_mx2w0;
  wire [11:0] return_add_generic_AC_RND_CONV_false_6_exp_plus_1_12_1_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_2;
  wire [8:0] BUTTERFLY_i_div_psp_sva_1;
  wire BUTTERFLY_1_i_9_0_sva_mx0c3;
  wire return_add_generic_AC_RND_CONV_false_6_r_nan_and_2;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx8c1;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx8c2;
  wire [10:0] drf_qr_lval_1_smx_lpi_3_dfm_mx0;
  wire return_extract_41_return_extract_41_or_1_cse_sva_1;
  wire return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_1_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_3_res_mant_3_0_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_1_e_dif_sat_sva_1;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm_mx1w0;
  wire return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm_mx1w0;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx1w0;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx3;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx1w0;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx2;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx4;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx2;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx3;
  wire BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx0c8;
  wire return_extract_12_return_extract_12_or_1_cse_sva_1;
  wire return_extract_44_return_extract_44_or_1_cse_sva_1;
  wire [10:0] drf_qr_lval_10_smx_lpi_3_dfm_mx2;
  wire [10:0] drf_qr_lval_10_smx_lpi_3_dfm_mx6;
  wire return_add_generic_AC_RND_CONV_false_8_if_2_return_add_generic_AC_RND_CONV_false_8_if_2_and_1_mx2w0;
  wire return_add_generic_AC_RND_CONV_false_7_if_2_return_add_generic_AC_RND_CONV_false_7_if_2_and_1_mx4w0;
  wire return_add_generic_AC_RND_CONV_false_12_if_2_return_add_generic_AC_RND_CONV_false_12_if_2_nor_mx3w0;
  wire return_add_generic_AC_RND_CONV_false_11_if_2_return_add_generic_AC_RND_CONV_false_11_if_2_nor_mx5w0;
  wire return_add_generic_AC_RND_CONV_false_6_do_sub_sva_1;
  wire return_add_generic_AC_RND_CONV_false_19_do_sub_sva_1;
  wire return_add_generic_AC_RND_CONV_false_1_if_2_return_add_generic_AC_RND_CONV_false_1_if_2_and_1_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_10_if_2_return_add_generic_AC_RND_CONV_false_10_if_2_and_1_mx3w0;
  wire return_add_generic_AC_RND_CONV_false_13_if_2_return_add_generic_AC_RND_CONV_false_13_if_2_and_1_mx4w1;
  wire return_add_generic_AC_RND_CONV_false_9_if_2_return_add_generic_AC_RND_CONV_false_9_if_2_and_1_mx5w0;
  wire [5:0] return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_24_e_dif_sat_sva_1;
  wire [16:0] stage_u_add_acc_1_itm_1;
  wire [17:0] nl_stage_u_add_acc_1_itm_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm_mx1w0;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_mx1c2;
  wire return_add_generic_AC_RND_CONV_false_4_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_5_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_6_r_nan_or_mx6w0;
  wire return_add_generic_AC_RND_CONV_false_14_op1_nan_sva_mx0w5;
  wire return_add_generic_AC_RND_CONV_false_10_op1_nan_sva_mx0w9;
  wire [11:0] operator_6_false_7_acc_psp_sva_mx0w0;
  wire [12:0] nl_operator_6_false_7_acc_psp_sva_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_18_mux_1_itm_mx1c2;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_res_mant_3_0_sva_1;
  wire [51:0] return_add_generic_AC_RND_CONV_false_res_rounded_lpi_3_dfm_51_0_1;
  wire return_add_generic_AC_RND_CONV_false_2_res_mant_3_0_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_e_dif_sat_sva_1;
  wire return_add_generic_AC_RND_CONV_false_6_exp_plus_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_19_exp_plus_1_0_lpi_3_dfm_1;
  wire [51:0] return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1;
  wire return_add_generic_AC_RND_CONV_false_2_exp_plus_1_0_lpi_3_dfm_1;
  wire [10:0] operator_6_false_9_acc_psp_1_sva_1;
  wire [11:0] nl_operator_6_false_9_acc_psp_1_sva_1;
  wire return_add_generic_AC_RND_CONV_false_3_exp_plus_1_0_lpi_3_dfm_1;
  wire [10:0] operator_6_false_11_acc_psp_1_sva_1;
  wire [11:0] nl_operator_6_false_11_acc_psp_1_sva_1;
  wire return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_50_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0;
  wire return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_6_op1_smaller_lor_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_6_res_mant_3_0_sva_1;
  wire return_extract_15_return_extract_15_or_sva_1;
  wire return_add_generic_AC_RND_CONV_false_4_m_r_51_lpi_3_dfm_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_4_e_r_qr_10_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1;
  wire [11:0] operator_6_false_13_acc_psp_sva_1;
  wire [12:0] nl_operator_6_false_13_acc_psp_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_6_e_dif_sat_sva_1;
  wire return_add_generic_AC_RND_CONV_false_4_if_7_not_4;
  wire [11:0] return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_2_10_0_1;
  wire return_mult_generic_AC_RND_CONV_false_1_e_incr_lpi_3_dfm_2;
  wire return_extract_17_return_extract_17_or_sva_1;
  wire return_add_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_5_e_r_qr_10_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_if_1_and_1_tmp_1;
  wire return_add_generic_AC_RND_CONV_false_5_if_7_not_4;
  wire [9:0] return_add_generic_AC_RND_CONV_false_6_e_r_qelse_qr_10_1_lpi_3_dfm_1;
  wire return_extract_19_return_extract_19_or_sva_1;
  wire return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_tmp_1;
  wire return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_7_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_8_res_mant_3_0_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_2_if_1_and_1_tmp_1;
  wire [49:0] return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_9_res_mant_3_0_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_8_mux_20_mx0;
  wire [9:0] return_add_generic_AC_RND_CONV_false_8_e_r_qelse_qr_10_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_8_r_nan_or_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_10_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_12_res_mant_3_0_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_1;
  wire return_add_generic_AC_RND_CONV_false_11_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_14_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_16_res_mant_3_0_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_16_e_dif_sat_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_14_e_dif_sat_sva_1;
  wire return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_13_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_15_res_mant_3_0_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_15_e_dif_sat_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_13_e_dif_sat_sva_1;
  wire [17:0] operator_32_false_3_acc_psp_sva_1;
  wire [18:0] nl_operator_32_false_3_acc_psp_sva_1;
  wire return_add_generic_AC_RND_CONV_false_15_exp_plus_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_16_exp_plus_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_50_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0;
  wire return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_19_op1_smaller_lor_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_19_res_mant_3_0_sva_1;
  wire return_extract_47_return_extract_47_or_sva_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm_1;
  wire [11:0] operator_6_false_42_acc_psp_sva_1;
  wire [12:0] nl_operator_6_false_42_acc_psp_sva_1;
  wire return_extract_49_return_extract_49_or_sva_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_18_e_r_qr_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_3_if_1_and_1_tmp_1;
  wire return_extract_51_return_extract_51_or_sva_1;
  wire return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_4_if_1_and_1_tmp_1;
  wire return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_20_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_21_res_mant_3_0_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_5_if_1_and_1_tmp_1;
  wire return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_22_res_mant_3_0_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_22_e_dif_sat_sva_1;
  wire return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_23_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_25_res_mant_3_0_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_23_e_dif_sat_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1;
  wire [52:0] return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_6_if_1_and_1_tmp_1;
  wire [14:0] operator_32_false_2_acc_psp_1_sva_1;
  wire [15:0] nl_operator_32_false_2_acc_psp_1_sva_1;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_else_2_else_else_mux_2;
  wire return_add_generic_AC_RND_CONV_false_4_sticky_bit_and_158;
  wire return_add_generic_AC_RND_CONV_false_6_mux_36;
  wire return_add_generic_AC_RND_CONV_false_3_return_add_generic_AC_RND_CONV_false_3_and_9;
  reg return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_56;
  reg m_in_15_1_lpi_1_dfm_1_0;
  reg return_add_generic_AC_RND_CONV_false_18_op_bigger_mux_1_itm_50;
  reg [49:0] return_add_generic_AC_RND_CONV_false_18_op_bigger_mux_1_itm_49_0;
  wire drf_qr_lval_6_smx_lpi_3_dfm_mx0_0;
  wire drf_qr_lval_22_smx_lpi_3_dfm_mx0_0;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_0;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_0;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_0;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_0;
  wire leading_sign_57_0_1_0_19_out_2;
  wire [5:0] leading_sign_57_0_1_0_19_out_3;
  wire [5:0] leading_sign_53_0_6_out_1;
  wire [55:0] return_add_generic_AC_RND_CONV_false_6_res_mant_conc_2_itm_56_1;
  wire [55:0] return_add_generic_AC_RND_CONV_false_19_res_mant_conc_2_itm_56_1;
  reg [4:0] BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0;
  reg drf_qr_lval_10_smx_lpi_3_dfm_rsp_0;
  wire return_add_generic_AC_RND_CONV_false_7_exp_and_ssc;
  reg [3:0] return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_0;
  reg [51:0] return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1;
  wire return_add_generic_AC_RND_CONV_false_12_res_mant_and_1_ssc;
  wire or_1864_ssc;
  wire or_1866_ssc;
  wire drf_qr_lval_6_smx_lpi_3_dfm_mx0_10;
  wire [8:0] drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_1;
  wire drf_qr_lval_22_smx_lpi_3_dfm_mx0_10;
  wire [8:0] drf_qr_lval_22_smx_lpi_3_dfm_mx0_9_1;
  wire operator_6_false_3_or_1_ssc;
  wire return_add_generic_AC_RND_CONV_false_19_exp_plus_1_and_cse;
  wire return_add_generic_AC_RND_CONV_false_12_op_bigger_and_cse;
  wire stage_PE_1_tmp_re_d_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_2_if_5_return_add_generic_AC_RND_CONV_false_2_if_5_nor_cse;
  wire [11:0] return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_2_cse;
  wire [9:0] nor_182_cse;
  wire [9:0] nor_186_cse;
  wire return_add_generic_AC_RND_CONV_false_11_or_4_cse;
  wire BUTTERFLY_1_i_or_3_cse;
  wire BUTTERFLY_else_1_or_cse;
  wire or_1341_cse;
  wire return_add_generic_AC_RND_CONV_false_11_or_5_cse;
  wire or_2455_cse;
  wire [55:0] return_add_generic_AC_RND_CONV_false_9_mux_28_cse;
  wire [55:0] return_add_generic_AC_RND_CONV_false_7_mux_31_cse;
  wire [55:0] return_add_generic_AC_RND_CONV_false_10_mux_28_cse;
  wire return_mult_generic_AC_RND_CONV_false_mux1h_cse;
  wire return_mult_generic_AC_RND_CONV_false_mux1h_1_cse;
  wire return_add_generic_AC_RND_CONV_false_e_dif1_or_1_cse;
  wire return_add_generic_AC_RND_CONV_false_1_res_rounded_or_2_cse;
  wire return_add_generic_AC_RND_CONV_false_7_res_rounded_and_cse;
  wire [5:0] return_add_generic_AC_RND_CONV_false_7_mux_33_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse;
  wire return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse;
  wire return_add_generic_AC_RND_CONV_false_10_r_zero_or_2_cse;
  wire return_add_generic_AC_RND_CONV_false_10_ls_or_2_cse;
  wire nand_133_cse;
  wire return_mult_generic_AC_RND_CONV_false_if_or_3_cse;
  wire [3:0] return_mult_generic_AC_RND_CONV_false_if_nand_1_cse;
  wire return_mult_generic_AC_RND_CONV_false_if_or_cse;
  wire return_add_generic_AC_RND_CONV_false_3_if_5_nor_cse;
  wire [5:0] return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_cse;
  wire return_mult_generic_AC_RND_CONV_false_2_if_or_3_cse;
  wire [3:0] return_mult_generic_AC_RND_CONV_false_2_if_nand_1_cse;
  wire return_mult_generic_AC_RND_CONV_false_2_if_or_cse;
  wire [5:0] return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse;
  wire and_3379_cse;
  wire return_add_generic_AC_RND_CONV_false_12_or_9_cse;
  wire operator_6_false_33_or_5_cse;
  wire operator_6_false_33_or_7_cse;
  wire operator_6_false_33_or_1_cse;
  wire operator_6_false_33_or_3_cse;
  wire operator_6_false_3_or_6_cse;
  wire operator_6_false_3_or_8_cse;
  wire operator_6_false_3_or_2_cse;
  wire operator_6_false_3_or_4_cse;
  wire return_add_generic_AC_RND_CONV_false_6_e_dif1_or_1_cse;
  wire BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_4_cse;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_or_cse;
  wire return_add_generic_AC_RND_CONV_false_12_or_22_cse;
  wire operator_6_false_33_or_12_cse;
  wire operator_6_false_33_or_14_cse;
  wire operator_6_false_33_or_15_cse;
  wire operator_6_false_3_or_12_cse;
  wire nand_102_cse;
  wire return_add_generic_AC_RND_CONV_false_10_r_zero_or_3_cse;
  wire return_extract_22_or_2_cse;
  wire return_add_generic_AC_RND_CONV_false_21_r_sign_mux_1_cse;
  wire return_add_generic_AC_RND_CONV_false_8_r_sign_mux_1_cse;
  wire and_275_cse;
  wire return_add_generic_AC_RND_CONV_false_12_r_zero_or_1_cse;
  wire and_339_cse;
  wire return_add_generic_AC_RND_CONV_false_12_or_11_cse_1;
  wire return_add_generic_AC_RND_CONV_false_12_or_41_cse;
  wire return_add_generic_AC_RND_CONV_false_3_or_4_cse;
  wire operator_14_false_1_or_cse;
  wire return_add_generic_AC_RND_CONV_false_2_and_cse;
  wire return_add_generic_AC_RND_CONV_false_2_and_6_cse;
  wire return_add_generic_AC_RND_CONV_false_2_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_2_and_2_cse;
  wire return_add_generic_AC_RND_CONV_false_2_and_8_cse;
  wire return_add_generic_AC_RND_CONV_false_2_or_5_cse;
  wire return_add_generic_AC_RND_CONV_false_2_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_2_and_10_cse;
  wire return_add_generic_AC_RND_CONV_false_2_or_7_cse;
  wire return_add_generic_AC_RND_CONV_false_1_and_16_cse;
  wire return_add_generic_AC_RND_CONV_false_1_and_20_cse;
  wire return_add_generic_AC_RND_CONV_false_1_or_7_cse;
  wire return_add_generic_AC_RND_CONV_false_1_or_9_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_33_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_39_cse;
  wire return_add_generic_AC_RND_CONV_false_12_or_24_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_29_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_31_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_35_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_37_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_30_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_32_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_36_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_38_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_25_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_27_cse;
  wire and_2172_cse;
  wire and_2173_cse;
  wire return_add_generic_AC_RND_CONV_false_1_or_6_cse;
  wire return_add_generic_AC_RND_CONV_false_12_or_27_cse;
  wire return_add_generic_AC_RND_CONV_false_12_or_29_cse;
  wire return_add_generic_AC_RND_CONV_false_12_or_44_cse;
  wire return_add_generic_AC_RND_CONV_false_10_ls_or_cse;
  wire return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_ssc;
  reg [4:0] return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_5_1;
  reg return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_0;
  reg m_in_15_1_lpi_1_dfm_1_1;
  wire return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_4_cse;
  wire return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_6_cse;
  wire and_517_tmp;
  wire return_extract_33_or_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_17_and_2_m1c;
  wire return_add_generic_AC_RND_CONV_false_12_and_106_m1c;
  wire return_add_generic_AC_RND_CONV_false_12_and_108_m1c;
  wire return_add_generic_AC_RND_CONV_false_12_and_114_m1c;
  wire and_572_tmp;
  wire and_577_tmp;
  wire and_582_tmp;
  wire and_584_tmp;
  wire and_588_tmp;
  wire and_591_tmp;
  wire return_add_generic_AC_RND_CONV_false_11_and_12_m1c;
  wire return_add_generic_AC_RND_CONV_false_11_and_14_m1c;
  wire return_add_generic_AC_RND_CONV_false_11_and_16_m1c;
  wire return_add_generic_AC_RND_CONV_false_16_and_2_m1c;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_1;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_1;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_1;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_1;
  reg m_in_15_1_lpi_1_dfm_1_2;
  wire return_add_generic_AC_RND_CONV_false_17_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_13_or_cse;
  wire return_add_generic_AC_RND_CONV_false_13_or_3_cse;
  wire return_add_generic_AC_RND_CONV_false_10_res_rounded_and_cse;
  wire return_extract_41_and_1_cse;
  wire operator_6_false_17_or_8_cse;
  wire operator_6_false_7_or_rgt;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_2;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_2;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_2;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_2;
  reg m_in_15_1_lpi_1_dfm_1_3;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_7_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_8_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_9_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_10_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse;
  wire return_add_generic_AC_RND_CONV_false_18_exp_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_18_exp_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_18_exp_or_cse;
  wire return_add_generic_AC_RND_CONV_false_18_exp_and_6_cse;
  wire return_add_generic_AC_RND_CONV_false_17_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_17_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_105_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_111_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_107_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_112_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_109_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_110_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_113_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_13_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_13_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_11_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_13_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_15_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_32_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_10_cse;
  wire return_add_generic_AC_RND_CONV_false_18_exp_and_4_cse;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_3;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_3;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_3;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_3;
  reg m_in_15_1_lpi_1_dfm_1_4;
  wire t_in_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_115_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_117_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_116_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_118_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_119_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_120_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_95_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_103_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_96_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_104_cse;
  wire return_add_generic_AC_RND_CONV_false_13_and_2_cse;
  wire return_add_generic_AC_RND_CONV_false_13_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_13_or_4_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_19_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_21_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_17_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_18_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_20_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_22_cse;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_4;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_4;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_4;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_4;
  reg m_in_15_1_lpi_1_dfm_1_5;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_5;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_5;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_6;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_5;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_5;
  reg m_in_15_1_lpi_1_dfm_1_6;
  reg t_in_10_0_lpi_1_dfm_1_8;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_7;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_6;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_6;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_7;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_6;
  reg m_in_15_1_lpi_1_dfm_1_7;
  reg t_in_10_0_lpi_1_dfm_1_7;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_7;
  reg t_in_10_0_lpi_1_dfm_1_6;
  reg m_in_15_1_lpi_1_dfm_1_8;
  reg t_in_10_0_lpi_1_dfm_1_5;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_8;
  reg t_in_10_0_lpi_1_dfm_1_4;
  reg m_in_15_1_lpi_1_dfm_1_9;
  reg t_in_10_0_lpi_1_dfm_1_3;
  reg t_in_10_0_lpi_1_dfm_1_2;
  reg m_in_15_1_lpi_1_dfm_1_10;
  reg t_in_10_0_lpi_1_dfm_1_1;
  reg t_in_10_0_lpi_1_dfm_1_0;
  reg stage_PE_1_index_const_14_11_lpi_2_dfm_0;
  reg m_in_15_1_lpi_1_dfm_1_11;
  reg stage_PE_1_index_const_14_11_lpi_2_dfm_1;
  reg m_in_15_1_lpi_1_dfm_1_12;
  reg stage_PE_1_index_const_14_11_lpi_2_dfm_3;
  reg stage_PE_1_index_const_14_11_lpi_2_dfm_2;
  reg m_in_15_1_lpi_1_dfm_1_14;
  reg m_in_15_1_lpi_1_dfm_1_13;
  wire or_2748_cse;
  wire [50:0] return_extract_2_mux_4_cse;
  wire [50:0] return_extract_33_mux_3_cse;
  wire return_add_generic_AC_RND_CONV_false_18_exp_and_2_itm;
  wire return_add_generic_AC_RND_CONV_false_11_and_9_itm;
  wire or_1342_itm;
  wire or_2707_itm;
  wire [10:0] operator_32_false_2_acc_5_itm;
  wire [11:0] nl_operator_32_false_2_acc_5_itm;
  wire return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_1_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_9_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_10_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_12_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_14_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_13_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_19_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_22_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_itm_52;
  wire return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1;
  wire return_add_generic_AC_RND_CONV_false_17_acc_3_itm_10;
  wire return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_16_acc_3_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1;
  reg BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0;
  reg [9:0] BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1;
  wire and_3925_ssc;
  reg [8:0] drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0;
  reg drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1;
  wire return_add_generic_AC_RND_CONV_false_7_exp_and_2_ssc;
  wire [9:0] return_add_generic_AC_RND_CONV_false_7_exp_mux1h_4_itm_9_0;
  wire [4:0] return_add_generic_AC_RND_CONV_false_15_mux_4_itm_5_1;
  wire [4:0] return_add_generic_AC_RND_CONV_false_7_mux_24_mx0_5_1;
  wire [8:0] BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_1_9_1;
  wire BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_1_0;
  wire return_add_generic_AC_RND_CONV_false_12_return_add_generic_AC_RND_CONV_false_12_nor_1_ssc;
  wire return_add_generic_AC_RND_CONV_false_12_or_16_ssc;
  wire return_add_generic_AC_RND_CONV_false_12_and_6_ssc;
  wire return_add_generic_AC_RND_CONV_false_2_or_4_ssc;
  wire return_add_generic_AC_RND_CONV_false_2_or_6_ssc;
  wire return_add_generic_AC_RND_CONV_false_3_or_2_seb;
  wire return_add_generic_AC_RND_CONV_false_12_and_89_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_90_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_91_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_92_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_97_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_98_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_99_cse;
  wire return_add_generic_AC_RND_CONV_false_12_and_100_cse;
  wire BUTTERFLY_1_else_1_if_and_1_rgt;
  wire BUTTERFLY_1_else_1_if_or_rgt;
  wire z_out_53_52;
  wire z_out_54_52;
  wire z_out_57_52;
  wire [15:0] z_out_61_15_0;
  wire [16:0] nl_z_out_61_15_0;
  wire z_out_71_11;
  wire return_add_generic_AC_RND_CONV_false_4_or_8_tmp;
  wire [5:0] acc_18_cse_6_1;
  wire [6:0] nl_acc_18_cse_6_1;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_or_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_6_else_2_else_return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_6_else_2_else_mux_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl;
  wire BUTTERFLY_if_1_and_nl;
  wire BUTTERFLY_if_1_and_1_nl;
  wire[50:0] return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_oelse_3_not_1_nl;
  wire t_in_mux_nl;
  wire t_in_mux_2_nl;
  wire t_in_mux_3_nl;
  wire t_in_mux_4_nl;
  wire t_in_mux_5_nl;
  wire t_in_mux_6_nl;
  wire t_in_mux_7_nl;
  wire t_in_mux_8_nl;
  wire t_in_mux_9_nl;
  wire need_ovf_1_need_ovf_1_and_nl;
  wire need_ovf_1_need_ovf_1_and_1_nl;
  wire m_in_mux_nl;
  wire m_in_mux_14_nl;
  wire m_in_mux_13_nl;
  wire m_in_mux_12_nl;
  wire m_in_mux_11_nl;
  wire m_in_mux_10_nl;
  wire m_in_mux_9_nl;
  wire m_in_mux_8_nl;
  wire m_in_mux_7_nl;
  wire m_in_mux_6_nl;
  wire m_in_mux_5_nl;
  wire m_in_mux_4_nl;
  wire m_in_mux_3_nl;
  wire m_in_mux_2_nl;
  wire not_932_nl;
  wire and_994_nl;
  wire and_996_nl;
  wire stage_PE_qif_qelse_mux_nl;
  wire stage_PE_qif_qelse_mux_1_nl;
  wire stage_PE_qif_qelse_mux_14_nl;
  wire stage_PE_qif_qelse_mux_13_nl;
  wire stage_PE_qif_qelse_mux_12_nl;
  wire stage_PE_qif_qelse_mux_11_nl;
  wire[9:0] or_2026_nl;
  wire[9:0] and_2618_nl;
  wire[9:0] mux1h_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_3_return_add_generic_AC_RND_CONV_false_3_and_6_nl;
  wire or_2741_nl;
  wire and_2611_nl;
  wire or_2742_nl;
  wire BUTTERFLY_else_and_2_nl;
  wire or_2744_nl;
  wire and_2613_nl;
  wire and_2614_nl;
  wire BUTTERFLY_else_and_4_nl;
  wire and_2616_nl;
  wire and_2617_nl;
  wire nand_153_nl;
  wire and_1068_nl;
  wire BUTTERFLY_i_or_nl;
  wire return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_3_nl;
  wire return_extract_12_m_zero_return_extract_12_m_zero_nor_nl;
  wire return_extract_20_m_zero_return_extract_20_m_zero_nor_nl;
  wire return_extract_25_m_zero_return_extract_25_m_zero_nor_nl;
  wire return_extract_53_m_zero_return_extract_53_m_zero_nor_nl;
  wire return_extract_59_m_zero_return_extract_59_m_zero_nor_nl;
  wire operator_11_true_12_operator_11_true_12_and_nl;
  wire operator_11_true_52_operator_11_true_52_and_nl;
  wire operator_11_true_25_operator_11_true_25_and_nl;
  wire operator_11_true_44_operator_11_true_44_and_nl;
  wire operator_11_true_57_operator_11_true_57_and_nl;
  wire return_add_generic_AC_RND_CONV_false_25_r_nan_and_nl;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_or_6_nl;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_and_3_nl;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_or_8_nl;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_and_4_nl;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_and_5_nl;
  wire reg_return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_rgt_nl;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_or_3_nl;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_or_4_nl;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_18_exp_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_6_nl;
  wire return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_21_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_22_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_16_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_93_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_94_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_101_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_102_nl;
  wire return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_3_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_or_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_4_if_2_return_add_generic_AC_RND_CONV_false_4_if_2_nor_1_nl;
  wire or_756_nl;
  wire or_1538_nl;
  wire return_add_generic_AC_RND_CONV_false_5_if_2_return_add_generic_AC_RND_CONV_false_5_if_2_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_9_do_sub_return_add_generic_AC_RND_CONV_false_9_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_23_do_sub_return_add_generic_AC_RND_CONV_false_23_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_3_if_2_return_add_generic_AC_RND_CONV_false_3_if_2_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_15_if_2_return_add_generic_AC_RND_CONV_false_15_if_2_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_46_nl;
  wire return_add_generic_AC_RND_CONV_false_17_do_sub_return_add_generic_AC_RND_CONV_false_17_do_sub_return_add_generic_AC_RND_CONV_false_17_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_10_do_sub_return_add_generic_AC_RND_CONV_false_10_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_22_do_sub_return_add_generic_AC_RND_CONV_false_22_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_18_do_sub_return_add_generic_AC_RND_CONV_false_18_do_sub_xor_nl;
  wire return_mult_generic_AC_RND_CONV_false_r_nan_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_r_nan_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_11_r_nan_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_r_nan_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_r_nan_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_24_r_nan_and_nl;
  wire return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_8_do_sub_return_add_generic_AC_RND_CONV_false_8_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_21_do_sub_return_add_generic_AC_RND_CONV_false_21_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_10_r_zero_or_1_nl;
  wire return_extract_50_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_zero_m_return_mult_generic_AC_RND_CONV_false_2_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_2_r_zero_return_mult_generic_AC_RND_CONV_false_2_r_zero_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_zero_m_return_mult_generic_AC_RND_CONV_false_5_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_5_r_zero_return_mult_generic_AC_RND_CONV_false_5_r_zero_nor_nl;
  wire operator_11_true_53_operator_11_true_53_and_nl;
  wire operator_11_true_27_operator_11_true_27_and_nl;
  wire operator_11_true_59_operator_11_true_59_and_nl;
  wire return_extract_24_exception_or_1_nl;
  wire return_extract_21_m_zero_return_extract_21_m_zero_nor_nl;
  wire return_extract_27_m_zero_return_extract_27_m_zero_nor_nl;
  wire return_extract_44_m_zero_return_extract_44_m_zero_nor_nl;
  wire return_extract_52_m_zero_return_extract_52_m_zero_nor_nl;
  wire return_extract_57_m_zero_return_extract_57_m_zero_nor_nl;
  wire operator_33_true_12_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_5_e_dif_sat_or_2_nl;
  wire operator_6_false_17_and_2_nl;
  wire operator_6_false_17_or_9_nl;
  wire return_add_generic_AC_RND_CONV_false_10_ls_or_6_nl;
  wire operator_32_false_1_or_1_nl;
  wire operator_32_false_1_operator_32_false_1_nor_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_14_mux1h_11_nl;
  wire return_add_generic_AC_RND_CONV_false_14_or_5_nl;
  wire nor_245_nl;
  wire return_extract_22_or_nl;
  wire return_extract_22_or_1_nl;
  wire mux_24_nl;
  wire mux_23_nl;
  wire and_38_nl;
  wire or_70_nl;
  wire return_add_generic_AC_RND_CONV_false_11_or_nl;
  wire return_add_generic_AC_RND_CONV_false_11_or_6_nl;
  wire return_add_generic_AC_RND_CONV_false_11_or_7_nl;
  wire return_add_generic_AC_RND_CONV_false_11_or_8_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_18_ma1_lt_ma2_acc_2_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_18_ma1_lt_ma2_acc_2_nl;
  wire and_1245_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_1_r_nan_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_2_r_nan_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_3_r_nan_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_or_nl;
  wire return_add_generic_AC_RND_CONV_false_16_r_nan_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_11_exp_or_nl;
  wire return_add_generic_AC_RND_CONV_false_11_exp_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_11_exp_and_3_nl;
  wire return_add_generic_AC_RND_CONV_false_11_exp_or_3_nl;
  wire return_add_generic_AC_RND_CONV_false_11_exp_and_5_nl;
  wire return_add_generic_AC_RND_CONV_false_11_exp_or_4_nl;
  wire return_add_generic_AC_RND_CONV_false_11_exp_and_9_nl;
  wire return_add_generic_AC_RND_CONV_false_11_exp_and_11_nl;
  wire return_add_generic_AC_RND_CONV_false_12_exp_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_12_exp_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_r_return_add_generic_AC_RND_CONV_false_1_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_nl;
  wire or_352_nl;
  wire return_add_generic_AC_RND_CONV_false_2_e_r_return_add_generic_AC_RND_CONV_false_2_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_2_mux_13_nl;
  wire return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_1_nl;
  wire or_370_nl;
  wire return_add_generic_AC_RND_CONV_false_3_e_r_return_add_generic_AC_RND_CONV_false_3_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux_13_nl;
  wire return_add_generic_AC_RND_CONV_false_16_e_r_qelse_mux_1_nl;
  wire or_382_nl;
  wire return_add_generic_AC_RND_CONV_false_6_if_5_return_add_generic_AC_RND_CONV_false_6_if_5_and_nl;
  wire return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_4_nl;
  wire or_409_nl;
  wire return_add_generic_AC_RND_CONV_false_15_e_r_return_add_generic_AC_RND_CONV_false_15_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_15_mux_13_nl;
  wire return_add_generic_AC_RND_CONV_false_15_return_add_generic_AC_RND_CONV_false_15_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_15_e_r_qelse_mux_1_nl;
  wire or_426_nl;
  wire return_add_generic_AC_RND_CONV_false_16_e_r_return_add_generic_AC_RND_CONV_false_16_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_16_mux_13_nl;
  wire return_add_generic_AC_RND_CONV_false_16_e_r_qelse_mux_3_nl;
  wire or_434_nl;
  wire return_add_generic_AC_RND_CONV_false_19_if_5_return_add_generic_AC_RND_CONV_false_19_if_5_and_nl;
  wire return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_16_r_zero_or_nl;
  wire operator_11_true_54_operator_11_true_54_and_nl;
  wire return_extract_58_and_1_nl;
  wire or_1826_nl;
  wire return_add_generic_AC_RND_CONV_false_18_return_add_generic_AC_RND_CONV_false_18_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_18_and_9_nl;
  wire return_add_generic_AC_RND_CONV_false_6_or_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl;
  wire return_add_generic_AC_RND_CONV_false_2_if_2_return_add_generic_AC_RND_CONV_false_2_if_2_nor_1_nl;
  wire and_596_nl;
  wire return_add_generic_AC_RND_CONV_false_2_if_2_and_nl;
  wire return_add_generic_AC_RND_CONV_false_2_if_2_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_11_or_9_nl;
  wire return_add_generic_AC_RND_CONV_false_16_if_2_return_add_generic_AC_RND_CONV_false_16_if_2_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_16_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_16_and_9_nl;
  wire return_add_generic_AC_RND_CONV_false_16_or_nl;
  wire return_add_generic_AC_RND_CONV_false_7_do_sub_return_add_generic_AC_RND_CONV_false_7_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_20_do_sub_return_add_generic_AC_RND_CONV_false_20_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_or_1_nl;
  wire return_extract_56_and_1_nl;
  wire stage_PE_1_tmp_re_d_and_3_nl;
  wire stage_PE_1_tmp_re_d_and_4_nl;
  wire stage_PE_1_tmp_re_d_and_5_nl;
  wire stage_PE_1_tmp_re_d_and_6_nl;
  wire return_add_generic_AC_RND_CONV_false_2_mux_9_nl;
  wire return_add_generic_AC_RND_CONV_false_2_if_5_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_3_if_5_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_6_mux_33_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux_15_nl;
  wire return_add_generic_AC_RND_CONV_false_4_if_5_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_5_mux_9_nl;
  wire return_add_generic_AC_RND_CONV_false_5_if_5_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_15_mux_9_nl;
  wire return_add_generic_AC_RND_CONV_false_15_if_5_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_17_mux_15_nl;
  wire return_add_generic_AC_RND_CONV_false_17_if_5_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_18_mux_9_nl;
  wire return_add_generic_AC_RND_CONV_false_18_if_5_or_1_nl;
  wire[11:0] return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl;
  wire[12:0] nl_return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl;
  wire[11:0] operator_33_true_13_acc_nl;
  wire[12:0] nl_operator_33_true_13_acc_nl;
  wire[11:0] operator_33_true_39_acc_nl;
  wire[12:0] nl_operator_33_true_39_acc_nl;
  wire[8:0] return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_8_nl;
  wire return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_9_nl;
  wire return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif_sat_or_1_nl;
  wire and_543_nl;
  wire and_548_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_1_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_1_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_6_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_6_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_9_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_9_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_10_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_10_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_11_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_11_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_12_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_12_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_14_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_14_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_13_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_13_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_19_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_19_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_22_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_22_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_23_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_23_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_24_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_24_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_25_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_25_acc_2_nl;
  wire[53:0] acc_3_nl;
  wire[54:0] nl_acc_3_nl;
  wire return_add_generic_AC_RND_CONV_false_8_ma1_lt_ma2_mux_5_nl;
  wire nand_128_nl;
  wire[53:0] acc_2_nl;
  wire[54:0] nl_acc_2_nl;
  wire return_add_generic_AC_RND_CONV_false_21_ma1_lt_ma2_mux_5_nl;
  wire nand_129_nl;
  wire nand_130_nl;
  wire nand_131_nl;
  wire[5:0] operator_6_false_41_acc_nl;
  wire[6:0] nl_operator_6_false_41_acc_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_24_e_dif_sat_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_oelse_3_return_mult_generic_AC_RND_CONV_false_3_if_3_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_oelse_3_return_mult_generic_AC_RND_CONV_false_4_if_3_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_r_qelse_not_5_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_1_if_5_or_nl;
  wire and_592_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_e_dif_acc_1_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_e_dif_acc_1_nl;
  wire return_add_generic_AC_RND_CONV_false_not_3_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_2_not_3_nl;
  wire return_add_generic_AC_RND_CONV_false_2_mux_14_nl;
  wire return_add_generic_AC_RND_CONV_false_2_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux_14_nl;
  wire return_add_generic_AC_RND_CONV_false_3_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_6_mux_6_nl;
  wire return_add_generic_AC_RND_CONV_false_6_r_sign_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_and_nl;
  wire return_add_generic_AC_RND_CONV_false_19_mux_6_nl;
  wire return_add_generic_AC_RND_CONV_false_19_r_sign_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_and_nl;
  wire nor_179_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux_19_nl;
  wire return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_3_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_dif_sat_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_not_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_if_not_1_nl;
  wire nor_183_nl;
  wire return_add_generic_AC_RND_CONV_false_5_mux_13_nl;
  wire return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_2_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_6_mux_31_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_not_3_nl;
  wire and_600_nl;
  wire return_add_generic_AC_RND_CONV_false_6_if_7_return_add_generic_AC_RND_CONV_false_6_if_7_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_19_e_r_qelse_mux_nl;
  wire or_389_nl;
  wire return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_3_nl;
  wire return_add_generic_AC_RND_CONV_false_6_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_6_if_5_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_if_not_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_7_e_dif_qif_acc_1_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_7_e_dif_qif_acc_1_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_2_else_2_else_return_mult_generic_AC_RND_CONV_false_2_else_2_else_and_nl;
  wire and_602_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_oelse_3_return_mult_generic_AC_RND_CONV_false_5_if_3_nor_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_8_e_dif_qif_acc_1_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_8_e_dif_qif_acc_1_nl;
  wire return_add_generic_AC_RND_CONV_false_8_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_7_e_dif_sat_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_3_nl;
  wire or_396_nl;
  wire return_add_generic_AC_RND_CONV_false_7_if_7_return_add_generic_AC_RND_CONV_false_7_if_7_nor_nl;
  wire return_extract_25_return_extract_25_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_18_nl;
  wire return_add_generic_AC_RND_CONV_false_7_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_8_e_r_qelse_not_5_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_nl;
  wire or_404_nl;
  wire and_609_nl;
  wire return_add_generic_AC_RND_CONV_false_8_if_7_return_add_generic_AC_RND_CONV_false_8_if_7_nor_nl;
  wire return_extract_27_return_extract_27_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_10_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_8_mux_14_nl;
  wire return_add_generic_AC_RND_CONV_false_8_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_9_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_9_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_10_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_10_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_11_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_11_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_12_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_12_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_16_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_14_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_14_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_14_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_13_e_dif_sat_or_1_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl;
  wire return_add_generic_AC_RND_CONV_false_13_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_13_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_15_mux_14_nl;
  wire return_add_generic_AC_RND_CONV_false_15_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_16_mux_14_nl;
  wire return_add_generic_AC_RND_CONV_false_16_if_5_or_nl;
  wire nor_187_nl;
  wire return_add_generic_AC_RND_CONV_false_17_mux_19_nl;
  wire return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_and_3_nl;
  wire nor_191_nl;
  wire return_add_generic_AC_RND_CONV_false_18_mux_13_nl;
  wire return_add_generic_AC_RND_CONV_false_18_return_add_generic_AC_RND_CONV_false_18_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_5_nl;
  wire and_612_nl;
  wire return_add_generic_AC_RND_CONV_false_19_if_7_return_add_generic_AC_RND_CONV_false_19_if_7_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_19_e_r_qelse_mux_2_nl;
  wire or_438_nl;
  wire return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_6_nl;
  wire return_add_generic_AC_RND_CONV_false_19_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_19_if_5_or_nl;
  wire and_614_nl;
  wire return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_4_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_6_nl;
  wire or_443_nl;
  wire return_add_generic_AC_RND_CONV_false_20_r_nan_or_1_nl;
  wire and_615_nl;
  wire return_add_generic_AC_RND_CONV_false_20_if_7_return_add_generic_AC_RND_CONV_false_20_if_7_nor_nl;
  wire return_extract_57_return_extract_57_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_22_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_20_mux_18_nl;
  wire return_add_generic_AC_RND_CONV_false_20_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_1_nl;
  wire or_447_nl;
  wire and_616_nl;
  wire return_add_generic_AC_RND_CONV_false_21_if_7_return_add_generic_AC_RND_CONV_false_21_if_7_nor_nl;
  wire return_extract_59_return_extract_59_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_23_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_21_mux_14_nl;
  wire return_add_generic_AC_RND_CONV_false_21_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_22_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_22_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_23_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_23_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_24_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_24_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_25_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_25_if_5_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_if_if_not_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_mux_1_nl;
  wire[23:0] operator_32_false_2_acc_2_nl;
  wire[24:0] nl_operator_32_false_2_acc_2_nl;
  wire[12:0] return_mult_generic_AC_RND_CONV_false_1_if_acc_2_nl;
  wire[13:0] nl_return_mult_generic_AC_RND_CONV_false_1_if_acc_2_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_17_acc_3_nl;
  wire[11:0] nl_return_add_generic_AC_RND_CONV_false_17_acc_3_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_8_acc_3_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_8_acc_3_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_15_acc_3_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_15_acc_3_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_16_acc_3_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_16_acc_3_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_18_acc_3_nl;
  wire[11:0] nl_return_add_generic_AC_RND_CONV_false_18_acc_3_nl;
  wire mux_14_nl;
  wire mux_13_nl;
  wire mux_18_nl;
  wire mux_17_nl;
  wire mux_16_nl;
  wire mux_21_nl;
  wire mux_20_nl;
  wire mux_11_nl;
  wire mux_10_nl;
  wire or_76_nl;
  wire mux_9_nl;
  wire or_72_nl;
  wire[3:0] for_acc_nl;
  wire[4:0] nl_for_acc_nl;
  wire BUTTERFLY_1_i_mux1h_1_nl;
  wire[8:0] mux1h_6_nl;
  wire or_2033_nl;
  wire or_2009_nl;
  wire BUTTERFLY_if_1_if_mux1h_nl;
  wire BUTTERFLY_if_1_if_or_1_nl;
  wire[9:0] or_2027_nl;
  wire[9:0] and_2637_nl;
  wire[9:0] mux1h_1_nl;
  wire and_2629_nl;
  wire or_2745_nl;
  wire not_1022_nl;
  wire BUTTERFLY_if_1_if_mux1h_2_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_return_add_generic_AC_RND_CONV_false_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_2_nl;
  wire or_358_nl;
  wire return_add_generic_AC_RND_CONV_false_9_e_r_return_add_generic_AC_RND_CONV_false_9_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_nl;
  wire or_467_nl;
  wire return_add_generic_AC_RND_CONV_false_10_e_r_return_add_generic_AC_RND_CONV_false_10_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_7_nl;
  wire or_476_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_return_add_generic_AC_RND_CONV_false_11_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_2_nl;
  wire or_483_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_r_return_add_generic_AC_RND_CONV_false_12_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_3_nl;
  wire or_490_nl;
  wire BUTTERFLY_if_1_if_mux1h_3_nl;
  wire return_add_generic_AC_RND_CONV_false_9_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_10_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_11_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_12_r_nan_or_nl;
  wire BUTTERFLY_if_1_if_or_3_nl;
  wire BUTTERFLY_if_1_if_and_11_nl;
  wire[50:0] and_3934_nl;
  wire[50:0] mux1h_2_nl;
  wire nor_246_nl;
  wire BUTTERFLY_1_i_mux1h_nl;
  wire[8:0] BUTTERFLY_1_i_mux1h_6_nl;
  wire BUTTERFLY_else_1_if_or_nl;
  wire BUTTERFLY_if_1_mux1h_2_nl;
  wire[8:0] mux1h_7_nl;
  wire or_2034_nl;
  wire or_2010_nl;
  wire BUTTERFLY_if_1_mux1h_1_nl;
  wire BUTTERFLY_if_1_or_nl;
  wire BUTTERFLY_if_1_or_1_nl;
  wire[9:0] or_2028_nl;
  wire[9:0] and_2654_nl;
  wire[9:0] mux1h_3_nl;
  wire or_2746_nl;
  wire not_1025_nl;
  wire BUTTERFLY_if_1_mux1h_6_nl;
  wire return_add_generic_AC_RND_CONV_false_13_e_r_return_add_generic_AC_RND_CONV_false_13_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_5_nl;
  wire or_416_nl;
  wire return_add_generic_AC_RND_CONV_false_22_e_r_return_add_generic_AC_RND_CONV_false_22_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_8_nl;
  wire or_498_nl;
  wire return_add_generic_AC_RND_CONV_false_23_e_r_return_add_generic_AC_RND_CONV_false_23_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_4_nl;
  wire or_506_nl;
  wire return_add_generic_AC_RND_CONV_false_24_e_r_return_add_generic_AC_RND_CONV_false_24_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_9_nl;
  wire or_514_nl;
  wire return_add_generic_AC_RND_CONV_false_25_e_r_return_add_generic_AC_RND_CONV_false_25_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_3_nl;
  wire or_521_nl;
  wire BUTTERFLY_if_1_mux1h_7_nl;
  wire return_add_generic_AC_RND_CONV_false_22_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_23_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_24_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_25_r_nan_or_nl;
  wire[50:0] and_3935_nl;
  wire[50:0] mux1h_4_nl;
  wire nor_247_nl;
  wire BUTTERFLY_else_1_mux1h_nl;
  wire[8:0] BUTTERFLY_else_1_mux1h_1_nl;
  wire BUTTERFLY_else_1_if_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_7_exp_and_6_nl;
  wire return_add_generic_AC_RND_CONV_false_7_exp_and_7_nl;
  wire[51:0] and_2619_nl;
  wire nor_nl;
  wire or_1760_nl;
  wire or_1761_nl;
  wire return_mult_generic_AC_RND_CONV_false_return_mult_generic_AC_RND_CONV_false_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_return_mult_generic_AC_RND_CONV_false_1_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_return_mult_generic_AC_RND_CONV_false_2_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_return_mult_generic_AC_RND_CONV_false_3_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_return_mult_generic_AC_RND_CONV_false_4_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_return_mult_generic_AC_RND_CONV_false_5_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_4_nl;
  wire BUTTERFLY_1_else_1_if_and_4_nl;
  wire BUTTERFLY_1_else_1_if_and_5_nl;
  wire BUTTERFLY_1_else_1_if_and_6_nl;
  wire BUTTERFLY_1_else_1_if_and_7_nl;
  wire BUTTERFLY_1_else_1_if_and_8_nl;
  wire BUTTERFLY_1_else_1_if_and_9_nl;
  wire BUTTERFLY_1_else_1_if_and_10_nl;
  wire BUTTERFLY_1_else_1_if_and_11_nl;
  wire[8:0] BUTTERFLY_1_else_3_else_mux_2_nl;
  wire BUTTERFLY_1_else_3_else_mux_3_nl;
  wire[53:0] acc_nl;
  wire[54:0] nl_acc_nl;
  wire return_add_generic_AC_RND_CONV_false_22_ma1_lt_ma2_mux_4_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_22_ma1_lt_ma2_mux_5_nl;
  wire[53:0] acc_1_nl;
  wire[54:0] nl_acc_1_nl;
  wire return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_mux1h_4_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_mux1h_5_nl;
  wire[53:0] acc_4_nl;
  wire[54:0] nl_acc_4_nl;
  wire return_add_generic_AC_RND_CONV_false_6_ma1_lt_ma2_mux_5_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_6_ma1_lt_ma2_mux_6_nl;
  wire[15:0] BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_9_nl;
  wire[1:0] BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_10_nl;
  wire BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_or_1_nl;
  wire[1:0] BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_and_2_nl;
  wire[1:0] BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_11_nl;
  wire[10:0] BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_and_3_nl;
  wire BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_12_nl;
  wire[15:0] BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_13_nl;
  wire[17:0] acc_9_nl;
  wire[18:0] nl_acc_9_nl;
  wire[15:0] BUTTERFLY_else_1_if_mux_6_nl;
  wire[31:0] operator_32_false_acc_7_nl;
  wire[32:0] nl_operator_32_false_acc_7_nl;
  wire BUTTERFLY_else_mux_10_nl;
  wire stage_PE_stage_PE_stage_PE_mux_3_nl;
  wire BUTTERFLY_else_mux_11_nl;
  wire BUTTERFLY_else_mux_12_nl;
  wire BUTTERFLY_else_mux_13_nl;
  wire BUTTERFLY_else_mux_14_nl;
  wire BUTTERFLY_else_mux_15_nl;
  wire BUTTERFLY_else_mux_16_nl;
  wire BUTTERFLY_else_mux_17_nl;
  wire BUTTERFLY_else_mux_18_nl;
  wire BUTTERFLY_else_mux_19_nl;
  wire BUTTERFLY_fry_mux_10_nl;
  wire BUTTERFLY_fry_mux_11_nl;
  wire BUTTERFLY_fry_mux_12_nl;
  wire BUTTERFLY_fry_mux_13_nl;
  wire BUTTERFLY_fry_mux_14_nl;
  wire BUTTERFLY_fry_mux_15_nl;
  wire BUTTERFLY_fry_mux_16_nl;
  wire BUTTERFLY_fry_mux_17_nl;
  wire BUTTERFLY_fry_mux_18_nl;
  wire BUTTERFLY_fry_mux_19_nl;
  wire[13:0] acc_14_nl;
  wire[14:0] nl_acc_14_nl;
  wire[12:0] acc_10_nl;
  wire[13:0] nl_acc_10_nl;
  wire[9:0] return_mult_generic_AC_RND_CONV_false_2_exp_mux_7_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_exp_mux_8_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_exp_mux_9_nl;
  wire[12:0] acc_15_nl;
  wire[13:0] nl_acc_15_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_6_nl;
  wire[8:0] return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_7_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_8_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_9_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_10_nl;
  wire[12:0] acc_16_nl;
  wire[13:0] nl_acc_16_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_6_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_and_4_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_or_5_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_or_6_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_7_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_8_nl;
  wire[8:0] return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_9_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_10_nl;
  wire[12:0] acc_17_nl;
  wire[13:0] nl_acc_17_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_1_e_dif_mux_3_nl;
  wire[57:0] acc_19_nl;
  wire[58:0] nl_acc_19_nl;
  wire[55:0] return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_1_or_17_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_15_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux_35_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_16_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_1_mux1h_17_nl;
  wire return_add_generic_AC_RND_CONV_false_1_or_18_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_18_nl;
  wire[57:0] acc_20_nl;
  wire[58:0] nl_acc_20_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_12_mux1h_26_nl;
  wire[1:0] return_add_generic_AC_RND_CONV_false_12_mux1h_27_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_12_mux1h_28_nl;
  wire return_add_generic_AC_RND_CONV_false_12_mux1h_29_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_47_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_121_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_122_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_123_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_124_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_125_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_126_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_127_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_128_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_129_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_130_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_131_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_132_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_133_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_134_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_135_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_136_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_137_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_138_nl;
  wire return_add_generic_AC_RND_CONV_false_12_mux1h_30_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_48_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_49_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_50_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_51_nl;
  wire return_add_generic_AC_RND_CONV_false_12_mux1h_31_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_52_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_53_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_54_nl;
  wire return_add_generic_AC_RND_CONV_false_12_mux1h_32_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_12_mux1h_33_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_55_nl;
  wire return_add_generic_AC_RND_CONV_false_12_mux1h_34_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_56_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_57_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_58_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_59_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_60_nl;
  wire[10:0] operator_6_false_2_mux1h_3_nl;
  wire[5:0] operator_6_false_2_mux1h_4_nl;
  wire[5:0] operator_6_false_2_acc_1_nl;
  wire[6:0] nl_operator_6_false_2_acc_1_nl;
  wire[5:0] operator_6_false_acc_1_nl;
  wire[6:0] nl_operator_6_false_acc_1_nl;
  wire[5:0] operator_6_false_31_acc_1_nl;
  wire[6:0] nl_operator_6_false_31_acc_1_nl;
  wire[5:0] operator_6_false_29_acc_1_nl;
  wire[6:0] nl_operator_6_false_29_acc_1_nl;
  wire operator_6_false_33_mux1h_6_nl;
  wire[7:0] operator_6_false_33_mux1h_7_nl;
  wire operator_6_false_33_mux1h_8_nl;
  wire operator_6_false_33_mux1h_9_nl;
  wire operator_6_false_33_or_22_nl;
  wire[5:0] operator_6_false_33_mux1h_10_nl;
  wire[5:0] operator_6_false_23_acc_3_nl;
  wire[6:0] nl_operator_6_false_23_acc_3_nl;
  wire[5:0] operator_6_false_27_acc_3_nl;
  wire[6:0] nl_operator_6_false_27_acc_3_nl;
  wire operator_6_false_33_mux1h_11_nl;
  wire[13:0] acc_25_nl;
  wire[14:0] nl_acc_25_nl;
  wire[12:0] acc_22_nl;
  wire[13:0] nl_acc_22_nl;
  wire[9:0] return_mult_generic_AC_RND_CONV_false_exp_mux1h_6_nl;
  wire return_mult_generic_AC_RND_CONV_false_exp_mux1h_7_nl;
  wire return_mult_generic_AC_RND_CONV_false_exp_mux1h_8_nl;
  wire mux1h_29_nl;
  wire mux1h_23_nl;
  wire mux1h_34_nl;
  wire mux1h_27_nl;
  wire mux1h_31_nl;
  wire mux1h_24_nl;
  wire mux1h_22_nl;
  wire mux1h_33_nl;
  wire mux1h_26_nl;
  wire mux1h_36_nl;
  wire mux1h_35_nl;
  wire mux1h_56_nl;
  wire mux1h_57_nl;
  wire mux1h_38_nl;
  wire mux1h_58_nl;
  wire mux1h_55_nl;
  wire mux1h_45_nl;
  wire mux1h_54_nl;
  wire mux1h_60_nl;
  wire mux1h_59_nl;
  wire mux1h_32_nl;
  wire mux1h_28_nl;
  wire mux1h_51_nl;
  wire mux1h_46_nl;
  wire mux1h_8_nl;
  wire mux1h_9_nl;
  wire mux1h_10_nl;
  wire mux1h_11_nl;
  wire mux1h_30_nl;
  wire mux1h_20_nl;
  wire mux1h_19_nl;
  wire mux1h_18_nl;
  wire mux1h_17_nl;
  wire mux1h_16_nl;
  wire mux1h_15_nl;
  wire mux1h_14_nl;
  wire mux1h_13_nl;
  wire mux1h_12_nl;
  wire mux1h_49_nl;
  wire mux1h_44_nl;
  wire mux1h_41_nl;
  wire mux1h_52_nl;
  wire mux1h_53_nl;
  wire mux1h_47_nl;
  wire mux1h_42_nl;
  wire mux1h_39_nl;
  wire mux1h_43_nl;
  wire mux1h_50_nl;
  wire mux1h_48_nl;
  wire mux1h_40_nl;
  wire mux1h_37_nl;
  wire return_mult_generic_AC_RND_CONV_false_and_3_nl;
  wire mux1h_25_nl;
  wire return_mult_generic_AC_RND_CONV_false_mux_16_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_1_or_3_nl;
  wire return_add_generic_AC_RND_CONV_false_1_res_rounded_return_add_generic_AC_RND_CONV_false_1_res_rounded_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_1_res_rounded_mux_1_nl;
  wire[51:0] return_add_generic_AC_RND_CONV_false_1_res_rounded_mux1h_3_nl;
  wire return_add_generic_AC_RND_CONV_false_1_res_rounded_mux1h_4_nl;
  wire return_add_generic_AC_RND_CONV_false_1_res_rounded_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_mux_12_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_if_1_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_or_1_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_10_res_rounded_return_add_generic_AC_RND_CONV_false_10_res_rounded_mux_3_nl;
  wire return_add_generic_AC_RND_CONV_false_10_res_rounded_return_add_generic_AC_RND_CONV_false_10_res_rounded_mux_4_nl;
  wire return_add_generic_AC_RND_CONV_false_12_res_rounded_and_1_nl;
  wire[12:0] acc_29_nl;
  wire[13:0] nl_acc_29_nl;
  wire operator_6_false_3_mux1h_6_nl;
  wire[7:0] operator_6_false_3_mux1h_7_nl;
  wire operator_6_false_3_mux1h_8_nl;
  wire operator_6_false_3_mux1h_9_nl;
  wire operator_6_false_3_or_16_nl;
  wire operator_6_false_3_or_17_nl;
  wire[5:0] operator_6_false_3_mux1h_10_nl;
  wire operator_6_false_3_or_18_nl;
  wire operator_6_false_3_or_19_nl;
  wire[12:0] acc_30_nl;
  wire[13:0] nl_acc_30_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_dif1_return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_3_nl;
  wire[8:0] return_add_generic_AC_RND_CONV_false_6_e_dif1_return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_4_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_dif1_return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_5_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_6_e_dif1_mux1h_5_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_dif1_mux1h_6_nl;
  wire[12:0] acc_31_nl;
  wire[13:0] nl_acc_31_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_or_2_nl;
  wire[9:0] return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_mux1h_5_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_mux1h_6_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_or_1_nl;
  wire[9:0] return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_nor_1_nl;
  wire[9:0] return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_mux_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_or_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_mux_3_nl;
  wire[18:0] acc_33_nl;
  wire[19:0] nl_acc_33_nl;
  wire[4:0] stage_u_add_or_6_nl;
  wire[4:0] stage_u_add_stage_u_add_mux_2_nl;
  wire stage_u_add_or_7_nl;
  wire stage_u_add_stage_u_add_mux_3_nl;
  wire[9:0] stage_u_add_mux1h_7_nl;
  wire stage_u_add_mux1h_8_nl;
  wire stage_u_add_or_8_nl;
  wire[4:0] stage_u_add_and_1_nl;
  wire[4:0] stage_u_add_mux1h_9_nl;
  wire not_1086_nl;
  wire stage_u_add_mux1h_10_nl;
  wire[9:0] stage_u_add_mux1h_11_nl;
  wire BUTTERFLY_BUTTERFLY_or_2_nl;
  wire[3:0] BUTTERFLY_BUTTERFLY_or_3_nl;
  wire[3:0] BUTTERFLY_mux_1546_nl;
  wire[4:0] BUTTERFLY_mux1h_3_nl;
  wire[9:0] operator_6_false_10_mux_3_nl;
  wire[10:0] operator_33_true_7_mux1h_1_nl;
  wire operator_33_true_7_or_1_nl;
  wire BUTTERFLY_i_and_5_nl;
  wire BUTTERFLY_i_BUTTERFLY_i_mux_3_nl;
  wire BUTTERFLY_i_and_6_nl;
  wire BUTTERFLY_i_BUTTERFLY_i_mux_4_nl;
  wire[41:0] BUTTERFLY_i_BUTTERFLY_i_and_1_nl;
  wire[41:0] BUTTERFLY_i_mux_1_nl;
  wire not_1089_nl;
  wire[8:0] BUTTERFLY_i_mux1h_17_nl;
  wire BUTTERFLY_i_and_7_nl;
  wire BUTTERFLY_i_mux1h_18_nl;
  wire BUTTERFLY_i_and_8_nl;
  wire BUTTERFLY_i_mux1h_19_nl;
  wire[40:0] BUTTERFLY_i_and_9_nl;
  wire[40:0] BUTTERFLY_i_mux1h_20_nl;
  wire not_1092_nl;
  wire BUTTERFLY_i_mux1h_21_nl;
  wire BUTTERFLY_i_mux1h_22_nl;
  wire BUTTERFLY_i_mux1h_23_nl;
  wire BUTTERFLY_i_mux1h_24_nl;
  wire BUTTERFLY_i_mux1h_25_nl;
  wire BUTTERFLY_i_mux1h_26_nl;
  wire BUTTERFLY_i_mux1h_27_nl;
  wire BUTTERFLY_i_mux1h_28_nl;
  wire BUTTERFLY_i_mux1h_29_nl;
  wire BUTTERFLY_i_mux1h_30_nl;
  wire[13:0] BUTTERFLY_else_2_mux_4_nl;
  wire[1:0] BUTTERFLY_else_1_BUTTERFLY_else_1_and_1_nl;
  wire[4:0] BUTTERFLY_else_1_mux_9_nl;
  wire BUTTERFLY_else_1_mux_10_nl;
  wire[9:0] BUTTERFLY_else_1_mux_11_nl;
  wire[17:0] acc_39_nl;
  wire[18:0] nl_acc_39_nl;
  wire[4:0] operator_6_false_15_operator_6_false_15_or_2_nl;
  wire not_1093_nl;
  wire[5:0] operator_6_false_15_operator_6_false_15_or_3_nl;
  wire not_1094_nl;
  wire[5:0] operator_6_false_15_mux_4_nl;
  wire operator_6_false_15_or_1_nl;
  wire operator_6_false_15_mux_5_nl;
  wire[1:0] operator_6_false_15_operator_6_false_15_and_2_nl;
  wire not_1096_nl;
  wire[8:0] operator_6_false_15_operator_6_false_15_and_3_nl;
  wire not_1097_nl;
  wire operator_6_false_15_mux_6_nl;
  wire[9:0] operator_33_true_11_mux_1_nl;
  wire operator_32_false_2_operator_32_false_2_and_1_nl;
  wire[9:0] operator_32_false_2_mux_3_nl;
  wire return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_3_nl;
  wire [53:0] nl_return_mult_generic_AC_RND_CONV_false_6_else_1_rshift_rg_a;
  assign nl_return_mult_generic_AC_RND_CONV_false_6_else_1_rshift_rg_a = {1'b0 ,
      return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp
      , (out_f_d_rsci_q_d[51:1]) , 1'b0};
  wire [3:0] nl_return_mult_generic_AC_RND_CONV_false_6_else_1_rshift_rg_s;
  assign nl_return_mult_generic_AC_RND_CONV_false_6_else_1_rshift_rg_s = ~ (return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp[3:0]);
  wire[51:0] return_mult_generic_AC_RND_CONV_false_6_if_return_mult_generic_AC_RND_CONV_false_6_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_op1_normal_not_5_nl;
  wire [52:0] nl_leading_sign_53_0_6_rg_mantissa;
  assign return_mult_generic_AC_RND_CONV_false_6_op1_normal_not_5_nl = ~ return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp;
  assign return_mult_generic_AC_RND_CONV_false_6_if_return_mult_generic_AC_RND_CONV_false_6_if_and_nl
      = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000, (out_f_d_rsci_q_d[51:0]),
      return_mult_generic_AC_RND_CONV_false_6_op1_normal_not_5_nl);
  assign nl_leading_sign_53_0_6_rg_mantissa = {return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp
      , return_mult_generic_AC_RND_CONV_false_6_if_return_mult_generic_AC_RND_CONV_false_6_if_and_nl};
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_return_mult_generic_AC_RND_CONV_false_1_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_if_return_mult_generic_AC_RND_CONV_false_2_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_if_return_mult_generic_AC_RND_CONV_false_3_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_if_return_mult_generic_AC_RND_CONV_false_4_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_if_return_mult_generic_AC_RND_CONV_false_5_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_5_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_5_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_7_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_3_nl;
  wire[50:0] return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_9_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_if_and_1_nl;
  wire [52:0] nl_leading_sign_53_0_rg_mantissa;
  assign return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_nl
      = return_extract_15_return_extract_15_or_sva_1 & BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm;
  assign return_mult_generic_AC_RND_CONV_false_1_if_return_mult_generic_AC_RND_CONV_false_1_if_and_nl
      = return_extract_17_return_extract_17_or_sva_1 & BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm;
  assign return_mult_generic_AC_RND_CONV_false_2_if_return_mult_generic_AC_RND_CONV_false_2_if_and_nl
      = return_extract_19_return_extract_19_or_sva_1 & return_extract_41_return_extract_41_or_1_cse_sva;
  assign return_mult_generic_AC_RND_CONV_false_3_if_return_mult_generic_AC_RND_CONV_false_3_if_and_nl
      = return_extract_47_return_extract_47_or_sva_1 & BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm;
  assign return_mult_generic_AC_RND_CONV_false_4_if_return_mult_generic_AC_RND_CONV_false_4_if_and_nl
      = return_extract_49_return_extract_49_or_sva_1 & BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm;
  assign return_mult_generic_AC_RND_CONV_false_5_if_return_mult_generic_AC_RND_CONV_false_5_if_and_nl
      = return_extract_51_return_extract_51_or_sva_1 & return_extract_41_return_extract_41_or_1_cse_sva;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_nl
      = MUX1HOT_s_1_6_2(return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_nl,
      return_mult_generic_AC_RND_CONV_false_1_if_return_mult_generic_AC_RND_CONV_false_1_if_and_nl,
      return_mult_generic_AC_RND_CONV_false_2_if_return_mult_generic_AC_RND_CONV_false_2_if_and_nl,
      return_mult_generic_AC_RND_CONV_false_3_if_return_mult_generic_AC_RND_CONV_false_3_if_and_nl,
      return_mult_generic_AC_RND_CONV_false_4_if_return_mult_generic_AC_RND_CONV_false_4_if_and_nl,
      return_mult_generic_AC_RND_CONV_false_5_if_return_mult_generic_AC_RND_CONV_false_5_if_and_nl,
      {(fsm_output[11]) , (fsm_output[12]) , (fsm_output[13]) , (fsm_output[36])
      , (fsm_output[37]) , (fsm_output[38])});
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_5_nl =
      ((~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm) & or_dcpl_680) | ((~
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm) & or_dcpl_484);
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_5_nl
      = BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm & or_dcpl_680;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_7_nl
      = BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm & or_dcpl_484;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_2_nl =
      ((~ return_extract_41_return_extract_41_or_1_cse_sva) & (fsm_output[13])) |
      ((~ return_extract_41_return_extract_41_or_1_cse_sva) & (fsm_output[38]));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_1_nl
      = return_extract_41_return_extract_41_or_1_cse_sva & (fsm_output[13]);
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_3_nl
      = return_extract_41_return_extract_41_or_1_cse_sva & (fsm_output[38]);
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_1_nl
      = MUX1HOT_s_1_6_2(stage_PE_1_tmp_im_d_1_lpi_3_dfm_51, return_add_generic_AC_RND_CONV_false_4_m_r_51_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_1, (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[51]),
      return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0,
      {return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_5_nl , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_5_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_7_nl ,
      return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_2_nl , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_1_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_3_nl});
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_nor_nl
      = ~(BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm | return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse);
  assign return_mult_generic_AC_RND_CONV_false_1_if_and_nl = (~ or_dcpl_680) & BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm
      & (~ return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse);
  assign return_mult_generic_AC_RND_CONV_false_1_if_and_1_nl = or_dcpl_680 & BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm
      & (~ return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse);
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_9_nl
      = (~ return_extract_41_return_extract_41_or_1_cse_sva) & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse;
  assign return_mult_generic_AC_RND_CONV_false_2_if_and_nl = (~ (fsm_output[38]))
      & return_extract_41_return_extract_41_or_1_cse_sva & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse;
  assign return_mult_generic_AC_RND_CONV_false_2_if_and_1_nl = (fsm_output[38]) &
      return_extract_41_return_extract_41_or_1_cse_sva & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_nl
      = MUX1HOT_v_51_6_2(return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm,
      return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1,
      (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[50:0]), return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1, {return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_nor_nl
      , return_mult_generic_AC_RND_CONV_false_1_if_and_nl , return_mult_generic_AC_RND_CONV_false_1_if_and_1_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_9_nl ,
      return_mult_generic_AC_RND_CONV_false_2_if_and_nl , return_mult_generic_AC_RND_CONV_false_2_if_and_1_nl});
  assign nl_leading_sign_53_0_rg_mantissa = {return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_1_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_nl};
  wire [53:0] nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_a;
  assign nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_a = {(z_out_104[105:53])
      , 1'b0};
  wire return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_nl;
  wire[3:0] return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_2_nl;
  wire [5:0] nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_s;
  assign return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_nl
      = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_if_or_3_cse, return_mult_generic_AC_RND_CONV_false_2_if_or_3_cse,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse);
  assign return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_1_nl
      = MUX_v_4_2_2(return_mult_generic_AC_RND_CONV_false_if_nand_1_cse, return_mult_generic_AC_RND_CONV_false_2_if_nand_1_cse,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse);
  assign return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_2_nl
      = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_if_or_cse, return_mult_generic_AC_RND_CONV_false_2_if_or_cse,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse);
  assign nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_s = {return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_nl
      , return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_1_nl
      , return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_2_nl};
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_11_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_1_mux1h_13_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_12_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_13_rshift_rg_a;
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_nl = MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_op_smaller_qr_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_52_lpi_3_dfm_mx0,
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[11]) , (fsm_output[30]) ,
      (fsm_output[32])});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_11_nl = MUX1HOT_s_1_5_2((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      (return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_50_mx0,
      (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[11]) , (fsm_output[30]) ,
      (fsm_output[32])});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_13_nl = MUX1HOT_v_50_5_2((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      (return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0,
      (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[11]) , (fsm_output[30]) ,
      (fsm_output[32])});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_12_nl = MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_op_smaller_qr_0_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_0_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_0_lpi_3_dfm_mx0,
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[11]) , (fsm_output[30]) ,
      (fsm_output[32])});
  assign nl_return_add_generic_AC_RND_CONV_false_13_rshift_rg_a = {1'b0 , return_add_generic_AC_RND_CONV_false_1_mux1h_nl
      , return_add_generic_AC_RND_CONV_false_1_mux1h_11_nl , return_add_generic_AC_RND_CONV_false_1_mux1h_13_nl
      , return_add_generic_AC_RND_CONV_false_1_mux1h_12_nl , 3'b000};
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_13_rshift_rg_s;
  assign nl_return_add_generic_AC_RND_CONV_false_13_rshift_rg_s = MUX1HOT_v_6_5_2(return_add_generic_AC_RND_CONV_false_1_e_dif_sat_sva_1,
      return_add_generic_AC_RND_CONV_false_e_dif_sat_sva_1, return_add_generic_AC_RND_CONV_false_6_e_dif_sat_sva_1,
      return_add_generic_AC_RND_CONV_false_14_e_dif_sat_sva_1, return_add_generic_AC_RND_CONV_false_13_e_dif_sat_sva_1,
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[11]) , (fsm_output[30]) ,
      (fsm_output[32])});
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_6_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_3_mux1h_7_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_8_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_a;
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_nl = MUX1HOT_s_1_10_2(return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_op_smaller_qr_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx2,
      return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_52_lpi_3_dfm_mx0,
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm, {(fsm_output[5]) , (fsm_output[7])
      , (fsm_output[16]) , (fsm_output[18]) , (fsm_output[30]) , (fsm_output[32])
      , (fsm_output[36]) , (fsm_output[41]) , (fsm_output[43]) , BUTTERFLY_else_or_cse});
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_6_nl = MUX1HOT_s_1_10_2((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      (return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx2, return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_51_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_50_mx0,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx4, return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_51_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[50]),
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[16]) , (fsm_output[18]) ,
      (fsm_output[30]) , (fsm_output[32]) , (fsm_output[36]) , (fsm_output[41]) ,
      (fsm_output[43]) , BUTTERFLY_else_or_cse});
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_7_nl = MUX1HOT_v_50_10_2((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      (return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0,
      return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[49:0]),
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[16]) , (fsm_output[18]) ,
      (fsm_output[30]) , (fsm_output[32]) , (fsm_output[36]) , (fsm_output[41]) ,
      (fsm_output[43]) , BUTTERFLY_else_or_cse});
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_8_nl = MUX1HOT_s_1_10_2(return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_op_smaller_qr_0_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2,
      return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_0_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_0_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx3, return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm, {(fsm_output[5])
      , (fsm_output[7]) , (fsm_output[16]) , (fsm_output[18]) , (fsm_output[30])
      , (fsm_output[32]) , (fsm_output[36]) , (fsm_output[41]) , (fsm_output[43])
      , BUTTERFLY_else_or_cse});
  assign nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_a = {1'b0 , return_add_generic_AC_RND_CONV_false_3_mux1h_nl
      , return_add_generic_AC_RND_CONV_false_3_mux1h_6_nl , return_add_generic_AC_RND_CONV_false_3_mux1h_7_nl
      , return_add_generic_AC_RND_CONV_false_3_mux1h_8_nl , 3'b000};
  wire return_add_generic_AC_RND_CONV_false_3_or_3_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_s;
  assign return_add_generic_AC_RND_CONV_false_3_or_3_nl = (fsm_output[16]) | (fsm_output[36]);
  assign nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_s = MUX1HOT_v_6_9_2(return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse,
      return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1, return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_cse,
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_1, return_add_generic_AC_RND_CONV_false_16_e_dif_sat_sva_1,
      return_add_generic_AC_RND_CONV_false_15_e_dif_sat_sva_1, return_add_generic_AC_RND_CONV_false_22_e_dif_sat_sva_1,
      return_add_generic_AC_RND_CONV_false_23_e_dif_sat_sva_1, operator_6_false_17_acc_itm_6_1,
      {(fsm_output[5]) , (fsm_output[7]) , return_add_generic_AC_RND_CONV_false_3_or_3_nl
      , (fsm_output[18]) , (fsm_output[30]) , (fsm_output[32]) , (fsm_output[41])
      , (fsm_output[43]) , BUTTERFLY_else_or_cse});
  wire return_add_generic_AC_RND_CONV_false_7_mux_35_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_36_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_7_mux_37_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_38_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_20_rshift_rg_a;
  assign return_add_generic_AC_RND_CONV_false_7_mux_35_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_52_lpi_3_dfm_mx0, fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_7_mux_36_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_51_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_51_lpi_3_dfm_mx0, fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_7_mux_37_nl = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0, fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_7_mux_38_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_0_lpi_3_dfm_mx0, fsm_output[39]);
  assign nl_return_add_generic_AC_RND_CONV_false_20_rshift_rg_a = {1'b0 , return_add_generic_AC_RND_CONV_false_7_mux_35_nl
      , return_add_generic_AC_RND_CONV_false_7_mux_36_nl , return_add_generic_AC_RND_CONV_false_7_mux_37_nl
      , return_add_generic_AC_RND_CONV_false_7_mux_38_nl , 3'b000};
  wire return_add_generic_AC_RND_CONV_false_8_mux1h_nl;
  wire return_add_generic_AC_RND_CONV_false_8_mux1h_2_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_8_mux1h_3_nl;
  wire return_add_generic_AC_RND_CONV_false_8_mux1h_4_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_11_rshift_rg_a;
  assign return_add_generic_AC_RND_CONV_false_8_mux1h_nl = MUX1HOT_s_1_7_2(return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx2, return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx3,
      return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm,
      {(fsm_output[14]) , (fsm_output[16]) , (fsm_output[18]) , (fsm_output[39])
      , (fsm_output[41]) , (fsm_output[43]) , BUTTERFLY_else_or_cse});
  assign return_add_generic_AC_RND_CONV_false_8_mux1h_2_nl = MUX1HOT_s_1_7_2(return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_51_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx2, return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_51_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx4,
      return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_51_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[50]),
      {(fsm_output[14]) , (fsm_output[16]) , (fsm_output[18]) , (fsm_output[39])
      , (fsm_output[41]) , (fsm_output[43]) , BUTTERFLY_else_or_cse});
  assign return_add_generic_AC_RND_CONV_false_8_mux1h_3_nl = MUX1HOT_v_50_7_2(return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[49:0]),
      {(fsm_output[14]) , (fsm_output[16]) , (fsm_output[18]) , (fsm_output[39])
      , (fsm_output[41]) , (fsm_output[43]) , BUTTERFLY_else_or_cse});
  assign return_add_generic_AC_RND_CONV_false_8_mux1h_4_nl = MUX1HOT_s_1_7_2(return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2, return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_0_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx3,
      return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_0_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm,
      {(fsm_output[14]) , (fsm_output[16]) , (fsm_output[18]) , (fsm_output[39])
      , (fsm_output[41]) , (fsm_output[43]) , BUTTERFLY_else_or_cse});
  assign nl_return_add_generic_AC_RND_CONV_false_11_rshift_rg_a = {1'b0 , return_add_generic_AC_RND_CONV_false_8_mux1h_nl
      , return_add_generic_AC_RND_CONV_false_8_mux1h_2_nl , return_add_generic_AC_RND_CONV_false_8_mux1h_3_nl
      , return_add_generic_AC_RND_CONV_false_8_mux1h_4_nl , 3'b000};
  wire[4:0] return_add_generic_AC_RND_CONV_false_8_mux1h_1_nl;
  wire return_add_generic_AC_RND_CONV_false_8_mux1h_5_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_11_rshift_rg_s;
  assign return_add_generic_AC_RND_CONV_false_8_mux1h_1_nl = MUX1HOT_v_5_7_2((return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1[5:1]),
      (return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1[5:1]), (return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1[5:1]),
      (return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1[5:1]), (return_add_generic_AC_RND_CONV_false_24_e_dif_sat_sva_1[5:1]),
      (return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse[5:1]), return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_5_1,
      {(fsm_output[14]) , (fsm_output[16]) , (fsm_output[18]) , (fsm_output[39])
      , (fsm_output[41]) , (fsm_output[43]) , BUTTERFLY_else_or_cse});
  assign return_add_generic_AC_RND_CONV_false_8_mux1h_5_nl = MUX1HOT_s_1_7_2((return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1[0]),
      (return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1[0]), (return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1[0]),
      (return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1[0]), (return_add_generic_AC_RND_CONV_false_24_e_dif_sat_sva_1[0]),
      (return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse[0]), return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_0,
      {(fsm_output[14]) , (fsm_output[16]) , (fsm_output[18]) , (fsm_output[39])
      , (fsm_output[41]) , (fsm_output[43]) , BUTTERFLY_else_or_cse});
  assign nl_return_add_generic_AC_RND_CONV_false_11_rshift_rg_s = {return_add_generic_AC_RND_CONV_false_8_mux1h_1_nl
      , return_add_generic_AC_RND_CONV_false_8_mux1h_5_nl};
  wire return_add_generic_AC_RND_CONV_false_1_and_nl;
  wire return_add_generic_AC_RND_CONV_false_1_or_3_nl;
  wire return_add_generic_AC_RND_CONV_false_1_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_1_and_4_nl;
  wire return_add_generic_AC_RND_CONV_false_1_and_6_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_13_lshift_1_rg_s;
  assign return_add_generic_AC_RND_CONV_false_1_and_nl = (~ return_add_generic_AC_RND_CONV_false_1_acc_2_itm_11_1)
      & (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_1_or_3_nl = (return_add_generic_AC_RND_CONV_false_1_acc_2_itm_11_1
      & (fsm_output[5])) | (return_add_generic_AC_RND_CONV_false_acc_2_itm_11_1 &
      (fsm_output[7])) | (return_add_generic_AC_RND_CONV_false_14_acc_2_itm_11_1
      & (fsm_output[30])) | (return_add_generic_AC_RND_CONV_false_13_acc_2_itm_11_1
      & (fsm_output[32]));
  assign return_add_generic_AC_RND_CONV_false_1_and_2_nl = (~ return_add_generic_AC_RND_CONV_false_acc_2_itm_11_1)
      & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_1_and_4_nl = (~ return_add_generic_AC_RND_CONV_false_14_acc_2_itm_11_1)
      & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_1_and_6_nl = (~ return_add_generic_AC_RND_CONV_false_13_acc_2_itm_11_1)
      & (fsm_output[32]);
  assign nl_return_add_generic_AC_RND_CONV_false_13_lshift_1_rg_s = MUX1HOT_v_6_5_2((drf_qr_lval_1_smx_lpi_3_dfm_mx0[5:0]),
      rtn_out_1, (drf_qr_lval_10_smx_lpi_3_dfm_mx2[5:0]), (return_extract_32_mux_cse[5:0]),
      (drf_qr_lval_10_smx_lpi_3_dfm_mx6[5:0]), {return_add_generic_AC_RND_CONV_false_1_and_nl
      , return_add_generic_AC_RND_CONV_false_1_or_3_nl , return_add_generic_AC_RND_CONV_false_1_and_2_nl
      , return_add_generic_AC_RND_CONV_false_1_and_4_nl , return_add_generic_AC_RND_CONV_false_1_and_6_nl});
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_12_lshift_1_rg_a;
  assign nl_return_add_generic_AC_RND_CONV_false_12_lshift_1_rg_a = {return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_56
      , return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_0 , return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1};
  wire[3:0] return_add_generic_AC_RND_CONV_false_12_return_add_generic_AC_RND_CONV_false_12_mux1h_nl;
  wire return_add_generic_AC_RND_CONV_false_12_return_add_generic_AC_RND_CONV_false_12_mux1h_1_nl;
  wire return_add_generic_AC_RND_CONV_false_12_mux_22_nl;
  wire return_add_generic_AC_RND_CONV_false_12_exp_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_12_exp_mux_1_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_12_lshift_1_rg_s;
  assign return_add_generic_AC_RND_CONV_false_12_return_add_generic_AC_RND_CONV_false_12_mux1h_nl
      = MUX1HOT_v_4_3_2((drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0[3:0]), (operator_6_false_17_acc_itm_6_1[5:2]),
      (drf_qr_lval_21_smx_9_0_lpi_3_dfm[4:1]), {return_add_generic_AC_RND_CONV_false_12_return_add_generic_AC_RND_CONV_false_12_nor_1_ssc
      , return_add_generic_AC_RND_CONV_false_12_or_16_ssc , return_add_generic_AC_RND_CONV_false_12_and_6_ssc});
  assign return_add_generic_AC_RND_CONV_false_12_return_add_generic_AC_RND_CONV_false_12_mux1h_1_nl
      = MUX1HOT_s_1_3_2(drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1, (operator_6_false_17_acc_itm_6_1[1]),
      (drf_qr_lval_21_smx_9_0_lpi_3_dfm[0]), {return_add_generic_AC_RND_CONV_false_12_return_add_generic_AC_RND_CONV_false_12_nor_1_ssc
      , return_add_generic_AC_RND_CONV_false_12_or_16_ssc , return_add_generic_AC_RND_CONV_false_12_and_6_ssc});
  assign return_add_generic_AC_RND_CONV_false_12_exp_mux_nl = MUX_s_1_2_2(drf_qr_lval_15_smx_0_lpi_3_dfm,
      (operator_6_false_17_acc_itm_6_1[0]), return_add_generic_AC_RND_CONV_false_12_acc_2_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_12_exp_mux_1_nl = MUX_s_1_2_2(drf_qr_lval_15_smx_0_lpi_3_dfm,
      (operator_6_false_17_acc_itm_6_1[0]), return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_12_mux_22_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_12_exp_mux_nl,
      return_add_generic_AC_RND_CONV_false_12_exp_mux_1_nl, fsm_output[50]);
  assign nl_return_add_generic_AC_RND_CONV_false_12_lshift_1_rg_s = {return_add_generic_AC_RND_CONV_false_12_return_add_generic_AC_RND_CONV_false_12_mux1h_nl
      , return_add_generic_AC_RND_CONV_false_12_return_add_generic_AC_RND_CONV_false_12_mux1h_1_nl
      , return_add_generic_AC_RND_CONV_false_12_mux_22_nl};
  wire return_add_generic_AC_RND_CONV_false_2_or_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_a;
  assign return_add_generic_AC_RND_CONV_false_2_or_nl = operator_6_false_17_or_cse
      | or_dcpl_484 | (fsm_output[19]) | (fsm_output[23]) | (fsm_output[42]) | (fsm_output[46]);
  assign nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_a = MUX_v_57_2_2(return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva,
      return_add_generic_AC_RND_CONV_false_11_res_mant_4_sva, return_add_generic_AC_RND_CONV_false_2_or_nl);
  wire[3:0] return_add_generic_AC_RND_CONV_false_2_mux1h_nl;
  wire return_add_generic_AC_RND_CONV_false_2_mux1h_2_nl;
  wire return_add_generic_AC_RND_CONV_false_2_mux1h_1_nl;
  wire return_add_generic_AC_RND_CONV_false_2_or_13_nl;
  wire return_add_generic_AC_RND_CONV_false_2_or_14_nl;
  wire return_add_generic_AC_RND_CONV_false_2_or_8_nl;
  wire return_add_generic_AC_RND_CONV_false_2_or_9_nl;
  wire return_add_generic_AC_RND_CONV_false_2_or_11_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_s;
  assign return_add_generic_AC_RND_CONV_false_2_mux1h_nl = MUX1HOT_v_4_14_2((return_add_generic_AC_RND_CONV_false_2_mux_4_itm[5:2]),
      (return_add_generic_AC_RND_CONV_false_3_mux_15_itm[5:2]), (return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_5_1[4:1]),
      (operator_6_false_17_acc_itm_6_1[5:2]), (return_add_generic_AC_RND_CONV_false_7_mux_24_mx0_5_1[4:1]),
      (return_add_generic_AC_RND_CONV_false_8_mux_20_mx0[5:2]), (operator_14_false_1_acc_psp_sva_9_0[4:1]),
      (return_add_generic_AC_RND_CONV_false_9_ls_sva[5:2]), (drf_qr_lval_21_smx_9_0_lpi_3_dfm[4:1]),
      (return_add_generic_AC_RND_CONV_false_10_ls_sva[5:2]), (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[4:1]),
      (return_add_generic_AC_RND_CONV_false_11_ls_sva[5:2]), (return_add_generic_AC_RND_CONV_false_15_mux_4_itm_5_1[4:1]),
      (drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0[3:0]), {(fsm_output[9]) , operator_6_false_17_or_cse
      , or_2455_cse , or_dcpl_484 , or_dcpl_493 , or_dcpl_485 , return_add_generic_AC_RND_CONV_false_2_or_4_ssc
      , return_add_generic_AC_RND_CONV_false_2_and_1_cse , return_add_generic_AC_RND_CONV_false_2_and_2_cse
      , return_add_generic_AC_RND_CONV_false_2_or_5_cse , return_add_generic_AC_RND_CONV_false_2_or_6_ssc
      , return_add_generic_AC_RND_CONV_false_2_or_7_cse , (fsm_output[34]) , return_add_generic_AC_RND_CONV_false_2_and_8_cse});
  assign return_add_generic_AC_RND_CONV_false_2_mux1h_2_nl = MUX1HOT_s_1_14_2((return_add_generic_AC_RND_CONV_false_2_mux_4_itm[1]),
      (return_add_generic_AC_RND_CONV_false_3_mux_15_itm[1]), (return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_5_1[0]),
      (operator_6_false_17_acc_itm_6_1[1]), (return_add_generic_AC_RND_CONV_false_7_mux_24_mx0_5_1[0]),
      (return_add_generic_AC_RND_CONV_false_8_mux_20_mx0[1]), (operator_14_false_1_acc_psp_sva_9_0[0]),
      (return_add_generic_AC_RND_CONV_false_9_ls_sva[1]), (drf_qr_lval_21_smx_9_0_lpi_3_dfm[0]),
      (return_add_generic_AC_RND_CONV_false_10_ls_sva[1]), (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[0]),
      (return_add_generic_AC_RND_CONV_false_11_ls_sva[1]), (return_add_generic_AC_RND_CONV_false_15_mux_4_itm_5_1[0]),
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1, {(fsm_output[9]) , operator_6_false_17_or_cse
      , or_2455_cse , or_dcpl_484 , or_dcpl_493 , or_dcpl_485 , return_add_generic_AC_RND_CONV_false_2_or_4_ssc
      , return_add_generic_AC_RND_CONV_false_2_and_1_cse , return_add_generic_AC_RND_CONV_false_2_and_2_cse
      , return_add_generic_AC_RND_CONV_false_2_or_5_cse , return_add_generic_AC_RND_CONV_false_2_or_6_ssc
      , return_add_generic_AC_RND_CONV_false_2_or_7_cse , (fsm_output[34]) , return_add_generic_AC_RND_CONV_false_2_and_8_cse});
  assign return_add_generic_AC_RND_CONV_false_2_or_13_nl = ((~ return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1)
      & or_dcpl_493) | ((~ return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1)
      & (fsm_output[34]));
  assign return_add_generic_AC_RND_CONV_false_2_or_14_nl = (return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1
      & or_dcpl_493) | return_add_generic_AC_RND_CONV_false_2_or_5_cse | (return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1
      & (fsm_output[34]));
  assign return_add_generic_AC_RND_CONV_false_2_or_8_nl = return_add_generic_AC_RND_CONV_false_2_and_cse
      | return_add_generic_AC_RND_CONV_false_2_and_6_cse;
  assign return_add_generic_AC_RND_CONV_false_2_or_9_nl = return_add_generic_AC_RND_CONV_false_2_and_2_cse
      | return_add_generic_AC_RND_CONV_false_2_and_8_cse;
  assign return_add_generic_AC_RND_CONV_false_2_or_11_nl = return_add_generic_AC_RND_CONV_false_2_and_4_cse
      | return_add_generic_AC_RND_CONV_false_2_and_10_cse;
  assign return_add_generic_AC_RND_CONV_false_2_mux1h_1_nl = MUX1HOT_s_1_12_2((return_add_generic_AC_RND_CONV_false_2_mux_4_itm[0]),
      (return_add_generic_AC_RND_CONV_false_3_mux_15_itm[0]), return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_0,
      (operator_6_false_17_acc_itm_6_1[0]), drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1,
      (return_add_generic_AC_RND_CONV_false_10_ls_sva[0]), (return_add_generic_AC_RND_CONV_false_8_mux_20_mx0[0]),
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm, (return_add_generic_AC_RND_CONV_false_9_ls_sva[0]),
      drf_qr_lval_13_smx_0_lpi_3_dfm, drf_qr_lval_14_smx_0_lpi_3_dfm, (return_add_generic_AC_RND_CONV_false_11_ls_sva[0]),
      {(fsm_output[9]) , operator_6_false_17_or_cse , or_2455_cse , or_dcpl_484 ,
      return_add_generic_AC_RND_CONV_false_2_or_13_nl , return_add_generic_AC_RND_CONV_false_2_or_14_nl
      , or_dcpl_485 , return_add_generic_AC_RND_CONV_false_2_or_8_nl , return_add_generic_AC_RND_CONV_false_2_and_1_cse
      , return_add_generic_AC_RND_CONV_false_2_or_9_nl , return_add_generic_AC_RND_CONV_false_2_or_11_nl
      , return_add_generic_AC_RND_CONV_false_2_or_7_cse});
  assign nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_s = {return_add_generic_AC_RND_CONV_false_2_mux1h_nl
      , return_add_generic_AC_RND_CONV_false_2_mux1h_2_nl , return_add_generic_AC_RND_CONV_false_2_mux1h_1_nl};
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_mux_2_nl;
  wire[51:0] return_mult_generic_AC_RND_CONV_false_1_if_1_mux_3_nl;
  wire[51:0] return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_not_3_nl;
  wire [105:0] nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_a;
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_and_nl
      = (return_mult_generic_AC_RND_CONV_false_1_p_1_sva[105]) & (~ (fsm_output[54]));
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_mux_2_nl = MUX_s_1_2_2((return_mult_generic_AC_RND_CONV_false_1_p_1_sva[104]),
      return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp,
      fsm_output[54]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_mux_3_nl = MUX_v_52_2_2((return_mult_generic_AC_RND_CONV_false_1_p_1_sva[103:52]),
      (out_f_d_rsci_q_d[51:0]), fsm_output[54]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_not_3_nl = ~ (fsm_output[54]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_nl
      = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000, (return_mult_generic_AC_RND_CONV_false_1_p_1_sva[51:0]),
      return_mult_generic_AC_RND_CONV_false_1_if_1_not_3_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_a = {return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_and_nl
      , return_mult_generic_AC_RND_CONV_false_1_if_1_mux_2_nl , return_mult_generic_AC_RND_CONV_false_1_if_1_mux_3_nl
      , return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_nl};
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_and_4_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_and_5_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_and_6_nl;
  wire [5:0] nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_s;
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_nor_nl
      = ~((z_out_111[12]) | (fsm_output[54]));
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_and_4_nl = (z_out_111[12])
      & (~ (fsm_output[54]));
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_and_5_nl = (~ (operator_6_false_58_acc_psp_sva_1[11]))
      & (fsm_output[54]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_and_6_nl = (operator_6_false_58_acc_psp_sva_1[11])
      & (fsm_output[54]);
  assign nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_s = MUX1HOT_v_6_4_2(return_add_generic_AC_RND_CONV_false_10_ls_sva,
      (operator_14_false_1_acc_psp_sva_9_0[5:0]), leading_sign_53_0_6_out_1, (return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp[5:0]),
      {return_mult_generic_AC_RND_CONV_false_1_if_1_return_mult_generic_AC_RND_CONV_false_1_if_1_nor_nl
      , return_mult_generic_AC_RND_CONV_false_1_if_1_and_4_nl , return_mult_generic_AC_RND_CONV_false_1_if_1_and_5_nl
      , return_mult_generic_AC_RND_CONV_false_1_if_1_and_6_nl});
  wire return_add_generic_AC_RND_CONV_false_3_or_nl;
  wire [54:0] nl_return_add_generic_AC_RND_CONV_false_12_lshift_rg_a;
  assign return_add_generic_AC_RND_CONV_false_3_or_nl = (fsm_output[11]) | (fsm_output[12])
      | (fsm_output[13]) | (fsm_output[36]) | (fsm_output[37]) | (fsm_output[38])
      | return_add_generic_AC_RND_CONV_false_3_or_2_seb;
  assign nl_return_add_generic_AC_RND_CONV_false_12_lshift_rg_a = signext_55_54({return_add_generic_AC_RND_CONV_false_3_or_2_seb
      , return_add_generic_AC_RND_CONV_false_3_or_nl , 52'b1111111111111111111111111111111111111111111111111111});
  wire return_add_generic_AC_RND_CONV_false_3_and_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_3_nl;
  wire return_add_generic_AC_RND_CONV_false_3_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_4_nl;
  wire[2:0] return_add_generic_AC_RND_CONV_false_3_mux1h_9_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux1h_5_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_12_lshift_rg_s;
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_3_nl = MUX1HOT_s_1_10_2((return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse[5]),
      (return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1[5]), return_mult_generic_AC_RND_CONV_false_if_or_3_cse,
      return_mult_generic_AC_RND_CONV_false_2_if_or_3_cse, (return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1[5]),
      (return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1[5]), (return_add_generic_AC_RND_CONV_false_16_e_dif_sat_sva_1[5]),
      (return_add_generic_AC_RND_CONV_false_15_e_dif_sat_sva_1[5]), (return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1[5]),
      (operator_6_false_17_acc_itm_6_1[5]), {return_add_generic_AC_RND_CONV_false_3_or_4_cse
      , (fsm_output[7]) , operator_14_false_1_or_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse
      , (fsm_output[14]) , (fsm_output[18]) , (fsm_output[30]) , (fsm_output[32])
      , (fsm_output[39]) , BUTTERFLY_else_or_cse});
  assign return_add_generic_AC_RND_CONV_false_3_and_nl = return_add_generic_AC_RND_CONV_false_3_mux1h_3_nl
      & (~ (fsm_output[54]));
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_4_nl = MUX1HOT_s_1_10_2((return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse[4]),
      (return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1[4]), (return_mult_generic_AC_RND_CONV_false_if_nand_1_cse[3]),
      (return_mult_generic_AC_RND_CONV_false_2_if_nand_1_cse[3]), (return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1[4]),
      (return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1[4]), (return_add_generic_AC_RND_CONV_false_16_e_dif_sat_sva_1[4]),
      (return_add_generic_AC_RND_CONV_false_15_e_dif_sat_sva_1[4]), (return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1[4]),
      (operator_6_false_17_acc_itm_6_1[4]), {return_add_generic_AC_RND_CONV_false_3_or_4_cse
      , (fsm_output[7]) , operator_14_false_1_or_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse
      , (fsm_output[14]) , (fsm_output[18]) , (fsm_output[30]) , (fsm_output[32])
      , (fsm_output[39]) , BUTTERFLY_else_or_cse});
  assign return_add_generic_AC_RND_CONV_false_3_and_1_nl = return_add_generic_AC_RND_CONV_false_3_mux1h_4_nl
      & (~ (fsm_output[54]));
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_9_nl = MUX1HOT_v_3_11_2((return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse[3:1]),
      (return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1[3:1]), (return_mult_generic_AC_RND_CONV_false_if_nand_1_cse[2:0]),
      (return_mult_generic_AC_RND_CONV_false_2_if_nand_1_cse[2:0]), (return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1[3:1]),
      (return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1[3:1]), (return_add_generic_AC_RND_CONV_false_16_e_dif_sat_sva_1[3:1]),
      (return_add_generic_AC_RND_CONV_false_15_e_dif_sat_sva_1[3:1]), (return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1[3:1]),
      (~ (return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp[3:1])), (operator_6_false_17_acc_itm_6_1[3:1]),
      {return_add_generic_AC_RND_CONV_false_3_or_4_cse , (fsm_output[7]) , operator_14_false_1_or_cse
      , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse , (fsm_output[14])
      , (fsm_output[18]) , (fsm_output[30]) , (fsm_output[32]) , (fsm_output[39])
      , (fsm_output[54]) , BUTTERFLY_else_or_cse});
  assign return_add_generic_AC_RND_CONV_false_3_mux1h_5_nl = MUX1HOT_s_1_11_2((return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse[0]),
      (return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1[0]), return_mult_generic_AC_RND_CONV_false_if_or_cse,
      return_mult_generic_AC_RND_CONV_false_2_if_or_cse, (return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1[0]),
      (return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1[0]), (return_add_generic_AC_RND_CONV_false_16_e_dif_sat_sva_1[0]),
      (return_add_generic_AC_RND_CONV_false_15_e_dif_sat_sva_1[0]), (return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1[0]),
      (~ (return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp[0])), (operator_6_false_17_acc_itm_6_1[0]),
      {return_add_generic_AC_RND_CONV_false_3_or_4_cse , (fsm_output[7]) , operator_14_false_1_or_cse
      , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse , (fsm_output[14])
      , (fsm_output[18]) , (fsm_output[30]) , (fsm_output[32]) , (fsm_output[39])
      , (fsm_output[54]) , BUTTERFLY_else_or_cse});
  assign nl_return_add_generic_AC_RND_CONV_false_12_lshift_rg_s = {return_add_generic_AC_RND_CONV_false_3_and_nl
      , return_add_generic_AC_RND_CONV_false_3_and_1_nl , return_add_generic_AC_RND_CONV_false_3_mux1h_9_nl
      , return_add_generic_AC_RND_CONV_false_3_mux1h_5_nl};
  wire[4:0] return_add_generic_AC_RND_CONV_false_1_mux1h_6_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux1h_14_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_13_lshift_rg_s;
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_6_nl = MUX1HOT_v_5_7_2((return_add_generic_AC_RND_CONV_false_1_e_dif_sat_sva_1[5:1]),
      (return_add_generic_AC_RND_CONV_false_e_dif_sat_sva_1[5:1]), (return_add_generic_AC_RND_CONV_false_6_e_dif_sat_sva_1[5:1]),
      (return_add_generic_AC_RND_CONV_false_14_e_dif_sat_sva_1[5:1]), (return_add_generic_AC_RND_CONV_false_13_e_dif_sat_sva_1[5:1]),
      (return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_cse[5:1]), return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_5_1,
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[11]) , (fsm_output[30]) ,
      (fsm_output[32]) , (fsm_output[36]) , or_2707_itm});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_14_nl = MUX1HOT_s_1_7_2((return_add_generic_AC_RND_CONV_false_1_e_dif_sat_sva_1[0]),
      (return_add_generic_AC_RND_CONV_false_e_dif_sat_sva_1[0]), (return_add_generic_AC_RND_CONV_false_6_e_dif_sat_sva_1[0]),
      (return_add_generic_AC_RND_CONV_false_14_e_dif_sat_sva_1[0]), (return_add_generic_AC_RND_CONV_false_13_e_dif_sat_sva_1[0]),
      (return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_cse[0]), return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_0,
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[11]) , (fsm_output[30]) ,
      (fsm_output[32]) , (fsm_output[36]) , or_2707_itm});
  assign nl_return_add_generic_AC_RND_CONV_false_13_lshift_rg_s = {return_add_generic_AC_RND_CONV_false_1_mux1h_6_nl
      , return_add_generic_AC_RND_CONV_false_1_mux1h_14_nl};
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_10_lshift_rg_s;
  assign nl_return_add_generic_AC_RND_CONV_false_10_lshift_rg_s = MUX1HOT_v_6_4_2(return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_cse,
      return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_1, return_add_generic_AC_RND_CONV_false_22_e_dif_sat_sva_1,
      return_add_generic_AC_RND_CONV_false_23_e_dif_sat_sva_1, {(fsm_output[16])
      , (fsm_output[18]) , (fsm_output[41]) , (fsm_output[43])});
  wire [79:0] nl_stage_run_out1_rsci_inst_out1_rsci_idat;
  assign nl_stage_run_out1_rsci_inst_out1_rsci_idat = {out1_rsci_idat_79_64 , out1_rsci_idat_63
      , out1_rsci_idat_62_52 , out1_rsci_idat_51 , out1_rsci_idat_50_0};
  wire nl_stage_run_run_fsm_inst_for_C_0_tr0;
  assign nl_stage_run_run_fsm_inst_for_C_0_tr0 = for_i_3_0_sva[0];
  wire nl_stage_run_run_fsm_inst_for_1_C_2_tr0;
  assign nl_stage_run_run_fsm_inst_for_1_C_2_tr0 = z_out_113[10];
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd16)) mode1_rsci (
      .dat(mode1_rsc_dat),
      .idat(mode1_rsci_idat)
    );
  leading_sign_57_0_1_0 leading_sign_57_0_1_0_19_rg (
      .mantissa(z_out_81),
      .all_same(leading_sign_57_0_1_0_19_out_2),
      .rtn(leading_sign_57_0_1_0_19_out_3)
    );
  mgc_shift_r_v5 #(.width_a(32'sd54),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd54)) return_mult_generic_AC_RND_CONV_false_6_else_1_rshift_rg (
      .a(nl_return_mult_generic_AC_RND_CONV_false_6_else_1_rshift_rg_a[53:0]),
      .s(nl_return_mult_generic_AC_RND_CONV_false_6_else_1_rshift_rg_s[3:0]),
      .z(return_mult_generic_AC_RND_CONV_false_6_else_1_rshift_itm)
    );
  leading_sign_53_0 leading_sign_53_0_6_rg (
      .mantissa(nl_leading_sign_53_0_6_rg_mantissa[52:0]),
      .rtn(leading_sign_53_0_6_out_1)
    );
  leading_sign_53_0 leading_sign_53_0_rg (
      .mantissa(nl_leading_sign_53_0_rg_mantissa[52:0]),
      .rtn(rtn_out)
    );
  mgc_shift_r_v5 #(.width_a(32'sd54),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd54)) return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg (
      .a(nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_a[53:0]),
      .s(nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_s[5:0]),
      .z(z_out_65)
    );
  mgc_shift_r_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_13_rshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_13_rshift_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_13_rshift_rg_s[5:0]),
      .z(z_out_73)
    );
  mgc_shift_r_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_10_rshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_s[5:0]),
      .z(z_out_74)
    );
  mgc_shift_r_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_20_rshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_20_rshift_rg_a[56:0]),
      .s(return_add_generic_AC_RND_CONV_false_7_mux_33_cse),
      .z(z_out_75)
    );
  mgc_shift_r_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_11_rshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_11_rshift_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_11_rshift_rg_s[5:0]),
      .z(z_out_76)
    );
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_13_lshift_1_rg (
      .a(z_out_80),
      .s(nl_return_add_generic_AC_RND_CONV_false_13_lshift_1_rg_s[5:0]),
      .z(z_out_77)
    );
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_12_lshift_1_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_12_lshift_1_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_12_lshift_1_rg_s[5:0]),
      .z(z_out_78)
    );
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_10_lshift_1_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_s[5:0]),
      .z(z_out_79)
    );
  leading_sign_57_0_1_0 leading_sign_57_0_1_0_rg (
      .mantissa(z_out_80),
      .all_same(all_same_out),
      .rtn(rtn_out_1)
    );
  leading_sign_57_0_1_0 leading_sign_57_0_1_0_10_rg (
      .mantissa(z_out_81),
      .all_same(all_same_out_1),
      .rtn(rtn_out_2)
    );
  mgc_shift_l_v5 #(.width_a(32'sd106),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd106)) return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg (
      .a(nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_a[105:0]),
      .s(nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_s[5:0]),
      .z(z_out_106)
    );
  mgc_shift_l_v5 #(.width_a(32'sd55),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd55)) return_add_generic_AC_RND_CONV_false_12_lshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_12_lshift_rg_a[54:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_12_lshift_rg_s[5:0]),
      .z(z_out_107)
    );
  mgc_shift_l_v5 #(.width_a(32'sd55),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd55)) return_add_generic_AC_RND_CONV_false_20_lshift_rg (
      .a(55'b1111111111111111111111111111111111111111111111111111111),
      .s(return_add_generic_AC_RND_CONV_false_7_mux_33_cse),
      .z(z_out_108)
    );
  mgc_shift_l_v5 #(.width_a(32'sd55),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd55)) return_add_generic_AC_RND_CONV_false_13_lshift_rg (
      .a(55'b1111111111111111111111111111111111111111111111111111111),
      .s(nl_return_add_generic_AC_RND_CONV_false_13_lshift_rg_s[5:0]),
      .z(z_out_109)
    );
  mgc_shift_l_v5 #(.width_a(32'sd55),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd55)) return_add_generic_AC_RND_CONV_false_10_lshift_rg (
      .a(55'b1111111111111111111111111111111111111111111111111111111),
      .s(nl_return_add_generic_AC_RND_CONV_false_10_lshift_rg_s[5:0]),
      .z(z_out_110)
    );
  stage_run_ap_start_rsci stage_run_ap_start_rsci_inst (
      .ap_start_rsc_dat(ap_start_rsc_dat),
      .ap_start_rsc_vld(ap_start_rsc_vld),
      .ap_start_rsc_rdy(ap_start_rsc_rdy),
      .ap_start_rsci_oswt(reg_ap_start_rsci_iswt0_cse),
      .ap_start_rsci_wen_comp(ap_start_rsci_wen_comp)
    );
  stage_run_ap_done_rsci stage_run_ap_done_rsci_inst (
      .ap_done_rsc_dat(ap_done_rsc_dat),
      .ap_done_rsc_vld(ap_done_rsc_vld),
      .ap_done_rsc_rdy(ap_done_rsc_rdy),
      .ap_done_rsci_oswt(reg_out_u_triosy_obj_iswt0_cse),
      .ap_done_rsci_wen_comp(ap_done_rsci_wen_comp)
    );
  stage_run_wait_dp stage_run_wait_dp_inst (
      .in_f_d_rsci_en_d(in_f_d_rsci_en_d),
      .in_u_rsci_en_d(in_u_rsci_en_d),
      .out_f_d_rsci_en_d(out_f_d_rsci_en_d),
      .out_u_rsci_en_d(out_u_rsci_en_d),
      .BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en),
      .BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en(BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en),
      .BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en),
      .BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en(BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en),
      .r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en),
      .run_wen(run_wen),
      .in_f_d_rsci_cgo(reg_in_f_d_rsci_cgo_ir_cse),
      .in_f_d_rsci_cgo_ir_unreg(or_1122_rmff),
      .in_u_rsci_cgo(reg_in_u_rsci_cgo_ir_cse),
      .in_u_rsci_cgo_ir_unreg(or_1121_rmff),
      .out_f_d_rsci_cgo(reg_out_f_d_rsci_cgo_ir_cse),
      .out_f_d_rsci_cgo_ir_unreg(or_1120_rmff),
      .out_u_rsci_cgo(reg_out_u_rsci_cgo_ir_cse),
      .out_u_rsci_cgo_ir_unreg(or_1119_rmff),
      .BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo),
      .BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo(BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo),
      .BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo),
      .BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo(BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo),
      .r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_cgo(reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_cgo_cse)
    );
  stage_run_out1_rsci stage_run_out1_rsci_inst (
      .out1_rsc_dat(out1_rsc_dat),
      .out1_rsc_vld(out1_rsc_vld),
      .out1_rsc_rdy(out1_rsc_rdy),
      .out1_rsci_oswt(reg_out1_rsci_iswt0_cse),
      .out1_rsci_wen_comp(out1_rsci_wen_comp),
      .out1_rsci_idat(nl_stage_run_out1_rsci_inst_out1_rsci_idat[79:0])
    );
  stage_run_mode1_triosy_obj stage_run_mode1_triosy_obj_inst (
      .mode1_triosy_lz(mode1_triosy_lz),
      .run_wten(run_wten),
      .mode1_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_in_f_d_triosy_obj stage_run_in_f_d_triosy_obj_inst (
      .in_f_d_triosy_lz(in_f_d_triosy_lz),
      .run_wten(run_wten),
      .in_f_d_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_in_u_triosy_obj stage_run_in_u_triosy_obj_inst (
      .in_u_triosy_lz(in_u_triosy_lz),
      .run_wten(run_wten),
      .in_u_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_out_f_d_triosy_obj stage_run_out_f_d_triosy_obj_inst (
      .out_f_d_triosy_lz(out_f_d_triosy_lz),
      .run_wten(run_wten),
      .out_f_d_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_out_u_triosy_obj stage_run_out_u_triosy_obj_inst (
      .out_u_triosy_lz(out_u_triosy_lz),
      .run_wten(run_wten),
      .out_u_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_staller stage_run_staller_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .ap_start_rsci_wen_comp(ap_start_rsci_wen_comp),
      .ap_done_rsci_wen_comp(ap_done_rsci_wen_comp),
      .out1_rsci_wen_comp(out1_rsci_wen_comp)
    );
  stage_run_run_fsm stage_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .for_C_0_tr0(nl_stage_run_run_fsm_inst_for_C_0_tr0),
      .BUTTERFLY_C_24_tr0(and_dcpl_159),
      .BUTTERFLY_C_24_tr1(and_dcpl_160),
      .BUTTERFLY_1_C_24_tr0(and_dcpl_159),
      .BUTTERFLY_1_C_24_tr1(and_dcpl_160),
      .for_1_C_2_tr0(nl_stage_run_run_fsm_inst_for_1_C_2_tr0)
    );
  assign for_1_if_and_ssc = run_wen & (or_tmp_64 | out1_rsci_idat_63_0_mx0c1 | out1_rsci_idat_63_0_mx0c2);
  assign or_1119_rmff = and_647_cse | (~(mode_lpi_1_dfm | (~(or_dcpl_204 | (fsm_output[33])
      | (fsm_output[6]) | (fsm_output[5]) | (fsm_output[32]))))) | (operator_16_false_operator_16_false_nor_cse_sva
      & or_dcpl_207) | (and_dcpl_185 & (fsm_output[34]));
  assign or_1120_rmff = (and_dcpl_18 & ((fsm_output[50]) | (fsm_output[51]) | (fsm_output[45])
      | (fsm_output[52]) | (fsm_output[47]) | (fsm_output[49]) | or_dcpl_209 | (fsm_output[9])
      | or_dcpl_208)) | (mode_lpi_1_dfm & (or_dcpl_204 | (fsm_output[7:6]!=2'b00)))
      | (stage_PE_1_and_1_tmp & (or_dcpl_224 | or_dcpl_223 | or_dcpl_221 | (fsm_output[33])
      | (fsm_output[5]))) | (or_dcpl_227 & or_dcpl_207);
  assign or_1121_rmff = (~(mode_lpi_1_dfm | (~(or_dcpl_230 | (fsm_output[7]) | or_dcpl_228
      | (fsm_output[31]))))) | (and_dcpl_183 & (fsm_output[55])) | and_660_cse |
      (and_dcpl_185 & (fsm_output[9])) | and_662_cse;
  assign or_1122_rmff = (mode_lpi_1_dfm & (or_dcpl_230 | or_dcpl_233)) | (and_dcpl_18
      & ((fsm_output[27]) | (fsm_output[26]) | (fsm_output[23]) | or_dcpl_240 | or_dcpl_236
      | (fsm_output[34]) | or_dcpl_235)) | (stage_PE_1_and_1_tmp & (or_dcpl_248 |
      (fsm_output[17:16]!=2'b00) | or_dcpl_245 | or_dcpl_228)) | and_660_cse;
  assign r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_addr = reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_addr_cse;
  assign BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr = reg_BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_addr_cse;
  assign or_1132_ssc = (fsm_output[5]) | (fsm_output[31]) | return_add_generic_AC_RND_CONV_false_12_and_112_cse;
  assign or_1133_ssc = (fsm_output[33]) | and_680_cse;
  assign and_317_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_13_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign and_368_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_22_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign and_374_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_23_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign and_382_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_24_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign and_389_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_25_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign or_1146_ssc = (fsm_output[4]) | (fsm_output[10]);
  assign or_1147_ssc = (fsm_output[49]) | (fsm_output[41]) | (fsm_output[9]) | (fsm_output[5]);
  assign or_1148_ssc = (fsm_output[45]) | (fsm_output[33]) | (fsm_output[6]);
  assign or_1150_ssc = (fsm_output[51]) | (fsm_output[47]) | (fsm_output[43]);
  assign or_1159_ssc = return_add_generic_AC_RND_CONV_false_11_and_10_cse | (fsm_output[30])
      | (fsm_output[6]);
  assign or_1160_ssc = and_746_cse | (fsm_output[8]);
  assign and_281_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign and_340_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_9_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign and_348_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_10_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign and_356_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign and_362_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_12_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign BUTTERFLY_if_1_if_or_cse = (fsm_output[8]) | (fsm_output[20]);
  assign return_add_generic_AC_RND_CONV_false_r_nan_or_cse = return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_mx2w0
      | return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0 | (return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0
      & return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0 & return_add_generic_AC_RND_CONV_false_20_do_sub_sva);
  assign and_2472_tmp = and_dcpl_231 & and_dcpl_503;
  assign or_1174_ssc = (fsm_output[20]) | (fsm_output[8]) | (fsm_output[31]);
  assign or_1176_ssc = (fsm_output[24]) | (fsm_output[16]) | (fsm_output[34]) | (fsm_output[30]);
  assign or_1177_ssc = or_dcpl_273 | (fsm_output[18]);
  assign or_1179_ssc = (fsm_output[29]) | (fsm_output[35]);
  assign nand_102_cse = ~(reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd
      & return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp);
  assign operator_16_false_and_cse = run_wen & (~ and_dcpl_323);
  assign t_in_and_cse = run_wen & ((fsm_output[1]) | (fsm_output[27]) | (fsm_output[52]));
  assign t_in_or_3_cse = (fsm_output[27]) | (fsm_output[52]);
  assign t_in_and_3_cse = t_in_and_cse & (~(and_dcpl_160 & t_in_or_3_cse));
  assign mode_and_cse = run_wen & (~(and_dcpl_323 & and_dcpl_327));
  assign or_2748_cse = and_225_cse | (z_out_101[9]);
  assign stage_PE_1_and_2_cse = run_wen & (~(and_dcpl_330 & and_dcpl_327));
  assign and_435_cse = return_add_generic_AC_RND_CONV_false_22_e1_eq_e2_equal_tmp
      & z_out_53_52;
  assign or_547_cse = and_435_cse | (z_out_96[11]);
  assign and_1046_cse = and_dcpl_340 & (fsm_output[41]);
  assign and_1057_cse = or_547_cse & (fsm_output[41]);
  assign or_1302_cse = and_1046_cse | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse;
  assign nor_174_m1c = ~(or_tmp | or_tmp_954 | or_tmp_955 | or_tmp_956);
  assign BUTTERFLY_else_or_cse = (fsm_output[6]) | (fsm_output[31]);
  assign return_add_generic_AC_RND_CONV_false_19_exp_plus_1_and_cse = run_wen & (~
      or_dcpl_484);
  assign BUTTERFLY_1_i_and_ssc = run_wen & ((inverse_lpi_1_dfm_1 & (~(and_dcpl_421
      & and_dcpl_323 & and_dcpl_389 & (~ (fsm_output[49])) & (~((fsm_output[55])
      | (fsm_output[46]) | (fsm_output[42]))) & (~((fsm_output[48]) | (fsm_output[23])
      | (fsm_output[22]))) & and_dcpl_382 & (~ (fsm_output[21])) & (~((fsm_output[17])
      | (fsm_output[54]) | (fsm_output[53])))))) | or_dcpl_198 | BUTTERFLY_1_i_9_0_sva_mx0c3);
  assign return_add_generic_AC_RND_CONV_false_10_and_cse = run_wen & ((inverse_lpi_1_dfm_1
      & (~((~((fsm_output[51]) | (fsm_output[45]))) & nor_34_cse & and_dcpl_420 &
      and_dcpl_330 & (~((fsm_output[55]) | (fsm_output[46]))) & and_dcpl_369 & and_dcpl_360
      & and_dcpl_382 & (~((fsm_output[43]) | (fsm_output[18]) | (fsm_output[54])))
      & and_dcpl_344 & (~ (fsm_output[31]))))) | (fsm_output[4]) | (fsm_output[20])
      | (fsm_output[29]) | (fsm_output[47]));
  assign or_1341_cse = (fsm_output[7]) | (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_13_or_cse = (fsm_output[7]) | (fsm_output[19])
      | (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_13_or_3_cse = (fsm_output[21]) | (fsm_output[23])
      | (fsm_output[25]) | (fsm_output[44]) | (fsm_output[46]) | (fsm_output[48])
      | (fsm_output[50]);
  assign return_add_generic_AC_RND_CONV_false_13_and_1_cse = (~ return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp)
      & (fsm_output[12]);
  assign return_add_generic_AC_RND_CONV_false_13_and_3_cse = (~ return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp)
      & (fsm_output[37]);
  assign return_add_generic_AC_RND_CONV_false_13_and_2_cse = return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp
      & (fsm_output[12]);
  assign return_add_generic_AC_RND_CONV_false_13_and_4_cse = return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp
      & (fsm_output[37]);
  assign return_add_generic_AC_RND_CONV_false_13_or_4_cse = return_add_generic_AC_RND_CONV_false_13_and_1_cse
      | return_add_generic_AC_RND_CONV_false_13_and_3_cse;
  assign return_add_generic_AC_RND_CONV_false_10_exp_mux1h_3_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1,
      (stage_PE_1_tmp_re_d_sva[52]), and_dcpl_446);
  assign return_add_generic_AC_RND_CONV_false_10_exp_mux1h_6_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1,
      (stage_PE_1_tmp_re_d_sva[52]), and_dcpl_447);
  assign return_add_generic_AC_RND_CONV_false_13_or_2_cse = (fsm_output[4]) | (fsm_output[6]);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse = (fsm_output[5])
      | (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_or_5_cse = (fsm_output[31:30]!=2'b00);
  assign and_517_tmp = (~ return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp)
      & inverse_lpi_1_dfm_1;
  assign return_extract_33_or_1_tmp = return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx8c1
      | ((~ return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp)
      & return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx8c2);
  assign return_extract_2_mux_4_cse = MUX_v_51_2_2((out_f_d_rsci_q_d[50:0]), (out_f_d_rsci_q_d[51:1]),
      return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp);
  assign return_extract_33_mux_3_cse = MUX_v_51_2_2((in_f_d_rsci_q_d[50:0]), (in_f_d_rsci_q_d[51:1]),
      return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp);
  assign stage_PE_1_tmp_re_d_or_3_cse = (fsm_output[29]) | (fsm_output[31]);
  assign return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse = (fsm_output[5]) |
      (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_18_exp_and_3_cse = (~ and_dcpl_446)
      & (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_18_exp_and_5_cse = (~ and_dcpl_447)
      & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_18_exp_and_6_cse = and_dcpl_447 & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_18_exp_and_4_cse = and_dcpl_446 & (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_18_exp_or_cse = return_add_generic_AC_RND_CONV_false_18_exp_and_4_cse
      | return_add_generic_AC_RND_CONV_false_18_exp_and_6_cse;
  assign return_add_generic_AC_RND_CONV_false_18_exp_and_2_itm = and_dcpl_460 & return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_6_nl = MUX_s_1_2_2(and_dcpl_467,
      and_dcpl_469, fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_cse = run_wen & ((~(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_6_nl
      | or_dcpl_628)) | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[13]) | (fsm_output[16])
      | (fsm_output[30]) | (fsm_output[32]) | (fsm_output[38]) | (fsm_output[41]));
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse = (fsm_output[13])
      | (fsm_output[38]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse = and_dcpl_466
      & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_7_cse = ((~ and_dcpl_448)
      & (fsm_output[5])) | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_8_cse = (and_dcpl_448
      & (fsm_output[5])) | (and_dcpl_452 & (fsm_output[30]));
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_9_cse = ((~ and_dcpl_466)
      & (fsm_output[7])) | ((~ and_dcpl_468) & (fsm_output[32]));
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse = (~ and_dcpl_341)
      & (fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse = and_dcpl_468
      & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_10_cse = ((~ and_dcpl_452)
      & (fsm_output[30])) | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse = (~ and_dcpl_340)
      & (fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse = and_dcpl_341
      & (fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse = and_dcpl_469
      & (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_32_cse = and_dcpl_467
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_12_and_95_cse = (~ return_add_generic_AC_RND_CONV_false_12_do_sub_sva)
      & (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_12_and_103_cse = (~ return_add_generic_AC_RND_CONV_false_12_do_sub_sva)
      & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_12_and_96_cse = return_add_generic_AC_RND_CONV_false_12_do_sub_sva
      & (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_12_and_104_cse = return_add_generic_AC_RND_CONV_false_12_do_sub_sva
      & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_12_and_89_cse = (~ return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1)
      & (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_12_and_90_cse = return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1
      & (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_12_and_91_cse = (~ return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1)
      & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_12_and_92_cse = return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1
      & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_12_and_97_cse = (~ return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1)
      & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_12_and_98_cse = return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1
      & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_12_and_99_cse = (~ return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1)
      & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_12_and_100_cse = return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1
      & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_12_op_bigger_and_cse = run_wen & (~
      or_dcpl_635);
  assign return_add_generic_AC_RND_CONV_false_12_op_bigger_and_1_cse = run_wen &
      (~(or_dcpl_585 | or_dcpl_269 | or_dcpl_597));
  assign return_extract_41_and_1_cse = run_wen & (~(or_dcpl_645 | (fsm_output[10])
      | (fsm_output[36]) | (fsm_output[11]) | or_dcpl_553 | or_dcpl_632 | or_dcpl_640))
      & mode_lpi_1_dfm;
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_cse = run_wen & (~
      or_dcpl_628);
  assign BUTTERFLY_1_fiy_mux1h_4_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1,
      (stage_PE_1_x_re_d_sva[52]), and_dcpl_341);
  assign BUTTERFLY_1_fiy_mux1h_10_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1,
      (stage_PE_1_x_re_d_sva[52]), and_dcpl_340);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_4_cse = return_add_generic_AC_RND_CONV_false_10_do_sub_sva
      & BUTTERFLY_else_or_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_3_cse = (~ return_add_generic_AC_RND_CONV_false_10_do_sub_sva)
      & BUTTERFLY_else_or_cse;
  assign and_606_cse = return_add_generic_AC_RND_CONV_false_23_e1_eq_e2_equal_tmp
      & z_out_54_52;
  assign or_1102_cse = and_606_cse | (z_out_70[11]);
  assign or_1993_cse = or_1102_cse & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_7_exp_mux1h_4_itm_9_0 = MUX_v_10_2_2((return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[9:0]),
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1, and_dcpl_469);
  assign return_add_generic_AC_RND_CONV_false_17_and_2_m1c = or_dcpl_684 & return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse;
  assign return_add_generic_AC_RND_CONV_false_17_and_1_cse = (~ or_dcpl_684) & return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse;
  assign return_add_generic_AC_RND_CONV_false_17_and_3_cse = (~ or_658_cse) & return_add_generic_AC_RND_CONV_false_17_and_2_m1c;
  assign return_add_generic_AC_RND_CONV_false_17_and_4_cse = or_658_cse & return_add_generic_AC_RND_CONV_false_17_and_2_m1c;
  assign return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_and_1_cse
      = z_out_54_52 & return_add_generic_AC_RND_CONV_false_1_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_and_1_cse
      | (z_out_70[11]);
  assign return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_and_cse
      = z_out_54_52 & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_and_cse
      | (z_out_95[11]);
  assign return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse
      = (return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_itm_52 & return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp)
      | (z_out_70[11]);
  assign return_add_generic_AC_RND_CONV_false_12_and_106_m1c = or_dcpl_708 & (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_12_and_108_m1c = or_dcpl_709 & (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_12_and_114_m1c = or_dcpl_711 & (fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_12_and_105_cse = (~ or_dcpl_708) &
      (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_12_and_111_cse = return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse
      & and_dcpl_501 & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_12_and_107_cse = (~ or_dcpl_709) &
      (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_12_and_112_cse = (~ inverse_lpi_1_dfm_1)
      & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_12_and_109_cse = return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp
      & return_add_generic_AC_RND_CONV_false_15_aif_equal_tmp & inverse_lpi_1_dfm_1
      & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_12_and_110_cse = (~ return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse)
      & and_dcpl_501 & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_12_and_113_cse = (~ or_dcpl_711) &
      (fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_12_and_115_cse = (~ return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse)
      & return_add_generic_AC_RND_CONV_false_12_and_106_m1c;
  assign return_add_generic_AC_RND_CONV_false_12_and_117_cse = (~ return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse)
      & return_add_generic_AC_RND_CONV_false_12_and_108_m1c;
  assign return_add_generic_AC_RND_CONV_false_12_and_116_cse = return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse
      & return_add_generic_AC_RND_CONV_false_12_and_106_m1c;
  assign return_add_generic_AC_RND_CONV_false_12_and_118_cse = return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse
      & return_add_generic_AC_RND_CONV_false_12_and_108_m1c;
  assign return_add_generic_AC_RND_CONV_false_12_and_119_cse = (~ or_547_cse) & return_add_generic_AC_RND_CONV_false_12_and_114_m1c;
  assign return_add_generic_AC_RND_CONV_false_12_and_120_cse = or_547_cse & return_add_generic_AC_RND_CONV_false_12_and_114_m1c;
  assign return_add_generic_AC_RND_CONV_false_12_do_sub_mux1h_1_cse = ~((out_f_d_rsci_q_d[63])
      ^ (stage_PE_1_tmp_re_d_sva[63]));
  assign return_add_generic_AC_RND_CONV_false_12_do_sub_mux1h_6_cse = ~((in_f_d_rsci_q_d[63])
      ^ (stage_PE_1_tmp_re_d_sva[63]));
  assign return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse = (fsm_output[5])
      | (fsm_output[7]) | (fsm_output[30]) | (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_10_r_zero_or_2_cse = (fsm_output[18])
      | (fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_10_r_zero_or_3_cse = return_add_generic_AC_RND_CONV_false_10_r_zero_or_2_cse
      | (fsm_output[45]);
  assign return_extract_19_and_cse = return_extract_19_return_extract_19_nor_tmp
      & return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp;
  assign return_extract_51_and_cse = return_extract_51_return_extract_51_nor_tmp
      & return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp;
  assign return_add_generic_AC_RND_CONV_false_5_e_dif_sat_or_2_nl = (return_add_generic_AC_RND_CONV_false_4_e_dif_qif_acc_pmx_lpi_3_dfm_mx0_9_0[9:6]!=4'b0000)
      | ((return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt[10]) & (return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp[10]));
  assign operator_6_false_17_mux1h_cse_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_4_e_dif_qif_acc_pmx_lpi_3_dfm_mx0_9_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_5_e_dif_sat_or_2_nl);
  assign operator_6_false_17_or_cse = (fsm_output[10]) | (fsm_output[35]);
  assign operator_6_false_17_or_8_cse = or_dcpl_553 | (fsm_output[14]) | or_dcpl_493
      | (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse = (fsm_output[9])
      | (fsm_output[34]);
  assign return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_ssc = run_wen & (~(or_dcpl_627
      | or_dcpl_625 | (fsm_output[17]) | (fsm_output[35]) | (fsm_output[10]) | or_dcpl_484));
  assign return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_1_cse = (~ return_add_generic_AC_RND_CONV_false_17_acc_3_itm_10)
      & return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse;
  assign return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_4_cse = (return_add_generic_AC_RND_CONV_false_17_acc_3_itm_10
      & return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse) | (return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1
      & (fsm_output[11]));
  assign return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_4_cse = (~ return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1)
      & (fsm_output[11]);
  assign return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_5_cse = (~ return_add_generic_AC_RND_CONV_false_19_acc_2_itm_11_1)
      & (fsm_output[36]);
  assign return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_6_cse = return_add_generic_AC_RND_CONV_false_19_acc_2_itm_11_1
      & (fsm_output[36]);
  assign return_add_generic_AC_RND_CONV_false_10_ls_or_2_cse = (fsm_output[14]) |
      (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_10_ls_or_cse = (fsm_output[11]) | (fsm_output[12])
      | (fsm_output[13]) | (fsm_output[36]) | (fsm_output[37]) | (fsm_output[38]);
  assign and_6_cse = (~ mode_lpi_1_dfm) & inverse_lpi_1_dfm_1;
  assign or_32_cse = (~ mode_lpi_1_dfm) | inverse_lpi_1_dfm_1;
  assign operator_6_false_7_or_rgt = (fsm_output[10]) | (fsm_output[34]);
  assign and_2393_rgt = return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp
      & (fsm_output[13]);
  assign and_2395_rgt = (~ return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp)
      & (fsm_output[13]);
  assign and_2407_rgt = return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp
      & (fsm_output[38]);
  assign and_2409_rgt = (~ return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp)
      & (fsm_output[38]);
  assign return_extract_22_or_2_cse = and_2185_cse | and_2184_cse;
  assign and_38_nl = return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 &
      mux_tmp_22;
  assign mux_23_nl = MUX_s_1_2_2(and_38_nl, and_tmp_1, return_extract_19_and_cse);
  assign or_70_nl = (~ (z_out_68[12])) | operator_11_true_19_operator_11_true_19_and_tmp;
  assign mux_24_nl = MUX_s_1_2_2(mux_23_nl, and_tmp_1, or_70_nl);
  assign return_add_generic_AC_RND_CONV_false_10_res_rounded_and_cse = run_wen &
      (~ mux_24_nl) & mode_lpi_1_dfm;
  assign return_add_generic_AC_RND_CONV_false_11_or_4_cse = (fsm_output[16]) | (fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_11_or_5_cse = (fsm_output[30]) | (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_11_and_9_itm = return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1
      & return_add_generic_AC_RND_CONV_false_11_or_5_cse;
  assign and_528_cse = return_add_generic_AC_RND_CONV_false_9_e1_eq_e2_equal_tmp
      & z_out_53_52;
  assign or_673_cse = and_528_cse | (z_out_69[11]);
  assign nl_return_add_generic_AC_RND_CONV_false_18_ma1_lt_ma2_acc_2_nl = ({1'b1
      , (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[51:0])}) + conv_u2u_52_53(~
      (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[51:0])) +
      53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_18_ma1_lt_ma2_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_18_ma1_lt_ma2_acc_2_nl[52:0];
  assign and_526_cse = return_add_generic_AC_RND_CONV_false_17_e1_eq_e2_equal_tmp
      & (readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_18_ma1_lt_ma2_acc_2_nl));
  assign or_658_cse = and_526_cse | (return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp[10]);
  assign and_1251_cse = or_673_cse & (fsm_output[16]);
  assign operator_14_false_1_or_cse = (fsm_output[11]) | (fsm_output[12]) | (fsm_output[36])
      | (fsm_output[37]);
  assign return_add_generic_AC_RND_CONV_false_12_res_mant_and_ssc = run_wen & (~(or_dcpl_605
      | (fsm_output[49]) | or_dcpl_209 | or_dcpl_725 | (fsm_output[24]) | or_dcpl_236));
  assign or_1997_cse = (~ return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp)
      | (z_out_85[11]);
  assign return_add_generic_AC_RND_CONV_false_4_or_nl = return_add_generic_AC_RND_CONV_false_11_op_smaller_and_3_cse
      | return_add_generic_AC_RND_CONV_false_12_and_95_cse | return_add_generic_AC_RND_CONV_false_12_and_103_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_2_nl = return_add_generic_AC_RND_CONV_false_12_and_96_cse
      | return_add_generic_AC_RND_CONV_false_12_and_104_cse;
  assign return_add_generic_AC_RND_CONV_false_12_res_mant_mux1h_1_itm = MUX1HOT_v_56_3_2((~
      (z_out_76[56:1])), (z_out_76[56:1]), (~ (z_out_76[56:1])), {return_add_generic_AC_RND_CONV_false_11_op_smaller_and_4_cse
      , return_add_generic_AC_RND_CONV_false_4_or_nl , return_add_generic_AC_RND_CONV_false_4_or_2_nl});
  assign nand_133_cse = ~(return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp
      & (~ (z_out_85[11])));
  assign and_572_tmp = or_dcpl_284 & (~ operator_11_true_return_1_sva) & and_dcpl_503;
  assign and_577_tmp = (~(nand_133_cse & return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1))
      & (~(return_add_generic_AC_RND_CONV_false_2_if_5_return_add_generic_AC_RND_CONV_false_2_if_5_and_tmp
      & (z_out_89[53]))) & and_dcpl_285 & and_dcpl_64;
  assign and_582_tmp = or_dcpl_854 & (~((z_out_89[53]) & return_add_generic_AC_RND_CONV_false_3_if_5_return_add_generic_AC_RND_CONV_false_3_if_5_and_tmp))
      & and_dcpl_223 & and_dcpl_57;
  assign and_584_tmp = or_dcpl_342 & (~ operator_11_true_return_1_sva) & and_dcpl_503;
  assign and_588_tmp = (~(nand_133_cse & return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1))
      & (~((z_out_89[53]) & return_add_generic_AC_RND_CONV_false_15_if_5_return_add_generic_AC_RND_CONV_false_15_if_5_and_tmp))
      & and_dcpl_223 & and_dcpl_64;
  assign and_591_tmp = or_dcpl_854 & (~((z_out_89[53]) & return_add_generic_AC_RND_CONV_false_16_if_5_return_add_generic_AC_RND_CONV_false_16_if_5_and_tmp))
      & and_dcpl_285 & and_dcpl_57;
  assign and_276_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_1_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign and_311_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_14_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_10_op2_nan_and_cse = run_wen & (~(or_dcpl_809
      | (fsm_output[48]) | (fsm_output[23]) | (fsm_output[25]) | (fsm_output[24])
      | (fsm_output[17]) | (fsm_output[7]) | or_dcpl_269));
  assign return_add_generic_AC_RND_CONV_false_18_and_1_ssc = run_wen & (~(or_dcpl_586
      | or_dcpl_870));
  assign and_2325_rgt = return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp
      & (fsm_output[10]);
  assign and_2327_rgt = (~ return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp)
      & (fsm_output[10]);
  assign and_2339_rgt = return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp
      & (fsm_output[35]);
  assign and_2341_rgt = (~ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp)
      & (fsm_output[35]);
  assign return_add_generic_AC_RND_CONV_false_23_op1_mu_and_cse = run_wen & (~(or_dcpl_590
      | or_dcpl_933 | (fsm_output[9]) | or_dcpl_584 | or_dcpl_511 | (fsm_output[30])
      | (fsm_output[36]) | (fsm_output[40]) | or_dcpl_509 | or_dcpl_466 | (fsm_output[12])
      | or_dcpl_744));
  assign nl_return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl = ({1'b1 ,
      (out_f_d_rsci_q_d[51:0])}) + conv_u2u_52_53(~ (stage_PE_1_tmp_re_d_sva[51:0]))
      + 53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl[52:0];
  assign return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_and_1_cse
      = (readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl))
      & return_add_generic_AC_RND_CONV_false_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_and_1_cse
      | (z_out_69[11]);
  assign and_597_m1c = or_dcpl_967 & inverse_lpi_1_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_11_and_12_m1c = or_dcpl_980 & (fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_11_and_14_m1c = or_dcpl_981 & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_11_and_16_m1c = or_dcpl_982 & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_11_and_11_cse = (~ or_dcpl_980) & (fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_11_and_13_cse = (~ or_dcpl_981) & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_11_and_15_cse = (~ or_dcpl_982) & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_11_and_10_cse = (~ inverse_lpi_1_dfm_1)
      & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_11_and_19_cse = (~ return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse)
      & return_add_generic_AC_RND_CONV_false_11_and_14_m1c;
  assign return_add_generic_AC_RND_CONV_false_11_and_21_cse = (~ or_1102_cse) & return_add_generic_AC_RND_CONV_false_11_and_16_m1c;
  assign return_add_generic_AC_RND_CONV_false_11_and_17_cse = (~ or_673_cse) & return_add_generic_AC_RND_CONV_false_11_and_12_m1c;
  assign return_add_generic_AC_RND_CONV_false_11_and_18_cse = or_673_cse & return_add_generic_AC_RND_CONV_false_11_and_12_m1c;
  assign return_add_generic_AC_RND_CONV_false_11_and_20_cse = return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse
      & return_add_generic_AC_RND_CONV_false_11_and_14_m1c;
  assign return_add_generic_AC_RND_CONV_false_11_and_22_cse = or_1102_cse & return_add_generic_AC_RND_CONV_false_11_and_16_m1c;
  assign return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_and_1_cse
      = z_out_54_52 & return_add_generic_AC_RND_CONV_false_14_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_and_1_cse
      | (z_out_95[11]);
  assign return_add_generic_AC_RND_CONV_false_16_and_2_m1c = or_dcpl_967 & (fsm_output[7]);
  assign stage_PE_1_tmp_re_d_and_1_cse = run_wen & (~(return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse
      | or_dcpl_484));
  assign return_add_generic_AC_RND_CONV_false_12_r_zero_or_1_cse = (fsm_output[19])
      | (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1 = return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_1_mux_28);
  assign return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_tmp
      = ~((z_out_84[11:0]==12'b011111111111));
  assign return_add_generic_AC_RND_CONV_false_2_if_5_return_add_generic_AC_RND_CONV_false_2_if_5_nor_cse
      = ~((z_out_85!=13'b0000000000000));
  assign return_add_generic_AC_RND_CONV_false_2_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1
      | return_add_generic_AC_RND_CONV_false_2_if_5_return_add_generic_AC_RND_CONV_false_2_if_5_nor_cse;
  assign return_add_generic_AC_RND_CONV_false_2_mux_9_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1,
      return_add_generic_AC_RND_CONV_false_2_if_5_or_1_nl, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0 = return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_2_mux_9_nl);
  assign return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp
      = ~((z_out_85[11:0]==12'b011111111111));
  assign return_add_generic_AC_RND_CONV_false_3_if_5_or_2_nl = return_add_generic_AC_RND_CONV_false_16_acc_3_itm_11_1
      | (~((operator_33_true_32_acc_tmp!=13'b0000000000000)));
  assign return_add_generic_AC_RND_CONV_false_3_mux_17_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_16_acc_3_itm_11_1,
      return_add_generic_AC_RND_CONV_false_3_if_5_or_2_nl, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs_mx0w0 = return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_3_mux_17_nl);
  assign return_add_generic_AC_RND_CONV_false_16_else_4_return_add_generic_AC_RND_CONV_false_16_else_4_nand_tmp
      = ~((operator_33_true_32_acc_tmp[11:0]==12'b011111111111));
  assign return_add_generic_AC_RND_CONV_false_6_mux_33_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva,
      return_add_generic_AC_RND_CONV_false_1_if_5_or_3, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1 = return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_6_mux_33_nl);
  assign return_add_generic_AC_RND_CONV_false_4_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva
      | return_add_generic_AC_RND_CONV_false_18_if_5_return_add_generic_AC_RND_CONV_false_18_if_5_nor_2;
  assign return_add_generic_AC_RND_CONV_false_4_mux_15_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva,
      return_add_generic_AC_RND_CONV_false_4_if_5_or_1_nl, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_or_svs_mx0w0 = return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_4_mux_15_nl);
  assign return_add_generic_AC_RND_CONV_false_5_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva
      | return_add_generic_AC_RND_CONV_false_17_if_5_return_add_generic_AC_RND_CONV_false_17_if_5_nor_2;
  assign return_add_generic_AC_RND_CONV_false_5_mux_9_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva,
      return_add_generic_AC_RND_CONV_false_5_if_5_or_1_nl, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qelse_or_svs_mx0w0 = return_add_generic_AC_RND_CONV_false_12_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_5_mux_9_nl);
  assign return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1 = return_add_generic_AC_RND_CONV_false_12_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_1_mux_28);
  assign return_add_generic_AC_RND_CONV_false_15_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1
      | return_add_generic_AC_RND_CONV_false_2_if_5_return_add_generic_AC_RND_CONV_false_2_if_5_nor_cse;
  assign return_add_generic_AC_RND_CONV_false_15_mux_9_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1,
      return_add_generic_AC_RND_CONV_false_15_if_5_or_1_nl, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs_mx0w0 = return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_15_mux_9_nl);
  assign return_add_generic_AC_RND_CONV_false_17_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva
      | return_add_generic_AC_RND_CONV_false_17_if_5_return_add_generic_AC_RND_CONV_false_17_if_5_nor_2;
  assign return_add_generic_AC_RND_CONV_false_17_mux_15_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva,
      return_add_generic_AC_RND_CONV_false_17_if_5_or_1_nl, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qelse_or_svs_mx0w0 = return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_17_mux_15_nl);
  assign return_add_generic_AC_RND_CONV_false_18_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva
      | return_add_generic_AC_RND_CONV_false_18_if_5_return_add_generic_AC_RND_CONV_false_18_if_5_nor_2;
  assign return_add_generic_AC_RND_CONV_false_18_mux_9_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva,
      return_add_generic_AC_RND_CONV_false_18_if_5_or_1_nl, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_svs_mx0w0 = return_add_generic_AC_RND_CONV_false_12_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_18_mux_9_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl = -operator_6_false_58_acc_psp_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl[11:0];
  assign return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1 = readslicef_12_1_11(return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl);
  assign return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w1 = return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_1_mux_28);
  assign operator_16_false_1_operator_16_false_1_and_mdf_sva_1 = (mode1_rsci_idat==16'b0000000000000001);
  assign operator_16_false_operator_16_false_nor_tmp = ~((mode1_rsci_idat!=16'b0000000000000000));
  assign t_in_10_0_lpi_1_dfm_1_10_mx0w0 = ~(operator_16_false_1_operator_16_false_1_and_mdf_sva_1
      | operator_16_false_operator_16_false_nor_tmp);
  assign mode_lpi_1_dfm_mx0w0 = operator_16_false_1_operator_16_false_1_and_mdf_sva_1
      | operator_16_false_operator_16_false_nor_tmp;
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_8 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_8,
      m_in_15_1_lpi_1_dfm_1_9, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_7 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_7,
      m_in_15_1_lpi_1_dfm_1_8, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_6 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_6,
      m_in_15_1_lpi_1_dfm_1_7, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_5 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_5,
      m_in_15_1_lpi_1_dfm_1_6, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_4 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_4,
      m_in_15_1_lpi_1_dfm_1_5, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_3 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_3,
      m_in_15_1_lpi_1_dfm_1_4, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_2 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_2,
      m_in_15_1_lpi_1_dfm_1_3, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_1 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_1,
      m_in_15_1_lpi_1_dfm_1_2, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_0 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_0,
      m_in_15_1_lpi_1_dfm_1_1, mode_lpi_1_dfm);
  assign stage_PE_1_and_1_tmp = mode_lpi_1_dfm & inverse_lpi_1_dfm_1;
  assign nl_for_i_3_0_sva_2 = for_i_3_0_sva + 4'b0001;
  assign for_i_3_0_sva_2 = nl_for_i_3_0_sva_2[3:0];
  assign return_extract_3_m_zero_sva_mx1w0 = ~((out_f_d_rsci_q_d[51:0]!=52'b0000000000000000000000000000000000000000000000000000));
  assign return_extract_56_m_zero_sva_mx2w0 = ~((in_f_d_rsci_q_d[51:0]!=52'b0000000000000000000000000000000000000000000000000000));
  assign nl_operator_33_true_13_acc_nl = conv_s2s_11_12(operator_6_false_13_acc_psp_sva_1[11:1])
      + 12'b000000000001;
  assign operator_33_true_13_acc_nl = nl_operator_33_true_13_acc_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_6_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      operator_33_true_13_acc_nl, return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1);
  assign nl_operator_33_true_39_acc_nl = conv_s2s_11_12(operator_6_false_42_acc_psp_sva_1[11:1])
      + 12'b000000000001;
  assign operator_33_true_39_acc_nl = nl_operator_33_true_39_acc_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_2 = MUX_v_12_2_2(12'b000000000000,
      operator_33_true_39_acc_nl, return_add_generic_AC_RND_CONV_false_19_acc_2_itm_11_1);
  assign BUTTERFLY_i_div_psp_sva_1 = div_9_u9_u16(BUTTERFLY_1_n_9_0_sva_8_0, {stage_PE_1_index_const_15_lpi_2_dfm
      , stage_PE_1_index_const_14_11_lpi_2_dfm_3 , stage_PE_1_index_const_14_11_lpi_2_dfm_2
      , stage_PE_1_index_const_14_11_lpi_2_dfm_1 , stage_PE_1_index_const_14_11_lpi_2_dfm_0
      , stage_PE_1_index_const_10_lpi_2_dfm , stage_PE_1_index_const_9_1_lpi_2_dfm_8
      , stage_PE_1_index_const_9_1_lpi_2_dfm_7 , stage_PE_1_index_const_9_1_lpi_2_dfm_6
      , stage_PE_1_index_const_9_1_lpi_2_dfm_5 , stage_PE_1_index_const_9_1_lpi_2_dfm_4
      , stage_PE_1_index_const_9_1_lpi_2_dfm_3 , stage_PE_1_index_const_9_1_lpi_2_dfm_2
      , stage_PE_1_index_const_9_1_lpi_2_dfm_1 , stage_PE_1_index_const_9_1_lpi_2_dfm_0
      , stage_PE_1_index_const_0_lpi_2_dfm});
  assign nl_BUTTERFLY_i_9_0_sva_1 = conv_u2u_9_10(BUTTERFLY_1_n_9_0_sva_8_0) + (z_out_104[9:0]);
  assign BUTTERFLY_i_9_0_sva_1 = nl_BUTTERFLY_i_9_0_sva_1[9:0];
  assign return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp
      = (out_f_d_rsci_q_d[62:52]!=11'b00000000000);
  assign return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0 = operator_11_true_return_1_sva
      & (~ return_extract_12_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp
      = (in_f_d_rsci_q_d[62:52]!=11'b00000000000);
  assign return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_mx2w0 = operator_11_true_return_21_sva
      & (~ return_extract_21_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0 = operator_11_true_return_1_sva
      & return_extract_12_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0 = operator_11_true_return_21_sva
      & return_extract_21_m_zero_sva;
  assign and_2172_cse = return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse
      & (fsm_output[7]);
  assign and_2173_cse = return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse
      & (fsm_output[32]);
  assign or_1864_ssc = and_2172_cse | and_2173_cse;
  assign or_1866_ssc = or_dcpl_485 | (fsm_output[41]) | or_dcpl_943 | or_dcpl_559
      | (fsm_output[15]) | or_dcpl_685 | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse;
  assign return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_8_nl
      = MUX_v_9_2_2(9'b000000000, (z_out_112[9:1]), return_add_generic_AC_RND_CONV_false_17_acc_3_itm_10);
  assign BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_1_9_1 = MUX1HOT_v_9_9_2((stage_PE_1_tmp_re_d_sva[61:53]),
      (out_f_d_rsci_q_d[61:53]), (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1[9:1]),
      return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_8_nl,
      (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1[9:1]),
      (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[9:1]),
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0, (in_f_d_rsci_q_d[61:53]), (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_1[9:1]),
      {or_1864_ssc , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
      , or_1866_ssc , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse ,
      (fsm_output[12]) , return_extract_22_or_2_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_32_cse
      , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse , (fsm_output[38])});
  assign return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_9_nl
      = (z_out_112[0]) & return_add_generic_AC_RND_CONV_false_17_acc_3_itm_10;
  assign BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_1_0 = MUX1HOT_s_1_9_2((stage_PE_1_tmp_re_d_sva[52]),
      (out_f_d_rsci_q_d[52]), (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1[0]),
      return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_9_nl,
      (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1[0]), (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[0]),
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1, (in_f_d_rsci_q_d[52]), (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_1[0]),
      {or_1864_ssc , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
      , or_1866_ssc , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse ,
      (fsm_output[12]) , return_extract_22_or_2_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_32_cse
      , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse , (fsm_output[38])});
  assign return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1 = (out_f_d_rsci_q_d[51])
      | return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm_mx1
      = MUX_s_1_2_2(stage_PE_tmp_re_d_1_lpi_3_dfm_51_mx0, stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50,
      return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm_mx3
      = MUX_s_1_2_2(stage_PE_1_tmp_im_d_1_lpi_3_dfm_51_mx1, stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50,
      return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_1 = (in_f_d_rsci_q_d[51])
      | return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp;
  assign drf_qr_lval_13_smx_0_lpi_3_dfm_mx3 = MUX_s_1_2_2(return_extract_44_return_extract_44_or_1_cse_sva_1,
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_51_mx1, return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp);
  assign operator_11_true_3_operator_11_true_3_and_tmp = (out_f_d_rsci_q_d[62:52]==11'b11111111111);
  assign return_add_generic_AC_RND_CONV_false_6_r_nan_and_2 = operator_11_true_return_22_sva
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva & return_add_generic_AC_RND_CONV_false_12_do_sub_sva;
  assign operator_11_true_35_operator_11_true_35_and_tmp = (in_f_d_rsci_q_d[62:52]==11'b11111111111);
  assign drf_qr_lval_1_smx_lpi_3_dfm_mx0 = MUX_v_11_2_2((out_f_d_rsci_q_d[62:52]),
      (stage_PE_1_tmp_re_d_sva[62:52]), and_dcpl_448);
  assign return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1 = (stage_PE_1_tmp_re_d_sva[63])
      ^ (out_f_d_rsci_q_d[63]);
  assign return_extract_41_return_extract_41_or_1_cse_sva_1 = (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[61:52]!=10'b0000000000);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_70,
      z_out_69, z_out_71_11);
  assign return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1 = (stage_PE_1_tmp_re_d_sva[0])
      & return_add_generic_AC_RND_CONV_false_10_unequal_tmp;
  assign return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1 = (out_f_d_rsci_q_d[0])
      & return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1, and_dcpl_448);
  assign return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0
      = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm,
      return_extract_2_mux_4_cse, and_dcpl_448);
  assign return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_0_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1, and_dcpl_448);
  assign return_add_generic_AC_RND_CONV_false_1_e1_eq_e2_equal_tmp = (stage_PE_1_tmp_re_d_sva[62:52])
      == (out_f_d_rsci_q_d[62:52]);
  assign return_add_generic_AC_RND_CONV_false_1_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_109[54]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_109[53]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_109[52]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_109[51]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_109[50]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_109[49]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_109[48]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_109[47]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_109[46]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_109[45]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_109[44]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_109[43]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_109[42]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_109[41]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_109[40]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_109[39]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_109[38]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_109[37]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_109[36]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_109[35]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_109[34]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_109[33]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_109[32]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_109[31]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_109[30]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_109[29]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_109[28]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_109[27]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_109[26]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_109[25]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_109[24]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_109[23]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_109[22]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_109[21]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_109[20]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_109[19]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_109[18]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_109[17]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_109[16]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_109[15]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_109[14]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_109[13]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_109[12]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_109[11]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_109[10]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_109[9]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_109[8]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_109[7]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_109[6]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_109[5]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_109[4]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_109[3]))) | (return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_109[2])));
  assign return_add_generic_AC_RND_CONV_false_3_e_dif_qr_lpi_3_dfm_mx0_10_0 = MUX_v_11_2_2((z_out_70[10:0]),
      (z_out_69[10:0]), z_out_70[11]);
  assign return_add_generic_AC_RND_CONV_false_3_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_107[54]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_107[53]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_107[52]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_107[51]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_107[50]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_107[49]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_107[48]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_107[47]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_107[46]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_107[45]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_107[44]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_107[43]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_107[42]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_107[41]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_107[40]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_107[39]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_107[38]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_107[37]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_107[36]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_107[35]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_107[34]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_107[33]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_107[32]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_107[31]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_107[30]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_107[29]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_107[28]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_107[27]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_107[26]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_107[25]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_107[24]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_107[23]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_107[22]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_107[21]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_107[20]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_107[19]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_107[18]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_107[17]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_107[16]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_107[15]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_107[14]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_107[13]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_107[12]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_107[11]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_107[10]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_107[9]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_107[8]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_107[7]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_107[6]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_107[5]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_107[4]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_107[3]))) | (return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_107[2])));
  assign return_add_generic_AC_RND_CONV_false_e_dif1_return_add_generic_AC_RND_CONV_false_e_dif1_and_cse
      = (z_out_69[11]) & (z_out_70[11]);
  assign return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_3_e_dif_qr_lpi_3_dfm_mx0_10_0[10:6]!=5'b00000)
      | return_add_generic_AC_RND_CONV_false_e_dif1_return_add_generic_AC_RND_CONV_false_e_dif1_and_cse;
  assign return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_cse = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_3_e_dif_qr_lpi_3_dfm_mx0_10_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_3_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_1_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_1_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_1_e_dif_sat_or_1_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt = ({1'b1 ,
      (~ (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[61:52]))}) + conv_u2s_10_11(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[61:52])
      + 11'b00000000001;
  assign return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt = nl_return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt[10:0];
  assign return_add_generic_AC_RND_CONV_false_4_e_dif_qif_acc_pmx_lpi_3_dfm_mx0_9_0
      = MUX_v_10_2_2((return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp[9:0]),
      (return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt[9:0]), return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp[10]);
  assign nl_return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp = ({1'b1 , (~ (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[61:52]))})
      + conv_u2s_10_11(BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[61:52])
      + 11'b00000000001;
  assign return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp = nl_return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp[10:0];
  assign return_add_generic_AC_RND_CONV_false_4_op1_mu_52_lpi_3_dfm_1 = (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[51])
      | return_add_generic_AC_RND_CONV_false_4_unequal_tmp_1;
  assign stage_PE_gm_re_d_mux_cse = MUX_v_51_2_2((BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[50:0]),
      (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[51:1]), return_add_generic_AC_RND_CONV_false_4_unequal_tmp_1);
  assign return_add_generic_AC_RND_CONV_false_4_op1_mu_0_lpi_3_dfm_1 = (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[0])
      & return_add_generic_AC_RND_CONV_false_4_unequal_tmp_1;
  assign stage_PE_gm_im_d_mux_cse = MUX_s_1_2_2(return_extract_41_return_extract_41_or_1_cse_sva_1,
      (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[51]), return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_if_1_return_add_generic_AC_RND_CONV_false_17_op2_normal_return_extract_41_nor_tmp);
  assign stage_PE_gm_im_d_mux_2_cse = MUX_v_51_2_2((r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[51:1]),
      (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[50:0]), return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_if_1_return_add_generic_AC_RND_CONV_false_17_op2_normal_return_extract_41_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_4_op2_mu_0_lpi_3_dfm_1 = (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[0])
      & (~ return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_if_1_return_add_generic_AC_RND_CONV_false_17_op2_normal_return_extract_41_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_17_e1_eq_e2_equal_tmp = (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[61:52])
      == (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[61:52]);
  assign return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_if_1_return_add_generic_AC_RND_CONV_false_17_op2_normal_return_extract_41_nor_tmp
      = ~((r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[61:52]!=10'b0000000000));
  assign return_add_generic_AC_RND_CONV_false_4_unequal_tmp_1 = (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[61:52]!=10'b0000000000);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm_mx1w0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_4_op2_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_4_op1_mu_0_lpi_3_dfm_1, and_dcpl_460);
  assign return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm_mx1w0 = MUX_s_1_2_2(stage_PE_gm_im_d_mux_cse,
      return_add_generic_AC_RND_CONV_false_4_op1_mu_52_lpi_3_dfm_1, and_dcpl_460);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx1w0
      = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_4_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_4_op2_mu_0_lpi_3_dfm_1, and_dcpl_460);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1,
      and_dcpl_341);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx3 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1,
      and_dcpl_340);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx1w0
      = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_4_op1_mu_52_lpi_3_dfm_1,
      stage_PE_gm_im_d_mux_cse, and_dcpl_460);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx2 =
      MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[50]),
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0, and_dcpl_341);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx4 =
      MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[50]),
      return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0, and_dcpl_340);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx1 =
      MUX_s_1_2_2(return_extract_12_return_extract_12_or_1_cse_sva_1, stage_PE_tmp_re_d_1_lpi_3_dfm_51_mx0,
      return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx2 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_23_op1_mu_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0,
      and_dcpl_341);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx3 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm, or_547_cse);
  assign return_extract_12_return_extract_12_or_1_cse_sva_1 = (drf_qr_lval_10_smx_lpi_3_dfm_mx3_10_1!=10'b0000000000)
      | drf_qr_lval_10_smx_lpi_3_dfm_mx3_0;
  assign and_543_nl = and_dcpl_475 & (~(return_add_generic_AC_RND_CONV_false_10_op2_inf_sva
      | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva | return_add_generic_AC_RND_CONV_false_10_do_sub_sva));
  assign BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx2 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_do_sub_sva,
      (z_out_87[51]), and_543_nl);
  assign return_extract_44_return_extract_44_or_1_cse_sva_1 = (drf_qr_lval_10_smx_lpi_3_dfm_mx7_10_1!=10'b0000000000)
      | drf_qr_lval_10_smx_lpi_3_dfm_mx7_0;
  assign and_548_nl = and_dcpl_479 & (~ return_add_generic_AC_RND_CONV_false_17_mux_6_itm)
      & and_dcpl_478;
  assign BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx5 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_do_sub_sva,
      (z_out_87[51]), and_548_nl);
  assign return_extract_32_mux_cse = MUX_v_11_2_2((in_f_d_rsci_q_d[62:52]), (stage_PE_1_tmp_re_d_sva[62:52]),
      and_dcpl_452);
  assign drf_qr_lval_10_smx_lpi_3_dfm_mx2 = MUX_v_11_2_2((stage_PE_1_tmp_re_d_sva[62:52]),
      (out_f_d_rsci_q_d[62:52]), and_dcpl_466);
  assign drf_qr_lval_10_smx_lpi_3_dfm_mx3_10_1 = MUX_v_10_2_2((out_f_d_rsci_q_d[62:53]),
      return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0, inverse_lpi_1_dfm_1);
  assign drf_qr_lval_10_smx_lpi_3_dfm_mx3_0 = MUX_s_1_2_2((out_f_d_rsci_q_d[52]),
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm,
      inverse_lpi_1_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_1 =
      MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_2_10_0_1,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_4_lor_lpi_3_dfm_1);
  assign drf_qr_lval_10_smx_lpi_3_dfm_mx6 = MUX_v_11_2_2((stage_PE_1_tmp_re_d_sva[62:52]),
      (in_f_d_rsci_q_d[62:52]), and_dcpl_468);
  assign drf_qr_lval_10_smx_lpi_3_dfm_mx7_10_1 = MUX_v_10_2_2((in_f_d_rsci_q_d[62:53]),
      return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0, inverse_lpi_1_dfm_1);
  assign drf_qr_lval_10_smx_lpi_3_dfm_mx7_0 = MUX_s_1_2_2((in_f_d_rsci_q_d[52]),
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm,
      inverse_lpi_1_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1 = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_2_10_0_1,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_3_lor_lpi_3_dfm_1);
  assign nl_return_add_generic_AC_RND_CONV_false_1_acc_2_nl = -(z_out_84[11:0]);
  assign return_add_generic_AC_RND_CONV_false_1_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_1_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_1_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_1_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_acc_2_nl = -(z_out_84[11:0]);
  assign return_add_generic_AC_RND_CONV_false_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_6_acc_2_nl = -(operator_33_true_12_acc_tmp[11:0]);
  assign return_add_generic_AC_RND_CONV_false_6_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_6_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_6_acc_2_nl);
  assign return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp
      = (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_1!=11'b00000000000);
  assign nl_return_add_generic_AC_RND_CONV_false_9_acc_2_nl = -(z_out_85[11:0]);
  assign return_add_generic_AC_RND_CONV_false_9_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_9_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_9_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_9_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_10_acc_2_nl = -(z_out_85[11:0]);
  assign return_add_generic_AC_RND_CONV_false_10_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_10_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_10_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_10_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_11_acc_2_nl = -(z_out_85[11:0]);
  assign return_add_generic_AC_RND_CONV_false_11_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_11_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_11_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_12_acc_2_nl = -(z_out_85[11:0]);
  assign return_add_generic_AC_RND_CONV_false_12_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_12_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_12_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_12_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_14_acc_2_nl = -(z_out_84[11:0]);
  assign return_add_generic_AC_RND_CONV_false_14_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_14_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_14_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_14_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_13_acc_2_nl = -(z_out_84[11:0]);
  assign return_add_generic_AC_RND_CONV_false_13_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_13_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_13_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_13_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_19_acc_2_nl = -(operator_33_true_38_acc_tmp[11:0]);
  assign return_add_generic_AC_RND_CONV_false_19_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_19_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_19_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_19_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_22_acc_2_nl = -(z_out_85[11:0]);
  assign return_add_generic_AC_RND_CONV_false_22_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_22_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_22_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_22_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_23_acc_2_nl = -(z_out_85[11:0]);
  assign return_add_generic_AC_RND_CONV_false_23_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_23_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_23_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_24_acc_2_nl = -(z_out_85[11:0]);
  assign return_add_generic_AC_RND_CONV_false_24_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_24_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_24_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_25_acc_2_nl = -(z_out_85[11:0]);
  assign return_add_generic_AC_RND_CONV_false_25_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_25_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_25_acc_2_nl);
  assign return_mult_generic_AC_RND_CONV_false_1_op1_zero_sva_1 = operator_11_true_return_21_sva
      & return_extract_12_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_8_if_2_return_add_generic_AC_RND_CONV_false_8_if_2_and_1_mx2w0
      = stage_d_mul_return_d_2_63_sva & stage_PE_1_tmp_re_d_1_lpi_3_dfm_63;
  assign return_add_generic_AC_RND_CONV_false_8_ma1_lt_ma2_mux_5_nl = MUX_s_1_2_2((~
      return_mult_generic_AC_RND_CONV_false_2_m_r_51_lpi_3_dfm_mx1), (~ return_mult_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_mx1),
      fsm_output[39]);
  assign nl_acc_3_nl = ({1'b1 , BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm
      , return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm
      , 1'b1}) + conv_u2u_53_54({return_add_generic_AC_RND_CONV_false_8_ma1_lt_ma2_mux_5_nl
      , (~ return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1) , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[53:0];
  assign return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_and_cse
      = (readslicef_54_1_53(acc_3_nl)) & return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_8_op1_smaller_return_add_generic_AC_RND_CONV_false_8_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp[11]);
  assign return_add_generic_AC_RND_CONV_false_8_r_sign_mux_1_cse = MUX_s_1_2_2(stage_PE_1_tmp_re_d_1_lpi_3_dfm_63,
      stage_d_mul_return_d_2_63_sva, return_add_generic_AC_RND_CONV_false_8_op1_smaller_return_add_generic_AC_RND_CONV_false_8_op1_smaller_or_cse);
  assign nand_128_nl = ~(return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm , return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm
      , return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_49_0 , return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_7_mux_27_cse
      , return_extract_21_mux_cse , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1})));
  assign return_add_generic_AC_RND_CONV_false_17_mux_6_itm_mx2 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_if_2_return_add_generic_AC_RND_CONV_false_8_if_2_and_1_mx2w0,
      return_add_generic_AC_RND_CONV_false_8_r_sign_mux_1_cse, nand_128_nl);
  assign return_add_generic_AC_RND_CONV_false_7_if_2_return_add_generic_AC_RND_CONV_false_7_if_2_and_1_mx4w0
      = stage_d_mul_return_d_2_63_sva & stage_d_mul_return_d_4_63_sva;
  assign return_add_generic_AC_RND_CONV_false_21_ma1_lt_ma2_mux_5_nl = MUX_s_1_2_2((~
      return_mult_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_mx1), (~ return_mult_generic_AC_RND_CONV_false_2_m_r_51_lpi_3_dfm_mx1),
      fsm_output[14]);
  assign nl_acc_2_nl = ({1'b1 , drf_qr_lval_15_smx_0_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm
      , 1'b1}) + conv_u2u_53_54({return_add_generic_AC_RND_CONV_false_21_ma1_lt_ma2_mux_5_nl
      , (~ return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1) , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[53:0];
  assign return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_and_cse
      = (readslicef_54_1_53(acc_2_nl)) & return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_21_op1_smaller_return_add_generic_AC_RND_CONV_false_21_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp[11]);
  assign return_add_generic_AC_RND_CONV_false_21_r_sign_mux_1_cse = MUX_s_1_2_2(stage_d_mul_return_d_4_63_sva,
      stage_d_mul_return_d_2_63_sva, return_add_generic_AC_RND_CONV_false_21_op1_smaller_return_add_generic_AC_RND_CONV_false_21_op1_smaller_or_cse);
  assign nand_129_nl = ~(return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm , return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm
      , return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_49_0 , return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_20_mux_27_cse
      , return_extract_21_mux_cse , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1})));
  assign return_add_generic_AC_RND_CONV_false_17_mux_6_itm_mx4 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_if_2_return_add_generic_AC_RND_CONV_false_7_if_2_and_1_mx4w0,
      return_add_generic_AC_RND_CONV_false_21_r_sign_mux_1_cse, nand_129_nl);
  assign return_add_generic_AC_RND_CONV_false_12_if_2_return_add_generic_AC_RND_CONV_false_12_if_2_nor_mx3w0
      = ~(return_add_generic_AC_RND_CONV_false_17_mux_6_itm | (~ (stage_PE_1_tmp_re_d_sva[63])));
  assign return_add_generic_AC_RND_CONV_false_11_if_2_return_add_generic_AC_RND_CONV_false_11_if_2_nor_mx5w0
      = ~(return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 | (~ (stage_PE_1_x_re_d_sva[63])));
  assign return_mult_generic_AC_RND_CONV_false_op2_zero_sva_1 = return_extract_15_return_extract_15_nor_tmp
      & return_extract_47_m_zero_return_extract_47_m_zero_nor_tmp;
  assign return_mult_generic_AC_RND_CONV_false_1_op2_zero_sva_1 = return_extract_17_return_extract_17_nor_tmp
      & return_extract_49_m_zero_return_extract_49_m_zero_nor_tmp;
  assign return_mult_generic_AC_RND_CONV_false_3_op2_zero_sva_1 = return_extract_47_return_extract_47_nor_tmp
      & return_extract_47_m_zero_return_extract_47_m_zero_nor_tmp;
  assign return_mult_generic_AC_RND_CONV_false_4_op2_zero_sva_1 = return_extract_49_return_extract_49_nor_tmp
      & return_extract_49_m_zero_return_extract_49_m_zero_nor_tmp;
  assign return_add_generic_AC_RND_CONV_false_6_do_sub_sva_1 = ~(stage_PE_1_tmp_re_d_1_lpi_3_dfm_63
      ^ stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0);
  assign return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1 = (stage_PE_1_tmp_re_d_sva[63])
      ^ (in_f_d_rsci_q_d[63]);
  assign return_add_generic_AC_RND_CONV_false_19_do_sub_sva_1 = ~(stage_PE_1_tmp_re_d_1_lpi_3_dfm_63
      ^ stage_PE_1_tmp_im_d_1_lpi_3_dfm_63_mx0);
  assign nand_130_nl = ~(return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm
      , return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0 , return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_7_mux_27_cse
      , return_extract_21_mux_cse , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1})));
  assign return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_if_2_return_add_generic_AC_RND_CONV_false_7_if_2_and_1_mx4w0,
      return_add_generic_AC_RND_CONV_false_21_r_sign_mux_1_cse, nand_130_nl);
  assign nand_131_nl = ~(return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp
      & (({drf_qr_lval_13_smx_0_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm
      , return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0 , return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_20_mux_27_cse
      , return_extract_21_mux_cse , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1})));
  assign return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_if_2_return_add_generic_AC_RND_CONV_false_8_if_2_and_1_mx2w0,
      return_add_generic_AC_RND_CONV_false_8_r_sign_mux_1_cse, nand_131_nl);
  assign return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp
      = ~((drf_qr_lval_10_smx_lpi_3_dfm_mx3_10_1!=10'b0000000000) | drf_qr_lval_10_smx_lpi_3_dfm_mx3_0);
  assign return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp
      = ~((drf_qr_lval_10_smx_lpi_3_dfm_mx7_10_1!=10'b0000000000) | drf_qr_lval_10_smx_lpi_3_dfm_mx7_0);
  assign return_add_generic_AC_RND_CONV_false_1_if_2_return_add_generic_AC_RND_CONV_false_1_if_2_and_1_mx0w0
      = (out_f_d_rsci_q_d[63]) & (stage_PE_1_tmp_re_d_sva[63]);
  assign return_add_generic_AC_RND_CONV_false_10_if_2_return_add_generic_AC_RND_CONV_false_10_if_2_and_1_mx3w0
      = return_add_generic_AC_RND_CONV_false_17_mux_6_itm & (stage_PE_1_tmp_re_d_sva[63]);
  assign return_add_generic_AC_RND_CONV_false_13_if_2_return_add_generic_AC_RND_CONV_false_13_if_2_and_1_mx4w1
      = (stage_PE_1_tmp_re_d_sva[63]) & (in_f_d_rsci_q_d[63]);
  assign return_add_generic_AC_RND_CONV_false_9_if_2_return_add_generic_AC_RND_CONV_false_9_if_2_and_1_mx5w0
      = return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 & (stage_PE_1_x_re_d_sva[63]);
  assign nl_operator_33_true_12_acc_tmp = conv_s2s_7_13({acc_18_cse_6_1 , (~ (rtn_out_2[0]))})
      + conv_u2s_11_13({drf_qr_lval_6_smx_lpi_3_dfm_mx0_10 , drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_1
      , drf_qr_lval_6_smx_lpi_3_dfm_mx0_0});
  assign operator_33_true_12_acc_tmp = nl_operator_33_true_12_acc_tmp[12:0];
  assign nl_operator_6_false_41_acc_nl = ({1'b1 , (~ (leading_sign_57_0_1_0_19_out_3[5:1]))})
      + 6'b000001;
  assign operator_6_false_41_acc_nl = nl_operator_6_false_41_acc_nl[5:0];
  assign nl_operator_33_true_38_acc_tmp = conv_s2s_7_13({operator_6_false_41_acc_nl
      , (~ (leading_sign_57_0_1_0_19_out_3[0]))}) + conv_u2s_11_13({drf_qr_lval_22_smx_lpi_3_dfm_mx0_10
      , drf_qr_lval_22_smx_lpi_3_dfm_mx0_9_1 , drf_qr_lval_22_smx_lpi_3_dfm_mx0_0});
  assign operator_33_true_38_acc_tmp = nl_operator_33_true_38_acc_tmp[12:0];
  assign return_add_generic_AC_RND_CONV_false_11_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_2_e_dif_qr_lpi_3_dfm_mx0_10_0[10:6]!=5'b00000)
      | return_add_generic_AC_RND_CONV_false_e_dif1_return_add_generic_AC_RND_CONV_false_e_dif1_and_cse;
  assign return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_2_e_dif_qr_lpi_3_dfm_mx0_10_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_11_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_24_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_24_e_dif_qr_lpi_3_dfm_mx0_10_0[10:6]!=5'b00000)
      | ((z_out_98[11]) & (z_out_96[11]));
  assign return_add_generic_AC_RND_CONV_false_24_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_24_e_dif_qr_lpi_3_dfm_mx0_10_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_24_e_dif_sat_or_1_nl);
  assign nl_stage_u_add_acc_1_itm_1 = conv_u2s_16_17({BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0
      , BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0 , BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1})
      + 17'b11100111111111111;
  assign stage_u_add_acc_1_itm_1 = nl_stage_u_add_acc_1_itm_1[16:0];
  assign return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm_mx1w0
      = MUX_v_51_2_2(stage_PE_gm_re_d_mux_cse, stage_PE_gm_im_d_mux_2_cse, and_dcpl_460);
  assign return_mult_generic_AC_RND_CONV_false_oelse_3_return_mult_generic_AC_RND_CONV_false_3_if_3_nor_nl
      = ~((~ return_mult_generic_AC_RND_CONV_false_1_zero_m_return_mult_generic_AC_RND_CONV_false_1_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_1_r_zero_return_mult_generic_AC_RND_CONV_false_1_r_zero_nor_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_3_lor_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (z_out_87[50:0]), return_mult_generic_AC_RND_CONV_false_oelse_3_return_mult_generic_AC_RND_CONV_false_3_if_3_nor_nl);
  assign return_mult_generic_AC_RND_CONV_false_1_oelse_3_return_mult_generic_AC_RND_CONV_false_4_if_3_nor_nl
      = ~((~ return_mult_generic_AC_RND_CONV_false_1_zero_m_return_mult_generic_AC_RND_CONV_false_1_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_1_r_zero_return_mult_generic_AC_RND_CONV_false_1_r_zero_nor_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_4_lor_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (z_out_87[50:0]), return_mult_generic_AC_RND_CONV_false_1_oelse_3_return_mult_generic_AC_RND_CONV_false_4_if_3_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_mx1w0 = MUX_v_51_2_2(stage_PE_gm_im_d_mux_2_cse,
      stage_PE_gm_re_d_mux_cse, and_dcpl_460);
  assign return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx1
      = MUX_v_51_2_2((out_f_d_rsci_q_d[50:0]), return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm,
      inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx2
      = MUX_v_51_2_2((in_f_d_rsci_q_d[50:0]), return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm,
      inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_1_e_r_qelse_not_5_nl = ~ return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1;
  assign return_add_generic_AC_RND_CONV_false_1_e_r_qelse_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(10'b0000000000,
      z_out_90, return_add_generic_AC_RND_CONV_false_1_e_r_qelse_not_5_nl);
  assign return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_5_cse
      = MUX_v_12_2_2(12'b000000000000, z_out_114, return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva);
  assign return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_2_cse
      = (z_out_94[0]) | (~ return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva);
  assign return_add_generic_AC_RND_CONV_false_1_if_5_or_nl = and_276_cse | return_add_generic_AC_RND_CONV_false_if_5_return_add_generic_AC_RND_CONV_false_if_5_and_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_1_mux_16_nl = MUX_s_1_2_2(and_276_cse,
      return_add_generic_AC_RND_CONV_false_1_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_1_exception_sva_1 = return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0
      | return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0 | return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_mx2w0 | return_add_generic_AC_RND_CONV_false_1_mux_16_nl;
  assign return_add_generic_AC_RND_CONV_false_4_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm
      & (~ (z_out_109[54]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[50])
      & (~ (z_out_109[53]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[49])
      & (~ (z_out_109[52]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[48])
      & (~ (z_out_109[51]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[47])
      & (~ (z_out_109[50]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[46])
      & (~ (z_out_109[49]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[45])
      & (~ (z_out_109[48]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[44])
      & (~ (z_out_109[47]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[43])
      & (~ (z_out_109[46]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[42])
      & (~ (z_out_109[45]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[41])
      & (~ (z_out_109[44]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[40])
      & (~ (z_out_109[43]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[39])
      & (~ (z_out_109[42]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[38])
      & (~ (z_out_109[41]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[37])
      & (~ (z_out_109[40]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[36])
      & (~ (z_out_109[39]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[35])
      & (~ (z_out_109[38]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[34])
      & (~ (z_out_109[37]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[33])
      & (~ (z_out_109[36]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[32])
      & (~ (z_out_109[35]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[31])
      & (~ (z_out_109[34]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[30])
      & (~ (z_out_109[33]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[29])
      & (~ (z_out_109[32]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[28])
      & (~ (z_out_109[31]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[27])
      & (~ (z_out_109[30]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[26])
      & (~ (z_out_109[29]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[25])
      & (~ (z_out_109[28]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[24])
      & (~ (z_out_109[27]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[23])
      & (~ (z_out_109[26]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[22])
      & (~ (z_out_109[25]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[21])
      & (~ (z_out_109[24]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[20])
      & (~ (z_out_109[23]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[19])
      & (~ (z_out_109[22]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[18])
      & (~ (z_out_109[21]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[17])
      & (~ (z_out_109[20]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[16])
      & (~ (z_out_109[19]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[15])
      & (~ (z_out_109[18]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[14])
      & (~ (z_out_109[17]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[13])
      & (~ (z_out_109[16]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[12])
      & (~ (z_out_109[15]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[11])
      & (~ (z_out_109[14]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[10])
      & (~ (z_out_109[13]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[9])
      & (~ (z_out_109[12]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[8])
      & (~ (z_out_109[11]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[7])
      & (~ (z_out_109[10]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[6])
      & (~ (z_out_109[9]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[5])
      & (~ (z_out_109[8]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[4])
      & (~ (z_out_109[7]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[3])
      & (~ (z_out_109[6]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[2])
      & (~ (z_out_109[5]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[1])
      & (~ (z_out_109[4]))) | ((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[0])
      & (~ (z_out_109[3]))) | return_add_generic_AC_RND_CONV_false_4_sticky_bit_and_158;
  assign return_add_generic_AC_RND_CONV_false_5_res_mant_3_0_sva_1 = (BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm
      & (~ (z_out_107[54]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[50])
      & (~ (z_out_107[53]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[49])
      & (~ (z_out_107[52]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[48])
      & (~ (z_out_107[51]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[47])
      & (~ (z_out_107[50]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[46])
      & (~ (z_out_107[49]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[45])
      & (~ (z_out_107[48]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[44])
      & (~ (z_out_107[47]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[43])
      & (~ (z_out_107[46]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[42])
      & (~ (z_out_107[45]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[41])
      & (~ (z_out_107[44]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[40])
      & (~ (z_out_107[43]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[39])
      & (~ (z_out_107[42]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[38])
      & (~ (z_out_107[41]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[37])
      & (~ (z_out_107[40]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[36])
      & (~ (z_out_107[39]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[35])
      & (~ (z_out_107[38]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[34])
      & (~ (z_out_107[37]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[33])
      & (~ (z_out_107[36]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[32])
      & (~ (z_out_107[35]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[31])
      & (~ (z_out_107[34]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[30])
      & (~ (z_out_107[33]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[29])
      & (~ (z_out_107[32]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[28])
      & (~ (z_out_107[31]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[27])
      & (~ (z_out_107[30]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[26])
      & (~ (z_out_107[29]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[25])
      & (~ (z_out_107[28]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[24])
      & (~ (z_out_107[27]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[23])
      & (~ (z_out_107[26]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[22])
      & (~ (z_out_107[25]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[21])
      & (~ (z_out_107[24]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[20])
      & (~ (z_out_107[23]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[19])
      & (~ (z_out_107[22]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[18])
      & (~ (z_out_107[21]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[17])
      & (~ (z_out_107[20]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[16])
      & (~ (z_out_107[19]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[15])
      & (~ (z_out_107[18]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[14])
      & (~ (z_out_107[17]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[13])
      & (~ (z_out_107[16]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[12])
      & (~ (z_out_107[15]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[11])
      & (~ (z_out_107[14]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[10])
      & (~ (z_out_107[13]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[9])
      & (~ (z_out_107[12]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[8])
      & (~ (z_out_107[11]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[7])
      & (~ (z_out_107[10]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[6])
      & (~ (z_out_107[9]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[5])
      & (~ (z_out_107[8]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[4])
      & (~ (z_out_107[7]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[3])
      & (~ (z_out_107[6]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[2])
      & (~ (z_out_107[5]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[1])
      & (~ (z_out_107[4]))) | ((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[0])
      & (~ (z_out_107[3]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm
      & (~ (z_out_107[2])));
  assign return_add_generic_AC_RND_CONV_false_6_r_nan_or_mx6w0 = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_6_r_nan_and_2;
  assign and_592_nl = and_dcpl_475 & and_dcpl_478;
  assign drf_qr_lval_15_smx_0_lpi_3_dfm_mx2 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_do_sub_sva,
      (z_out_87[51]), and_592_nl);
  assign return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 = operator_11_true_return_21_sva
      & (~ return_extract_12_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_14_op1_nan_sva_mx0w5 = operator_11_true_return_24_sva
      & (~ return_add_generic_AC_RND_CONV_false_12_mux_itm);
  assign return_add_generic_AC_RND_CONV_false_10_op1_nan_sva_mx0w9 = operator_11_true_return_26_sva
      & (~ return_extract_26_m_zero_sva);
  assign return_mult_generic_AC_RND_CONV_false_op2_inf_sva_1 = operator_11_true_15_operator_11_true_15_and_tmp
      & return_extract_47_m_zero_return_extract_47_m_zero_nor_tmp;
  assign return_mult_generic_AC_RND_CONV_false_1_op2_inf_sva_1 = operator_11_true_17_operator_11_true_17_and_tmp
      & return_extract_49_m_zero_return_extract_49_m_zero_nor_tmp;
  assign return_mult_generic_AC_RND_CONV_false_2_op2_inf_sva_1 = operator_11_true_19_operator_11_true_19_and_tmp
      & return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp;
  assign return_mult_generic_AC_RND_CONV_false_3_op2_inf_sva_1 = operator_11_true_47_operator_11_true_47_and_tmp
      & return_extract_47_m_zero_return_extract_47_m_zero_nor_tmp;
  assign return_mult_generic_AC_RND_CONV_false_4_op2_inf_sva_1 = operator_11_true_49_operator_11_true_49_and_tmp
      & return_extract_49_m_zero_return_extract_49_m_zero_nor_tmp;
  assign return_mult_generic_AC_RND_CONV_false_5_op2_inf_sva_1 = operator_11_true_51_operator_11_true_51_and_tmp
      & return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp;
  assign return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp
      = (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1!=11'b00000000000);
  assign return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1 = operator_11_true_return_1_sva
      & return_extract_21_m_zero_sva;
  assign nl_operator_6_false_7_acc_psp_sva_mx0w0 = conv_u2s_11_12(drf_qr_lval_19_smx_lpi_3_dfm)
      + conv_s2s_7_12({1'b1 , (~ rtn_out_2)}) + 12'b000000000001;
  assign operator_6_false_7_acc_psp_sva_mx0w0 = nl_operator_6_false_7_acc_psp_sva_mx0w0[11:0];
  assign nl_return_add_generic_AC_RND_CONV_false_e_dif_acc_1_nl = ({1'b1 , (out_f_d_rsci_q_d[62:52])})
      + conv_u2u_11_12(~ (stage_PE_1_tmp_re_d_sva[62:52])) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_e_dif_acc_1_nl = nl_return_add_generic_AC_RND_CONV_false_e_dif_acc_1_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_69,
      z_out_70, readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_e_dif_acc_1_nl));
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_0_lpi_3_dfm_1 = (stage_PE_1_tmp_re_d_sva[0])
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_op_smaller_qr_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1,
      drf_qr_lval_13_smx_0_lpi_3_dfm, and_dcpl_466);
  assign return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0 =
      MUX_v_51_2_2(return_extract_2_mux_4_cse, return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm,
      and_dcpl_466);
  assign return_add_generic_AC_RND_CONV_false_op_smaller_qr_0_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_0_lpi_3_dfm_1, and_dcpl_466);
  assign return_add_generic_AC_RND_CONV_false_e1_eq_e2_equal_tmp = (out_f_d_rsci_q_d[62:52])
      == (stage_PE_1_tmp_re_d_sva[62:52]);
  assign return_add_generic_AC_RND_CONV_false_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_109[54]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_109[53]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_109[52]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_109[51]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_109[50]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_109[49]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_109[48]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_109[47]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_109[46]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_109[45]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_109[44]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_109[43]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_109[42]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_109[41]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_109[40]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_109[39]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_109[38]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_109[37]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_109[36]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_109[35]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_109[34]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_109[33]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_109[32]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_109[31]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_109[30]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_109[29]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_109[28]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_109[27]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_109[26]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_109[25]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_109[24]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_109[23]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_109[22]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_109[21]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_109[20]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_109[19]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_109[18]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_109[17]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_109[16]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_109[15]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_109[14]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_109[13]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_109[12]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_109[11]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_109[10]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_109[9]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_109[8]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_109[7]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_109[6]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_109[5]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_109[4]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_109[3]))) | (return_add_generic_AC_RND_CONV_false_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_109[2])));
  assign return_add_generic_AC_RND_CONV_false_not_3_nl = ~ (z_out_88[53]);
  assign return_add_generic_AC_RND_CONV_false_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (z_out_88[51:0]), return_add_generic_AC_RND_CONV_false_not_3_nl);
  assign return_add_generic_AC_RND_CONV_false_2_e_dif_qr_lpi_3_dfm_mx0_10_0 = MUX_v_11_2_2((z_out_69[10:0]),
      (z_out_70[10:0]), z_out_69[11]);
  assign return_add_generic_AC_RND_CONV_false_2_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_107[54]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_107[53]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_107[52]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_107[51]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_107[50]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_107[49]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_107[48]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_107[47]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_107[46]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_107[45]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_107[44]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_107[43]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_107[42]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_107[41]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_107[40]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_107[39]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_107[38]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_107[37]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_107[36]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_107[35]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_107[34]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_107[33]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_107[32]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_107[31]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_107[30]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_107[29]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_107[28]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_107[27]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_107[26]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_107[25]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_107[24]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_107[23]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_107[22]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_107[21]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_107[20]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_107[19]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_107[18]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_107[17]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_107[16]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_107[15]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_107[14]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_107[13]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_107[12]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_107[11]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_107[10]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_107[9]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_107[8]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_107[7]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_107[6]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_107[5]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_107[4]))) | ((return_add_generic_AC_RND_CONV_false_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_107[3]))) | (return_add_generic_AC_RND_CONV_false_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_107[2])));
  assign return_add_generic_AC_RND_CONV_false_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_if_5_or_nl = and_281_cse | return_add_generic_AC_RND_CONV_false_if_5_return_add_generic_AC_RND_CONV_false_if_5_and_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_mux_16_nl = MUX_s_1_2_2(and_281_cse,
      return_add_generic_AC_RND_CONV_false_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_exception_sva_1 = return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0
      | return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0 | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_mx2w0
      | return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0 | return_add_generic_AC_RND_CONV_false_mux_16_nl;
  assign return_add_generic_AC_RND_CONV_false_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_6_exp_plus_1_0_lpi_3_dfm_1 = (operator_6_false_13_acc_psp_sva_1[0])
      | (~ return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_19_exp_plus_1_0_lpi_3_dfm_1 = (operator_6_false_42_acc_psp_sva_1[0])
      | (~ return_add_generic_AC_RND_CONV_false_19_acc_2_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1 = operator_11_true_return_1_sva
      & (~ return_extract_21_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_7_mux_27_cse = MUX_s_1_2_2((return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1[50]),
      return_mult_generic_AC_RND_CONV_false_2_m_r_51_lpi_3_dfm_mx1, return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp);
  assign return_extract_21_mux_cse = MUX_v_50_2_2((return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1[49:0]),
      (return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1[50:1]), return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp);
  assign return_add_generic_AC_RND_CONV_false_20_mux_27_cse = MUX_s_1_2_2((return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1[50]),
      return_mult_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_mx1, return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp);
  assign return_add_generic_AC_RND_CONV_false_2_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      z_out_103, return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_2_not_3_nl = ~ (z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (z_out_89[51:0]), return_add_generic_AC_RND_CONV_false_2_not_3_nl);
  assign return_add_generic_AC_RND_CONV_false_2_exp_plus_1_0_lpi_3_dfm_1 = (z_out_94[0])
      | (~ return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_2_if_5_return_add_generic_AC_RND_CONV_false_2_if_5_and_tmp
      = (return_add_generic_AC_RND_CONV_false_2_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_2_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_2_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_2_if_5_or_nl = return_add_generic_AC_RND_CONV_false_2_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_2_if_5_return_add_generic_AC_RND_CONV_false_2_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_2_mux_14_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_2_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_2_if_5_or_nl, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_2_exception_sva_1 = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      | operator_11_true_return_26_sva | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_unequal_tmp | return_add_generic_AC_RND_CONV_false_2_mux_14_nl;
  assign return_add_generic_AC_RND_CONV_false_2_r_inf_lpi_3_dfm_2 = or_1997_cse &
      return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_2_mux_4_itm = MUX_v_6_2_2((BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1[5:0]),
      return_add_generic_AC_RND_CONV_false_10_ls_sva, return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1);
  assign nl_operator_6_false_9_acc_psp_1_sva_1 = conv_u2s_10_11(operator_14_false_1_acc_psp_sva_9_0)
      + conv_s2s_7_11({1'b1 , (~ rtn_out_2)}) + 11'b00000000001;
  assign operator_6_false_9_acc_psp_1_sva_1 = nl_operator_6_false_9_acc_psp_1_sva_1[10:0];
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_51_mx0 = MUX_s_1_2_2((out_f_d_rsci_q_d[51]),
      drf_qr_lval_14_smx_0_lpi_3_dfm, inverse_lpi_1_dfm_1);
  assign nl_operator_33_true_32_acc_tmp = conv_s2s_7_13({operator_6_false_21_acc_itm_6_1
      , operator_6_false_21_acc_itm_0}) + conv_u2s_11_13(drf_qr_lval_19_smx_lpi_3_dfm);
  assign operator_33_true_32_acc_tmp = nl_operator_33_true_32_acc_tmp[12:0];
  assign return_add_generic_AC_RND_CONV_false_3_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      z_out_103, return_add_generic_AC_RND_CONV_false_16_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_3_exp_plus_1_0_lpi_3_dfm_1 = (operator_32_false_1_acc_psp_sva_11_0[0])
      | (~ return_add_generic_AC_RND_CONV_false_16_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_3_if_5_nor_cse = ~((return_add_generic_AC_RND_CONV_false_3_exp_plus_1_12_1_lpi_3_dfm_1[11:10]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_3_if_5_return_add_generic_AC_RND_CONV_false_3_if_5_and_tmp
      = (return_add_generic_AC_RND_CONV_false_3_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_3_exp_plus_1_0_lpi_3_dfm_1 & return_add_generic_AC_RND_CONV_false_3_if_5_nor_cse;
  assign return_add_generic_AC_RND_CONV_false_3_if_5_or_nl = return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_3_if_5_return_add_generic_AC_RND_CONV_false_3_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_3_mux_14_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_3_if_5_or_nl, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_3_exception_sva_1 = operator_11_true_return_22_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_3_mux_14_nl;
  assign return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2 = ((operator_33_true_32_acc_tmp[11])
      | (~ return_add_generic_AC_RND_CONV_false_16_else_4_return_add_generic_AC_RND_CONV_false_16_else_4_nand_tmp))
      & return_add_generic_AC_RND_CONV_false_16_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_3_mux_15_itm = MUX_v_6_2_2((drf_qr_lval_19_smx_lpi_3_dfm[5:0]),
      return_add_generic_AC_RND_CONV_false_11_ls_sva, return_add_generic_AC_RND_CONV_false_16_acc_3_itm_11_1);
  assign nl_operator_6_false_11_acc_psp_1_sva_1 = conv_u2s_10_11(drf_qr_lval_21_smx_9_0_lpi_3_dfm)
      + conv_s2s_7_11({1'b1 , (~ rtn_out_2)}) + 11'b00000000001;
  assign operator_6_false_11_acc_psp_1_sva_1 = nl_operator_6_false_11_acc_psp_1_sva_1[10:0];
  assign stage_d_mul_return_d_1_63_sva_1 = stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0 ^
      return_add_generic_AC_RND_CONV_false_18_mux_itm;
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_51_mx1 = MUX_s_1_2_2((in_f_d_rsci_q_d[51]),
      drf_qr_lval_14_smx_0_lpi_3_dfm, inverse_lpi_1_dfm_1);
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50 = MUX_s_1_2_2((out_f_d_rsci_q_d[50]),
      (return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[50]),
      inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_6_r_sign_mux_nl = MUX_s_1_2_2(stage_PE_1_tmp_re_d_1_lpi_3_dfm_63,
      (~ stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0), return_add_generic_AC_RND_CONV_false_6_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_nor_nl
      = ~(stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0 | (~ stage_PE_1_tmp_re_d_1_lpi_3_dfm_63));
  assign return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_and_nl
      = (({return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm
      , return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0 , return_add_generic_AC_RND_CONV_false_6_op1_mu_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx1
      , return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm_mx1
      , return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_49_0_mx0 , return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1}))
      & return_add_generic_AC_RND_CONV_false_6_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_6_mux_6_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_r_sign_mux_nl,
      return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_nor_nl,
      return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_and_nl);
  assign stage_d_mul_return_d_2_63_sva_1 = inverse_lpi_1_dfm_1 ^ return_add_generic_AC_RND_CONV_false_6_mux_6_nl;
  assign return_add_generic_AC_RND_CONV_false_19_r_sign_mux_nl = MUX_s_1_2_2(stage_PE_1_tmp_re_d_1_lpi_3_dfm_63,
      (~ stage_PE_1_tmp_im_d_1_lpi_3_dfm_63_mx0), return_add_generic_AC_RND_CONV_false_19_op1_smaller_lor_lpi_3_dfm_2);
  assign return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_nor_nl
      = ~(stage_PE_1_tmp_im_d_1_lpi_3_dfm_63_mx0 | (~ stage_PE_1_tmp_re_d_1_lpi_3_dfm_63));
  assign return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_and_nl
      = (({drf_qr_lval_13_smx_0_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm
      , return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0 , return_add_generic_AC_RND_CONV_false_6_op1_mu_0_lpi_3_dfm_1})
      == ({drf_qr_lval_13_smx_0_lpi_3_dfm_mx3 , return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm_mx3
      , return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0_mx0 ,
      return_add_generic_AC_RND_CONV_false_19_op2_mu_0_lpi_3_dfm_1})) & return_add_generic_AC_RND_CONV_false_19_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_19_mux_6_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_19_r_sign_mux_nl,
      return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_nor_nl,
      return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_and_nl);
  assign stage_d_mul_return_d_5_63_sva_1 = inverse_lpi_1_dfm_1 ^ return_add_generic_AC_RND_CONV_false_19_mux_6_nl;
  assign stage_d_mul_return_d_63_sva_1 = stage_PE_1_tmp_re_d_1_lpi_3_dfm_63 ^ return_add_generic_AC_RND_CONV_false_17_mux_6_itm;
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0 = MUX_s_1_2_2((out_f_d_rsci_q_d[63]),
      return_add_generic_AC_RND_CONV_false_12_mux_itm, inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_95,
      z_out_70, z_out_95[11]);
  assign return_add_generic_AC_RND_CONV_false_6_op1_mu_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[0])
      & (~ operator_11_true_return_21_sva);
  assign return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_49_0_mx0 =
      MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx1[50:1]),
      (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx1[49:0]),
      return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx1[0])
      & (~ return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp);
  assign drf_qr_lval_6_smx_lpi_3_dfm_mx0_10 = MUX_s_1_2_2((drf_qr_lval_10_smx_lpi_3_dfm_mx3_10_1[9]),
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_0, and_dcpl_531);
  assign drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_1 = MUX_v_9_2_2((drf_qr_lval_10_smx_lpi_3_dfm_mx3_10_1[8:0]),
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0, and_dcpl_531);
  assign drf_qr_lval_6_smx_lpi_3_dfm_mx0_0 = MUX_s_1_2_2(drf_qr_lval_10_smx_lpi_3_dfm_mx3_0,
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1, and_dcpl_531);
  assign return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx1, and_dcpl_531);
  assign return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_50_mx0
      = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm_mx1,
      and_dcpl_531);
  assign return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0
      = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0, return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_49_0_mx0,
      and_dcpl_531);
  assign return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_0_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1, and_dcpl_531);
  assign return_add_generic_AC_RND_CONV_false_6_e1_eq_e2_equal_tmp = ({drf_qr_lval_10_smx_lpi_3_dfm_rsp_0
      , drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0 , drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1})
      == ({drf_qr_lval_10_smx_lpi_3_dfm_mx3_10_1 , drf_qr_lval_10_smx_lpi_3_dfm_mx3_0});
  assign return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_and_cse
      = z_out_57_52 & return_add_generic_AC_RND_CONV_false_6_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_6_op1_smaller_lor_lpi_3_dfm_2 = return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_and_cse
      | (z_out_95[11]);
  assign return_add_generic_AC_RND_CONV_false_6_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_109[54]))) | (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_50_mx0
      & (~ (z_out_109[53]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[49])
      & (~ (z_out_109[52]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[48])
      & (~ (z_out_109[51]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[47])
      & (~ (z_out_109[50]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[46])
      & (~ (z_out_109[49]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[45])
      & (~ (z_out_109[48]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[44])
      & (~ (z_out_109[47]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[43])
      & (~ (z_out_109[46]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[42])
      & (~ (z_out_109[45]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[41])
      & (~ (z_out_109[44]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[40])
      & (~ (z_out_109[43]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[39])
      & (~ (z_out_109[42]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[38])
      & (~ (z_out_109[41]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[37])
      & (~ (z_out_109[40]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[36])
      & (~ (z_out_109[39]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[35])
      & (~ (z_out_109[38]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[34])
      & (~ (z_out_109[37]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[33])
      & (~ (z_out_109[36]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[32])
      & (~ (z_out_109[35]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[31])
      & (~ (z_out_109[34]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[30])
      & (~ (z_out_109[33]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[29])
      & (~ (z_out_109[32]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[28])
      & (~ (z_out_109[31]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[27])
      & (~ (z_out_109[30]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[26])
      & (~ (z_out_109[29]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[25])
      & (~ (z_out_109[28]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[24])
      & (~ (z_out_109[27]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[23])
      & (~ (z_out_109[26]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[22])
      & (~ (z_out_109[25]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[21])
      & (~ (z_out_109[24]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[20])
      & (~ (z_out_109[23]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[19])
      & (~ (z_out_109[22]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[18])
      & (~ (z_out_109[21]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[17])
      & (~ (z_out_109[20]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[16])
      & (~ (z_out_109[19]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[15])
      & (~ (z_out_109[18]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[14])
      & (~ (z_out_109[17]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[13])
      & (~ (z_out_109[16]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[12])
      & (~ (z_out_109[15]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[11])
      & (~ (z_out_109[14]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[10])
      & (~ (z_out_109[13]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[9])
      & (~ (z_out_109[12]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[8])
      & (~ (z_out_109[11]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[7])
      & (~ (z_out_109[10]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[6])
      & (~ (z_out_109[9]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[5])
      & (~ (z_out_109[8]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[4])
      & (~ (z_out_109[7]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[3])
      & (~ (z_out_109[6]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[2])
      & (~ (z_out_109[5]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[1])
      & (~ (z_out_109[4]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[0])
      & (~ (z_out_109[3]))) | (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_109[2])));
  assign return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1 = ~((z_out_86[9:6]==4'b1111));
  assign return_extract_15_return_extract_15_or_sva_1 = (return_add_generic_AC_RND_CONV_false_4_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_4_m_r_51_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1[51])
      & return_add_generic_AC_RND_CONV_false_4_if_7_not_4;
  assign return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_4_if_7_not_4);
  assign nor_182_cse = ~(MUX_v_10_2_2(z_out_91, 10'b1111111111, return_add_generic_AC_RND_CONV_false_17_if_5_return_add_generic_AC_RND_CONV_false_17_if_5_and_tmp));
  assign nor_179_nl = ~((~ return_add_generic_AC_RND_CONV_false_4_e_r_qelse_or_svs_mx0w0)
      | return_add_generic_AC_RND_CONV_false_17_if_5_return_add_generic_AC_RND_CONV_false_17_if_5_and_tmp);
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qr_10_1_lpi_3_dfm_1 = ~(MUX_v_10_2_2(nor_182_cse,
      10'b1111111111, nor_179_nl));
  assign return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_3_nl
      = (operator_33_true_36_acc_psp_1_sva[0]) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_4_mux_19_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_3_nl,
      operator_6_false_17_acc_itm_0, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_4_mux_19_nl
      & (~ return_add_generic_AC_RND_CONV_false_4_e_r_qelse_or_svs_mx0w0)) | return_add_generic_AC_RND_CONV_false_17_if_5_return_add_generic_AC_RND_CONV_false_17_if_5_and_tmp;
  assign return_extract_15_return_extract_15_nor_tmp = ~((return_add_generic_AC_RND_CONV_false_4_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1);
  assign operator_11_true_15_operator_11_true_15_and_tmp = (return_add_generic_AC_RND_CONV_false_4_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1;
  assign return_extract_47_m_zero_return_extract_47_m_zero_nor_tmp = ~(return_add_generic_AC_RND_CONV_false_4_m_r_51_lpi_3_dfm_1
      | (return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign nl_operator_6_false_13_acc_psp_sva_1 = conv_u2s_11_12({drf_qr_lval_6_smx_lpi_3_dfm_mx0_10
      , drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_1 , drf_qr_lval_6_smx_lpi_3_dfm_mx0_0})
      + conv_s2s_7_12({1'b1 , (~ rtn_out_2)}) + 12'b000000000001;
  assign operator_6_false_13_acc_psp_sva_1 = nl_operator_6_false_13_acc_psp_sva_1[11:0];
  assign return_add_generic_AC_RND_CONV_false_6_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_6_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_6_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_6_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_17_if_5_return_add_generic_AC_RND_CONV_false_17_if_5_and_tmp
      = (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1==10'b1111111111)
      & operator_6_false_17_acc_itm_0 & (~ BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0)
      & (z_out_89[53]);
  assign return_mult_generic_AC_RND_CONV_false_if_or_3_cse = (~ (z_out_86[5])) |
      return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_if_not_nl = ~ return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_if_nand_1_cse = ~(MUX_v_4_2_2(4'b0000,
      (z_out_86[4:1]), return_mult_generic_AC_RND_CONV_false_if_not_nl));
  assign return_mult_generic_AC_RND_CONV_false_if_or_cse = (~ (z_out_86[0])) | return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1;
  assign return_add_generic_AC_RND_CONV_false_4_if_7_not_4 = ~(return_add_generic_AC_RND_CONV_false_17_if_5_return_add_generic_AC_RND_CONV_false_17_if_5_and_tmp
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign stage_d_mul_return_d_4_63_sva_2 = stage_PE_1_tmp_im_d_1_lpi_3_dfm_63_mx0
      ^ return_add_generic_AC_RND_CONV_false_18_mux_itm;
  assign return_mult_generic_AC_RND_CONV_false_if_1_aelse_return_mult_generic_AC_RND_CONV_false_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1) | (z_out_106[105]);
  assign return_mult_generic_AC_RND_CONV_false_if_if_not_1_nl = ~ (z_out_111[12]);
  assign return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      (z_out_111[11:0]), return_mult_generic_AC_RND_CONV_false_if_if_not_1_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_acc_tmp = return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1
      + 12'b000000000001;
  assign return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_acc_tmp = nl_return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_acc_tmp[11:0];
  assign return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_2_10_0_1 = MUX_v_11_2_2(11'b00000000000,
      return_mult_generic_AC_RND_CONV_false_else_2_else_else_mux_2, return_mult_generic_AC_RND_CONV_false_1_zero_m_return_mult_generic_AC_RND_CONV_false_1_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_1_r_zero_return_mult_generic_AC_RND_CONV_false_1_r_zero_nor_mdf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_1_e_incr_lpi_3_dfm_2 = ~((~(((z_out_106[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((z_out_106[51]) | return_mult_generic_AC_RND_CONV_false_if_1_aelse_return_mult_generic_AC_RND_CONV_false_if_1_aelse_or_2))
      | (z_out_106[105]))) | (operator_14_false_1_acc_psp_sva_12_10[2]));
  assign return_mult_generic_AC_RND_CONV_false_1_zero_m_return_mult_generic_AC_RND_CONV_false_1_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_1_r_zero_return_mult_generic_AC_RND_CONV_false_1_r_zero_nor_mdf_sva_1
      = ~(return_add_generic_AC_RND_CONV_false_17_mux_6_itm | return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign return_extract_17_return_extract_17_or_sva_1 = (return_add_generic_AC_RND_CONV_false_5_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1[51])
      & return_add_generic_AC_RND_CONV_false_5_if_7_not_4;
  assign return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_5_if_7_not_4);
  assign nor_186_cse = ~(MUX_v_10_2_2(z_out_91, 10'b1111111111, return_add_generic_AC_RND_CONV_false_18_if_5_return_add_generic_AC_RND_CONV_false_18_if_5_and_tmp));
  assign nor_183_nl = ~((~ return_add_generic_AC_RND_CONV_false_5_e_r_qelse_or_svs_mx0w0)
      | return_add_generic_AC_RND_CONV_false_18_if_5_return_add_generic_AC_RND_CONV_false_18_if_5_and_tmp);
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qr_10_1_lpi_3_dfm_1 = ~(MUX_v_10_2_2(nor_186_cse,
      10'b1111111111, nor_183_nl));
  assign return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_and_1_nl
      = (operator_32_false_1_acc_psp_sva_11_0[0]) & return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_5_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_and_1_nl,
      operator_6_false_21_acc_itm_0, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_5_mux_13_nl
      & (~ return_add_generic_AC_RND_CONV_false_5_e_r_qelse_or_svs_mx0w0)) | return_add_generic_AC_RND_CONV_false_18_if_5_return_add_generic_AC_RND_CONV_false_18_if_5_and_tmp;
  assign return_extract_17_return_extract_17_nor_tmp = ~((return_add_generic_AC_RND_CONV_false_5_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1);
  assign operator_11_true_17_operator_11_true_17_and_tmp = (return_add_generic_AC_RND_CONV_false_5_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1;
  assign return_extract_49_m_zero_return_extract_49_m_zero_nor_tmp = ~(return_add_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_1
      | (return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_mult_generic_AC_RND_CONV_false_3_lor_lpi_3_dfm_1 = operator_11_true_return_22_sva
      | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva | return_mult_generic_AC_RND_CONV_false_1_exp_ovf_return_mult_generic_AC_RND_CONV_false_1_exp_ovf_or_tmp
      | return_add_generic_AC_RND_CONV_false_11_do_sub_sva;
  assign return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_2_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva, operator_14_false_1_acc_psp_sva_12_10[2]);
  assign return_mult_generic_AC_RND_CONV_false_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_2_nl
      & (~ (z_out_106[105]));
  assign return_add_generic_AC_RND_CONV_false_18_if_5_return_add_generic_AC_RND_CONV_false_18_if_5_and_tmp
      = (drf_qr_lval_19_smx_lpi_3_dfm[9:0]==10'b1111111111) & operator_6_false_21_acc_itm_0
      & (~ (drf_qr_lval_19_smx_lpi_3_dfm[10])) & (z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_5_if_7_not_4 = ~(return_add_generic_AC_RND_CONV_false_18_if_5_return_add_generic_AC_RND_CONV_false_18_if_5_and_tmp
      | return_add_generic_AC_RND_CONV_false_12_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_6_mux_31_nl = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_11,
      return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_not_3_nl = ~ return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1;
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(10'b0000000000,
      return_add_generic_AC_RND_CONV_false_6_mux_31_nl, return_add_generic_AC_RND_CONV_false_6_e_r_qelse_not_3_nl);
  assign return_mult_generic_AC_RND_CONV_false_2_if_nor_ovfl_sva_1 = ~((z_out_68[9:6]==4'b1111));
  assign return_extract_19_return_extract_19_nor_tmp = ~((return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1);
  assign return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp = ~(return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_19_return_extract_19_or_sva_1 = (return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1;
  assign and_600_nl = and_dcpl_224 & or_dcpl_320 & and_dcpl_64;
  assign return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_r_nan_or_mx6w0,
      (return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1[51]),
      and_600_nl);
  assign return_add_generic_AC_RND_CONV_false_6_if_7_return_add_generic_AC_RND_CONV_false_6_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_6_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_6_if_7_return_add_generic_AC_RND_CONV_false_6_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_6_exception_sva_1);
  assign and_293_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign or_389_nl = or_dcpl_324 | and_293_cse | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva;
  assign return_add_generic_AC_RND_CONV_false_19_e_r_qelse_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs, or_389_nl);
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_6_mux_36
      & (~ return_add_generic_AC_RND_CONV_false_19_e_r_qelse_mux_nl)) | return_add_generic_AC_RND_CONV_false_6_exception_sva_1;
  assign operator_11_true_19_operator_11_true_19_and_tmp = (return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1;
  assign return_mult_generic_AC_RND_CONV_false_4_lor_lpi_3_dfm_1 = return_add_generic_AC_RND_CONV_false_10_op2_inf_sva
      | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva | return_mult_generic_AC_RND_CONV_false_1_exp_ovf_return_mult_generic_AC_RND_CONV_false_1_exp_ovf_or_tmp
      | return_add_generic_AC_RND_CONV_false_11_do_sub_sva;
  assign return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_3_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva, operator_14_false_1_acc_psp_sva_12_10[2]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_3_nl
      & (~ (z_out_106[105]));
  assign return_add_generic_AC_RND_CONV_false_6_if_5_or_nl = and_293_cse | return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm;
  assign return_add_generic_AC_RND_CONV_false_6_mux_16_nl = MUX_s_1_2_2(and_293_cse,
      return_add_generic_AC_RND_CONV_false_6_if_5_or_nl, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_6_exception_sva_1 = operator_11_true_return_22_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_6_mux_16_nl;
  assign return_mult_generic_AC_RND_CONV_false_2_if_or_3_cse = (~ (z_out_68[5]))
      | return_mult_generic_AC_RND_CONV_false_2_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_2_if_not_nl = ~ return_mult_generic_AC_RND_CONV_false_2_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_2_if_nand_1_cse = ~(MUX_v_4_2_2(4'b0000,
      (z_out_68[4:1]), return_mult_generic_AC_RND_CONV_false_2_if_not_nl));
  assign return_mult_generic_AC_RND_CONV_false_2_if_or_cse = (~ (z_out_68[0])) |
      return_mult_generic_AC_RND_CONV_false_2_if_nor_ovfl_sva_1;
  assign nl_return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp = ({1'b1 , BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0
      , BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1}) + conv_u2s_11_12(~
      return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp = nl_return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp[11:0];
  assign nl_return_add_generic_AC_RND_CONV_false_7_e_dif_qif_acc_1_nl = ({1'b1 ,
      return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1}) + conv_u2s_11_12({(~
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0) , (~ BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1)})
      + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_7_e_dif_qif_acc_1_nl = nl_return_add_generic_AC_RND_CONV_false_7_e_dif_qif_acc_1_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_7_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp,
      return_add_generic_AC_RND_CONV_false_7_e_dif_qif_acc_1_nl, return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp[11]);
  assign return_mult_generic_AC_RND_CONV_false_2_else_2_else_return_mult_generic_AC_RND_CONV_false_2_else_2_else_and_nl
      = MUX_v_11_2_2(11'b00000000000, return_mult_generic_AC_RND_CONV_false_else_2_else_else_mux_2,
      return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1 =
      MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_2_else_2_else_return_mult_generic_AC_RND_CONV_false_2_else_2_else_and_nl,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_5_lor_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[0])
      & return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1 = return_mult_generic_AC_RND_CONV_false_2_m_r_51_lpi_3_dfm_mx1
      | return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1 = (return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1[0])
      & return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1, and_dcpl_469);
  assign return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_51_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_7_mux_27_cse, and_dcpl_469);
  assign return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0, return_extract_21_mux_cse,
      and_dcpl_469);
  assign return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_0_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_469);
  assign and_602_nl = and_dcpl_479 & and_dcpl_534;
  assign return_mult_generic_AC_RND_CONV_false_2_m_r_51_lpi_3_dfm_mx1 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_do_sub_sva,
      (z_out_87[51]), and_602_nl);
  assign return_mult_generic_AC_RND_CONV_false_2_oelse_3_return_mult_generic_AC_RND_CONV_false_5_if_3_nor_nl
      = ~((~ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1) | return_mult_generic_AC_RND_CONV_false_5_lor_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (z_out_87[50:0]), return_mult_generic_AC_RND_CONV_false_2_oelse_3_return_mult_generic_AC_RND_CONV_false_5_if_3_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp = ({BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0
      , BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1}) == (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1);
  assign return_add_generic_AC_RND_CONV_false_7_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_108[54]))) | (return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (z_out_108[53]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_108[52]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_108[51]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_108[50]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_108[49]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_108[48]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_108[47]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_108[46]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_108[45]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_108[44]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_108[43]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_108[42]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_108[41]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_108[40]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_108[39]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_108[38]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_108[37]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_108[36]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_108[35]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_108[34]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_108[33]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_108[32]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_108[31]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_108[30]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_108[29]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_108[28]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_108[27]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_108[26]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_108[25]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_108[24]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_108[23]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_108[22]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_108[21]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_108[20]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_108[19]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_108[18]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_108[17]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_108[16]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_108[15]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_108[14]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_108[13]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_108[12]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_108[11]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_108[10]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_108[9]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_108[8]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_108[7]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_108[6]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_108[5]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_108[4]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_108[3]))) | (return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_108[2])));
  assign nl_return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp = ({1'b1 , drf_qr_lval_10_smx_lpi_3_dfm_rsp_0
      , drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0 , drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1})
      + conv_u2s_11_12(~ return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1)
      + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp = nl_return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp[11:0];
  assign nl_return_add_generic_AC_RND_CONV_false_8_e_dif_qif_acc_1_nl = ({1'b1 ,
      return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1}) + conv_u2s_11_12({(~
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_0) , (~ drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0)
      , (~ drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1)}) + 12'b000000000001;
  assign return_add_generic_AC_RND_CONV_false_8_e_dif_qif_acc_1_nl = nl_return_add_generic_AC_RND_CONV_false_8_e_dif_qif_acc_1_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_8_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp,
      return_add_generic_AC_RND_CONV_false_8_e_dif_qif_acc_1_nl, return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp[11]);
  assign return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[0])
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1,
      and_dcpl_467);
  assign return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_51_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm, return_add_generic_AC_RND_CONV_false_7_mux_27_cse,
      and_dcpl_467);
  assign return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_49_0,
      return_extract_21_mux_cse, and_dcpl_467);
  assign return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_0_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_467);
  assign return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp = ({drf_qr_lval_10_smx_lpi_3_dfm_rsp_0
      , drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0 , drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1})
      == (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1);
  assign return_add_generic_AC_RND_CONV_false_8_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_107[54]))) | (return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (z_out_107[53]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_107[52]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_107[51]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_107[50]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_107[49]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_107[48]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_107[47]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_107[46]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_107[45]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_107[44]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_107[43]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_107[42]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_107[41]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_107[40]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_107[39]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_107[38]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_107[37]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_107[36]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_107[35]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_107[34]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_107[33]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_107[32]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_107[31]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_107[30]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_107[29]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_107[28]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_107[27]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_107[26]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_107[25]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_107[24]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_107[23]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_107[22]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_107[21]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_107[20]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_107[19]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_107[18]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_107[17]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_107[16]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_107[15]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_107[14]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_107[13]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_107[12]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_107[11]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_107[10]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_107[9]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_107[8]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_107[7]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_107[6]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_107[5]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_107[4]))) | ((return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_107[3]))) | (return_add_generic_AC_RND_CONV_false_8_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_107[2])));
  assign return_add_generic_AC_RND_CONV_false_8_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_8_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_8_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_8_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_7_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_7_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_7_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_7_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp
      = (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1!=11'b00000000000);
  assign return_mult_generic_AC_RND_CONV_false_5_lor_lpi_3_dfm_1 = return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | return_mult_generic_AC_RND_CONV_false_1_exp_ovf_return_mult_generic_AC_RND_CONV_false_1_exp_ovf_or_tmp
      | return_add_generic_AC_RND_CONV_false_11_do_sub_sva;
  assign return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva, operator_14_false_1_acc_psp_sva_12_10[2]);
  assign return_mult_generic_AC_RND_CONV_false_2_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_nl
      & (~ (z_out_106[105]));
  assign return_add_generic_AC_RND_CONV_false_7_mux_24_mx0_5_1 = MUX_v_5_2_2((drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0[4:0]),
      (return_add_generic_AC_RND_CONV_false_10_ls_sva[5:1]), return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_1_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_7_exception_sva_1);
  assign and_300_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_7_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign or_396_nl = and_300_cse | operator_11_true_return_1_sva | or_dcpl_285;
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_3_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs, or_396_nl);
  assign return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_1_mux_30
      & (~ return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_3_nl)) | return_add_generic_AC_RND_CONV_false_7_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_r_nan_or_cse,
      (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1[51]), and_2472_tmp);
  assign return_add_generic_AC_RND_CONV_false_7_if_7_return_add_generic_AC_RND_CONV_false_7_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_7_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1[50:0]),
      return_add_generic_AC_RND_CONV_false_7_if_7_return_add_generic_AC_RND_CONV_false_7_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_9_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_69,
      z_out_70, z_out_69[11]);
  assign return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1 = (stage_PE_1_x_re_d_sva[0])
      & return_add_generic_AC_RND_CONV_false_11_mux_itm;
  assign return_extract_25_return_extract_25_or_2_nl = (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_extract_25_return_extract_25_or_2_nl,
      return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1[50]), return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0 = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1[50:1]),
      (return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1[49:0]), return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1[0])
      & (~ return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[49:0]),
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_341);
  assign return_add_generic_AC_RND_CONV_false_9_e1_eq_e2_equal_tmp = (stage_PE_1_x_re_d_sva[62:52])
      == ({return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1});
  assign return_add_generic_AC_RND_CONV_false_9_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx2
      & (~ (z_out_110[54]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx2
      & (~ (z_out_110[53]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_110[52]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_110[51]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_110[50]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_110[49]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_110[48]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_110[47]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_110[46]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_110[45]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_110[44]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_110[43]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_110[42]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_110[41]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_110[40]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_110[39]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_110[38]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_110[37]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_110[36]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_110[35]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_110[34]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_110[33]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_110[32]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_110[31]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_110[30]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_110[29]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_110[28]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_110[27]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_110[26]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_110[25]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_110[24]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_110[23]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_110[22]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_110[21]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_110[20]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_110[19]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_110[18]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_110[17]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_110[16]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_110[15]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_110[14]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_110[13]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_110[12]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_110[11]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_110[10]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_110[9]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_110[8]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_110[7]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_110[6]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_110[5]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_110[4]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_110[3]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2
      & (~ (z_out_110[2])));
  assign return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_9_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_cse = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_9_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp
      = ~((return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_7_if_5_or_nl = and_300_cse | return_add_generic_AC_RND_CONV_false_if_5_return_add_generic_AC_RND_CONV_false_if_5_and_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_7_mux_18_nl = MUX_s_1_2_2(and_300_cse,
      return_add_generic_AC_RND_CONV_false_7_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_7_exception_sva_1 = return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0
      | return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0 | return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_mx2w0 | return_add_generic_AC_RND_CONV_false_7_mux_18_nl;
  assign return_add_generic_AC_RND_CONV_false_8_mux_20_mx0 = MUX_v_6_2_2((BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1[5:0]),
      return_add_generic_AC_RND_CONV_false_11_ls_sva, return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_8_e_r_qelse_not_5_nl = ~ return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1;
  assign return_add_generic_AC_RND_CONV_false_8_e_r_qelse_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(10'b0000000000,
      z_out_90, return_add_generic_AC_RND_CONV_false_8_e_r_qelse_not_5_nl);
  assign return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_8_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_8_exception_sva_1);
  assign and_307_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_8_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign or_404_nl = and_307_cse | operator_11_true_return_22_sva | or_dcpl_337;
  assign return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs, or_404_nl);
  assign return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_1_mux_30
      & (~ return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_nl)) | return_add_generic_AC_RND_CONV_false_8_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_8_r_nan_or_mx0w0 = return_add_generic_AC_RND_CONV_false_21_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | (return_add_generic_AC_RND_CONV_false_21_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva & return_add_generic_AC_RND_CONV_false_16_do_sub_sva);
  assign and_609_nl = and_dcpl_237 & and_dcpl_541;
  assign return_add_generic_AC_RND_CONV_false_8_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_r_nan_or_mx0w0,
      (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1[51]), and_609_nl);
  assign return_add_generic_AC_RND_CONV_false_8_if_7_return_add_generic_AC_RND_CONV_false_8_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_8_exception_sva_1 | return_add_generic_AC_RND_CONV_false_12_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1[50:0]),
      return_add_generic_AC_RND_CONV_false_8_if_7_return_add_generic_AC_RND_CONV_false_8_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_95,
      z_out_96, z_out_95[11]);
  assign return_extract_27_return_extract_27_or_2_nl = (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_extract_27_return_extract_27_or_2_nl,
      return_add_generic_AC_RND_CONV_false_8_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_10_op2_mu_1_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_m_r_51_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1[50]), return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_10_op2_mu_1_50_1_lpi_3_dfm_mx0 = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1[50:1]),
      (return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1[49:0]), return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1[0])
      & (~ return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(drf_qr_lval_13_smx_0_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx0,
      and_dcpl_446);
  assign return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_51_lpi_3_dfm_mx0 =
      MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[50]),
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_51_lpi_3_dfm_mx0, and_dcpl_446);
  assign return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49:0]),
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_446);
  assign return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1,
      and_dcpl_446);
  assign return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_equal_tmp = (stage_PE_1_tmp_re_d_sva[62:52])
      == ({return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1});
  assign return_add_generic_AC_RND_CONV_false_10_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_110[54]))) | (return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (z_out_110[53]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_110[52]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_110[51]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_110[50]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_110[49]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_110[48]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_110[47]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_110[46]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_110[45]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_110[44]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_110[43]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_110[42]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_110[41]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_110[40]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_110[39]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_110[38]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_110[37]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_110[36]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_110[35]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_110[34]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_110[33]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_110[32]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_110[31]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_110[30]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_110[29]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_110[28]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_110[27]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_110[26]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_110[25]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_110[24]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_110[23]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_110[22]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_110[21]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_110[20]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_110[19]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_110[18]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_110[17]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_110[16]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_110[15]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_110[14]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_110[13]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_110[12]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_110[11]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_110[10]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_110[9]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_110[8]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_110[7]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_110[6]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_110[5]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_110[4]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_110[3]))) | (return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_110[2])));
  assign return_add_generic_AC_RND_CONV_false_12_e_dif_qr_lpi_3_dfm_mx0_10_0 = MUX_v_11_2_2((z_out_95[10:0]),
      (z_out_96[10:0]), z_out_95[11]);
  assign return_add_generic_AC_RND_CONV_false_12_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_107[54]))) | (return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (z_out_107[53]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_107[52]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_107[51]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_107[50]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_107[49]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_107[48]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_107[47]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_107[46]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_107[45]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_107[44]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_107[43]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_107[42]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_107[41]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_107[40]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_107[39]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_107[38]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_107[37]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_107[36]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_107[35]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_107[34]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_107[33]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_107[32]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_107[31]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_107[30]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_107[29]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_107[28]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_107[27]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_107[26]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_107[25]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_107[24]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_107[23]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_107[22]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_107[21]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_107[20]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_107[19]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_107[18]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_107[17]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_107[16]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_107[15]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_107[14]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_107[13]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_107[12]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_107[11]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_107[10]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_107[9]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_107[8]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_107[7]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_107[6]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_107[5]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_107[4]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_107[3]))) | (return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_107[2])));
  assign return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_12_e_dif_qr_lpi_3_dfm_mx0_10_0[10:6]!=5'b00000)
      | ((z_out_96[11]) & (z_out_95[11]));
  assign return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_12_e_dif_qr_lpi_3_dfm_mx0_10_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_10_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_10_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_10_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_10_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp
      = ~((return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_21_op1_nan_sva_1 = operator_11_true_return_22_sva
      & (~ return_extract_22_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_21_op1_inf_sva_1 = operator_11_true_return_22_sva
      & return_extract_22_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_8_if_5_or_nl = and_307_cse | return_add_generic_AC_RND_CONV_false_if_5_return_add_generic_AC_RND_CONV_false_if_5_and_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_8_mux_14_nl = MUX_s_1_2_2(and_307_cse,
      return_add_generic_AC_RND_CONV_false_8_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_8_exception_sva_1 = return_add_generic_AC_RND_CONV_false_21_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_21_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_8_mux_14_nl;
  assign return_add_generic_AC_RND_CONV_false_9_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      z_out_103, return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva);
  assign return_add_generic_AC_RND_CONV_false_11_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm
      & (~ (z_out_109[54]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm
      & (~ (z_out_109[53]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[49])
      & (~ (z_out_109[52]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[48])
      & (~ (z_out_109[51]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[47])
      & (~ (z_out_109[50]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[46])
      & (~ (z_out_109[49]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[45])
      & (~ (z_out_109[48]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[44])
      & (~ (z_out_109[47]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[43])
      & (~ (z_out_109[46]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[42])
      & (~ (z_out_109[45]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[41])
      & (~ (z_out_109[44]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[40])
      & (~ (z_out_109[43]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[39])
      & (~ (z_out_109[42]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[38])
      & (~ (z_out_109[41]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[37])
      & (~ (z_out_109[40]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[36])
      & (~ (z_out_109[39]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[35])
      & (~ (z_out_109[38]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[34])
      & (~ (z_out_109[37]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[33])
      & (~ (z_out_109[36]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[32])
      & (~ (z_out_109[35]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[31])
      & (~ (z_out_109[34]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[30])
      & (~ (z_out_109[33]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[29])
      & (~ (z_out_109[32]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[28])
      & (~ (z_out_109[31]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[27])
      & (~ (z_out_109[30]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[26])
      & (~ (z_out_109[29]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[25])
      & (~ (z_out_109[28]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[24])
      & (~ (z_out_109[27]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[23])
      & (~ (z_out_109[26]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[22])
      & (~ (z_out_109[25]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[21])
      & (~ (z_out_109[24]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[20])
      & (~ (z_out_109[23]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[19])
      & (~ (z_out_109[22]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[18])
      & (~ (z_out_109[21]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[17])
      & (~ (z_out_109[20]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[16])
      & (~ (z_out_109[19]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[15])
      & (~ (z_out_109[18]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[14])
      & (~ (z_out_109[17]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[13])
      & (~ (z_out_109[16]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[12])
      & (~ (z_out_109[15]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[11])
      & (~ (z_out_109[14]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[10])
      & (~ (z_out_109[13]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[9])
      & (~ (z_out_109[12]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[8])
      & (~ (z_out_109[11]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[7])
      & (~ (z_out_109[10]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[6])
      & (~ (z_out_109[9]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[5])
      & (~ (z_out_109[8]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[4])
      & (~ (z_out_109[7]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[3])
      & (~ (z_out_109[6]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[2])
      & (~ (z_out_109[5]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[1])
      & (~ (z_out_109[4]))) | ((return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0[0])
      & (~ (z_out_109[3]))) | return_add_generic_AC_RND_CONV_false_4_sticky_bit_and_158;
  assign return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp
      = (return_add_generic_AC_RND_CONV_false_9_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_2_cse
      & (return_add_generic_AC_RND_CONV_false_9_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_9_if_5_or_nl = and_340_cse | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_9_mux_17_nl = MUX_s_1_2_2(and_340_cse,
      return_add_generic_AC_RND_CONV_false_9_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_9_exception_sva_1 = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0 | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0 | return_add_generic_AC_RND_CONV_false_9_mux_17_nl;
  assign return_add_generic_AC_RND_CONV_false_9_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_9_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_10_if_5_or_nl = and_348_cse | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_10_mux_17_nl = MUX_s_1_2_2(and_348_cse,
      return_add_generic_AC_RND_CONV_false_10_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_10_exception_sva_1 = operator_11_true_return_22_sva
      | return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0 | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_mx2w0 | return_add_generic_AC_RND_CONV_false_10_mux_17_nl;
  assign return_add_generic_AC_RND_CONV_false_10_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_10_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_11_if_5_or_nl = and_356_cse | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_11_mux_10_nl = MUX_s_1_2_2(and_356_cse,
      return_add_generic_AC_RND_CONV_false_11_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_11_exception_sva_1 = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      | operator_11_true_return_26_sva | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_unequal_tmp | return_add_generic_AC_RND_CONV_false_11_mux_10_nl;
  assign return_add_generic_AC_RND_CONV_false_11_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_11_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_12_if_5_or_nl = and_362_cse | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_12_mux_10_nl = MUX_s_1_2_2(and_362_cse,
      return_add_generic_AC_RND_CONV_false_12_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_12_exception_sva_1 = operator_11_true_return_22_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_12_mux_10_nl;
  assign return_add_generic_AC_RND_CONV_false_12_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_12_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_12_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_14_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_95,
      z_out_70, z_out_71_11);
  assign return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1 = (in_f_d_rsci_q_d[0])
      & return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_1, and_dcpl_452);
  assign return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0
      = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm,
      return_extract_33_mux_3_cse, and_dcpl_452);
  assign return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1,
      and_dcpl_452);
  assign return_add_generic_AC_RND_CONV_false_14_e1_eq_e2_equal_tmp = (stage_PE_1_tmp_re_d_sva[62:52])
      == (in_f_d_rsci_q_d[62:52]);
  assign return_add_generic_AC_RND_CONV_false_14_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_109[54]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_109[53]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_109[52]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_109[51]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_109[50]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_109[49]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_109[48]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_109[47]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_109[46]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_109[45]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_109[44]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_109[43]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_109[42]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_109[41]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_109[40]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_109[39]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_109[38]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_109[37]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_109[36]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_109[35]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_109[34]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_109[33]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_109[32]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_109[31]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_109[30]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_109[29]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_109[28]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_109[27]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_109[26]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_109[25]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_109[24]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_109[23]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_109[22]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_109[21]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_109[20]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_109[19]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_109[18]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_109[17]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_109[16]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_109[15]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_109[14]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_109[13]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_109[12]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_109[11]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_109[10]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_109[9]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_109[8]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_109[7]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_109[6]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_109[5]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_109[4]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_109[3]))) | (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_109[2])));
  assign return_add_generic_AC_RND_CONV_false_16_e_dif_qr_lpi_3_dfm_mx0_10_0 = MUX_v_11_2_2((z_out_95[10:0]),
      (z_out_70[10:0]), z_out_95[11]);
  assign return_add_generic_AC_RND_CONV_false_16_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_107[54]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_107[53]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_107[52]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_107[51]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_107[50]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_107[49]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_107[48]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_107[47]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_107[46]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_107[45]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_107[44]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_107[43]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_107[42]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_107[41]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_107[40]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_107[39]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_107[38]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_107[37]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_107[36]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_107[35]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_107[34]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_107[33]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_107[32]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_107[31]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_107[30]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_107[29]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_107[28]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_107[27]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_107[26]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_107[25]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_107[24]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_107[23]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_107[22]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_107[21]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_107[20]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_107[19]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_107[18]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_107[17]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_107[16]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_107[15]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_107[14]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_107[13]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_107[12]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_107[11]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_107[10]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_107[9]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_107[8]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_107[7]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_107[6]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_107[5]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_107[4]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_107[3]))) | (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_107[2])));
  assign return_add_generic_AC_RND_CONV_false_13_e_dif1_return_add_generic_AC_RND_CONV_false_13_e_dif1_and_cse
      = (z_out_70[11]) & (z_out_95[11]);
  assign return_add_generic_AC_RND_CONV_false_16_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_16_e_dif_qr_lpi_3_dfm_mx0_10_0[10:6]!=5'b00000)
      | return_add_generic_AC_RND_CONV_false_13_e_dif1_return_add_generic_AC_RND_CONV_false_13_e_dif1_and_cse;
  assign return_add_generic_AC_RND_CONV_false_16_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_16_e_dif_qr_lpi_3_dfm_mx0_10_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_16_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_14_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_14_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_14_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_14_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_14_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_14_if_5_or_nl = and_311_cse | return_add_generic_AC_RND_CONV_false_if_5_return_add_generic_AC_RND_CONV_false_if_5_and_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_14_mux_16_nl = MUX_s_1_2_2(and_311_cse,
      return_add_generic_AC_RND_CONV_false_14_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_14_exception_sva_1 = return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0
      | return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0 | return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_mx2w0 | return_add_generic_AC_RND_CONV_false_14_mux_16_nl;
  assign return_add_generic_AC_RND_CONV_false_13_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_70,
      z_out_95, z_out_69[11]);
  assign return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_1,
      drf_qr_lval_13_smx_0_lpi_3_dfm, and_dcpl_468);
  assign return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0
      = MUX_v_51_2_2(return_extract_33_mux_3_cse, return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm,
      and_dcpl_468);
  assign return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_13_op2_mu_0_lpi_3_dfm_1,
      and_dcpl_468);
  assign return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp = (in_f_d_rsci_q_d[62:52])
      == (stage_PE_1_tmp_re_d_sva[62:52]);
  assign return_add_generic_AC_RND_CONV_false_13_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_109[54]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_109[53]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_109[52]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_109[51]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_109[50]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_109[49]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_109[48]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_109[47]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_109[46]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_109[45]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_109[44]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_109[43]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_109[42]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_109[41]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_109[40]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_109[39]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_109[38]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_109[37]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_109[36]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_109[35]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_109[34]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_109[33]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_109[32]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_109[31]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_109[30]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_109[29]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_109[28]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_109[27]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_109[26]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_109[25]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_109[24]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_109[23]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_109[22]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_109[21]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_109[20]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_109[19]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_109[18]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_109[17]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_109[16]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_109[15]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_109[14]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_109[13]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_109[12]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_109[11]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_109[10]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_109[9]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_109[8]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_109[7]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_109[6]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_109[5]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_109[4]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_109[3]))) | (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_109[2])));
  assign return_add_generic_AC_RND_CONV_false_15_e_dif_qr_lpi_3_dfm_mx0_10_0 = MUX_v_11_2_2((z_out_70[10:0]),
      (z_out_95[10:0]), z_out_70[11]);
  assign return_add_generic_AC_RND_CONV_false_15_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_107[54]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_107[53]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_107[52]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_107[51]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_107[50]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_107[49]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_107[48]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_107[47]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_107[46]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_107[45]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_107[44]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_107[43]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_107[42]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_107[41]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_107[40]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_107[39]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_107[38]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_107[37]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_107[36]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_107[35]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_107[34]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_107[33]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_107[32]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_107[31]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_107[30]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_107[29]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_107[28]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_107[27]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_107[26]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_107[25]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_107[24]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_107[23]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_107[22]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_107[21]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_107[20]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_107[19]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_107[18]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_107[17]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_107[16]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_107[15]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_107[14]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_107[13]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_107[12]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_107[11]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_107[10]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_107[9]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_107[8]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_107[7]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_107[6]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_107[5]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_107[4]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_107[3]))) | (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_107[2])));
  assign return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_15_e_dif_qr_lpi_3_dfm_mx0_10_0[10:6]!=5'b00000)
      | return_add_generic_AC_RND_CONV_false_13_e_dif1_return_add_generic_AC_RND_CONV_false_13_e_dif1_and_cse;
  assign return_add_generic_AC_RND_CONV_false_15_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_15_e_dif_qr_lpi_3_dfm_mx0_10_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_13_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_13_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_13_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_13_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_13_e_dif_sat_or_1_nl);
  assign nl_operator_32_false_3_acc_psp_sva_1 = conv_s2s_17_18(stage_u_add_acc_1_itm_1)
      + conv_s2s_17_18(z_out_111);
  assign operator_32_false_3_acc_psp_sva_1 = nl_operator_32_false_3_acc_psp_sva_1[17:0];
  assign nl_return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl = ({1'b1
      , (in_f_d_rsci_q_d[51:0])}) + conv_u2u_52_53(~ (stage_PE_1_tmp_re_d_sva[51:0]))
      + 53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl[52:0];
  assign return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_itm_52 = readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl);
  assign return_add_generic_AC_RND_CONV_false_13_if_5_or_nl = and_317_cse | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_13_mux_16_nl = MUX_s_1_2_2(and_317_cse,
      return_add_generic_AC_RND_CONV_false_13_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_13_exception_sva_1 = return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0
      | return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0 | return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_mx2w0 | return_add_generic_AC_RND_CONV_false_13_mux_16_nl;
  assign return_add_generic_AC_RND_CONV_false_13_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_13_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_15_exp_plus_1_12_1_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      z_out_114, return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_15_exp_plus_1_0_lpi_3_dfm_1 = (z_out_94[0])
      | (~ return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_15_if_5_return_add_generic_AC_RND_CONV_false_15_if_5_and_tmp
      = (return_add_generic_AC_RND_CONV_false_15_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_15_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_15_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_15_if_5_or_nl = return_add_generic_AC_RND_CONV_false_15_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_15_if_5_return_add_generic_AC_RND_CONV_false_15_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_15_mux_14_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_15_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_15_if_5_or_nl, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_15_exception_sva_1 = operator_11_true_return_22_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_15_mux_14_nl;
  assign return_add_generic_AC_RND_CONV_false_15_r_inf_lpi_3_dfm_2 = or_1997_cse
      & return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_15_mux_4_itm_5_1 = MUX_v_5_2_2((drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0[4:0]),
      (return_add_generic_AC_RND_CONV_false_10_ls_sva[5:1]), return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_16_exp_plus_1_0_lpi_3_dfm_1 = (operator_33_true_36_acc_psp_1_sva[0])
      | (~ return_add_generic_AC_RND_CONV_false_16_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_16_if_5_return_add_generic_AC_RND_CONV_false_16_if_5_and_tmp
      = (return_add_generic_AC_RND_CONV_false_3_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_16_exp_plus_1_0_lpi_3_dfm_1 & return_add_generic_AC_RND_CONV_false_3_if_5_nor_cse;
  assign return_add_generic_AC_RND_CONV_false_16_if_5_or_nl = return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_16_if_5_return_add_generic_AC_RND_CONV_false_16_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_16_mux_14_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_16_if_5_or_nl, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_16_exception_sva_1 = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      | operator_11_true_return_26_sva | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_unequal_tmp | return_add_generic_AC_RND_CONV_false_16_mux_14_nl;
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50 = MUX_s_1_2_2((in_f_d_rsci_q_d[50]),
      (return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[50]),
      inverse_lpi_1_dfm_1);
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_63_mx0 = MUX_s_1_2_2((in_f_d_rsci_q_d[63]),
      return_add_generic_AC_RND_CONV_false_16_mux_itm, inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0_mx0 =
      MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx2[50:1]),
      (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx2[49:0]),
      return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_19_op2_mu_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx2[0])
      & (~ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp);
  assign drf_qr_lval_22_smx_lpi_3_dfm_mx0_10 = MUX_s_1_2_2((drf_qr_lval_10_smx_lpi_3_dfm_mx7_10_1[9]),
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_0, and_dcpl_543);
  assign drf_qr_lval_22_smx_lpi_3_dfm_mx0_9_1 = MUX_v_9_2_2((drf_qr_lval_10_smx_lpi_3_dfm_mx7_10_1[8:0]),
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0, and_dcpl_543);
  assign drf_qr_lval_22_smx_lpi_3_dfm_mx0_0 = MUX_s_1_2_2(drf_qr_lval_10_smx_lpi_3_dfm_mx7_0,
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1, and_dcpl_543);
  assign return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(drf_qr_lval_13_smx_0_lpi_3_dfm, drf_qr_lval_13_smx_0_lpi_3_dfm_mx3,
      and_dcpl_543);
  assign return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_50_mx0
      = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm_mx3,
      and_dcpl_543);
  assign return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0
      = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0, return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0_mx0,
      and_dcpl_543);
  assign return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_19_op2_mu_0_lpi_3_dfm_1,
      and_dcpl_543);
  assign return_add_generic_AC_RND_CONV_false_19_e1_eq_e2_equal_tmp = ({drf_qr_lval_10_smx_lpi_3_dfm_rsp_0
      , drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0 , drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1})
      == ({drf_qr_lval_10_smx_lpi_3_dfm_mx7_10_1 , drf_qr_lval_10_smx_lpi_3_dfm_mx7_0});
  assign return_add_generic_AC_RND_CONV_false_19_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_19_op1_smaller_oelse_and_cse
      = z_out_57_52 & return_add_generic_AC_RND_CONV_false_19_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_19_op1_smaller_lor_lpi_3_dfm_2 = return_add_generic_AC_RND_CONV_false_19_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_19_op1_smaller_oelse_and_cse
      | (z_out_69[11]);
  assign return_add_generic_AC_RND_CONV_false_19_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_109[54]))) | (return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_50_mx0
      & (~ (z_out_109[53]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[49])
      & (~ (z_out_109[52]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[48])
      & (~ (z_out_109[51]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[47])
      & (~ (z_out_109[50]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[46])
      & (~ (z_out_109[49]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[45])
      & (~ (z_out_109[48]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[44])
      & (~ (z_out_109[47]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[43])
      & (~ (z_out_109[46]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[42])
      & (~ (z_out_109[45]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[41])
      & (~ (z_out_109[44]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[40])
      & (~ (z_out_109[43]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[39])
      & (~ (z_out_109[42]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[38])
      & (~ (z_out_109[41]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[37])
      & (~ (z_out_109[40]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[36])
      & (~ (z_out_109[39]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[35])
      & (~ (z_out_109[38]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[34])
      & (~ (z_out_109[37]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[33])
      & (~ (z_out_109[36]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[32])
      & (~ (z_out_109[35]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[31])
      & (~ (z_out_109[34]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[30])
      & (~ (z_out_109[33]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[29])
      & (~ (z_out_109[32]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[28])
      & (~ (z_out_109[31]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[27])
      & (~ (z_out_109[30]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[26])
      & (~ (z_out_109[29]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[25])
      & (~ (z_out_109[28]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[24])
      & (~ (z_out_109[27]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[23])
      & (~ (z_out_109[26]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[22])
      & (~ (z_out_109[25]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[21])
      & (~ (z_out_109[24]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[20])
      & (~ (z_out_109[23]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[19])
      & (~ (z_out_109[22]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[18])
      & (~ (z_out_109[21]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[17])
      & (~ (z_out_109[20]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[16])
      & (~ (z_out_109[19]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[15])
      & (~ (z_out_109[18]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[14])
      & (~ (z_out_109[17]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[13])
      & (~ (z_out_109[16]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[12])
      & (~ (z_out_109[15]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[11])
      & (~ (z_out_109[14]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[10])
      & (~ (z_out_109[13]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[9])
      & (~ (z_out_109[12]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[8])
      & (~ (z_out_109[11]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[7])
      & (~ (z_out_109[10]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[6])
      & (~ (z_out_109[9]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[5])
      & (~ (z_out_109[8]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[4])
      & (~ (z_out_109[7]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[3])
      & (~ (z_out_109[6]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[2])
      & (~ (z_out_109[5]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[1])
      & (~ (z_out_109[4]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[0])
      & (~ (z_out_109[3]))) | (return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_109[2])));
  assign return_extract_47_return_extract_47_or_sva_1 = (return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm_1;
  assign nor_187_nl = ~((~ return_add_generic_AC_RND_CONV_false_17_e_r_qelse_or_svs_mx0w0)
      | return_add_generic_AC_RND_CONV_false_17_if_5_return_add_generic_AC_RND_CONV_false_17_if_5_and_tmp);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_1 = ~(MUX_v_10_2_2(nor_182_cse,
      10'b1111111111, nor_187_nl));
  assign return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_and_3_nl
      = (operator_32_false_1_acc_psp_sva_11_0[0]) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_17_mux_19_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_and_3_nl,
      operator_6_false_17_acc_itm_0, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_17_mux_19_nl
      & (~ return_add_generic_AC_RND_CONV_false_17_e_r_qelse_or_svs_mx0w0)) | return_add_generic_AC_RND_CONV_false_17_if_5_return_add_generic_AC_RND_CONV_false_17_if_5_and_tmp;
  assign return_extract_47_return_extract_47_nor_tmp = ~((return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm_1);
  assign operator_11_true_47_operator_11_true_47_and_tmp = (return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm_1;
  assign nl_operator_6_false_42_acc_psp_sva_1 = conv_u2s_11_12({drf_qr_lval_22_smx_lpi_3_dfm_mx0_10
      , drf_qr_lval_22_smx_lpi_3_dfm_mx0_9_1 , drf_qr_lval_22_smx_lpi_3_dfm_mx0_0})
      + conv_s2s_7_12({1'b1 , (~ leading_sign_57_0_1_0_19_out_3)}) + 12'b000000000001;
  assign operator_6_false_42_acc_psp_sva_1 = nl_operator_6_false_42_acc_psp_sva_1[11:0];
  assign return_extract_49_return_extract_49_or_sva_1 = (return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_18_e_r_qr_0_lpi_3_dfm_1;
  assign nor_191_nl = ~((~ return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_svs_mx0w0)
      | return_add_generic_AC_RND_CONV_false_18_if_5_return_add_generic_AC_RND_CONV_false_18_if_5_and_tmp);
  assign return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1 = ~(MUX_v_10_2_2(nor_186_cse,
      10'b1111111111, nor_191_nl));
  assign return_add_generic_AC_RND_CONV_false_18_return_add_generic_AC_RND_CONV_false_18_and_1_nl
      = (operator_33_true_36_acc_psp_1_sva[0]) & return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_18_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_18_return_add_generic_AC_RND_CONV_false_18_and_1_nl,
      operator_6_false_21_acc_itm_0, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_18_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_18_mux_13_nl
      & (~ return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_svs_mx0w0)) | return_add_generic_AC_RND_CONV_false_18_if_5_return_add_generic_AC_RND_CONV_false_18_if_5_and_tmp;
  assign return_extract_49_return_extract_49_nor_tmp = ~((return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_18_e_r_qr_0_lpi_3_dfm_1);
  assign operator_11_true_49_operator_11_true_49_and_tmp = (return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_18_e_r_qr_0_lpi_3_dfm_1;
  assign return_mult_generic_AC_RND_CONV_false_1_exp_ovf_return_mult_generic_AC_RND_CONV_false_1_exp_ovf_or_tmp
      = return_mult_generic_AC_RND_CONV_false_1_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_1_exp_ovf_oif_aelse_and_1_tmp
      | (return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_acc_tmp[11]);
  assign return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_5_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva, operator_14_false_1_acc_psp_sva_12_10[2]);
  assign return_mult_generic_AC_RND_CONV_false_3_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_5_nl
      & (~ (z_out_106[105]));
  assign return_extract_51_return_extract_51_nor_tmp = ~((return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1);
  assign return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp = ~(return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_51_return_extract_51_or_sva_1 = (return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1;
  assign and_612_nl = and_dcpl_224 & or_dcpl_371 & and_dcpl_64;
  assign return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_r_nan_or_mx6w0,
      (return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1[51]),
      and_612_nl);
  assign return_add_generic_AC_RND_CONV_false_19_if_7_return_add_generic_AC_RND_CONV_false_19_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_19_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_add_generic_AC_RND_CONV_false_19_if_7_return_add_generic_AC_RND_CONV_false_19_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_19_exception_sva_1);
  assign and_324_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign or_438_nl = or_dcpl_324 | and_324_cse | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva;
  assign return_add_generic_AC_RND_CONV_false_19_e_r_qelse_mux_2_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs, or_438_nl);
  assign return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_6_mux_36
      & (~ return_add_generic_AC_RND_CONV_false_19_e_r_qelse_mux_2_nl)) | return_add_generic_AC_RND_CONV_false_19_exception_sva_1;
  assign operator_11_true_51_operator_11_true_51_and_tmp = (return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1;
  assign return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_6_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva, operator_14_false_1_acc_psp_sva_12_10[2]);
  assign return_mult_generic_AC_RND_CONV_false_4_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_6_nl
      & (~ (z_out_106[105]));
  assign return_add_generic_AC_RND_CONV_false_19_if_5_or_nl = and_324_cse | return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm;
  assign return_add_generic_AC_RND_CONV_false_19_mux_16_nl = MUX_s_1_2_2(and_324_cse,
      return_add_generic_AC_RND_CONV_false_19_if_5_or_nl, z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_19_exception_sva_1 = operator_11_true_return_22_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_19_mux_16_nl;
  assign return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[0])
      & return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1 = return_mult_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_mx1
      | return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(drf_qr_lval_13_smx_0_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1,
      and_dcpl_467);
  assign return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_51_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_20_mux_27_cse, and_dcpl_467);
  assign return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0, return_extract_21_mux_cse,
      and_dcpl_467);
  assign return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_467);
  assign and_614_nl = and_dcpl_474 & (~ (return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_acc_tmp[11]))
      & and_dcpl_534;
  assign return_mult_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_mx1 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_do_sub_sva,
      (z_out_87[51]), and_614_nl);
  assign return_add_generic_AC_RND_CONV_false_20_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_108[54]))) | (return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (z_out_108[53]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_108[52]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_108[51]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_108[50]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_108[49]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_108[48]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_108[47]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_108[46]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_108[45]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_108[44]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_108[43]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_108[42]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_108[41]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_108[40]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_108[39]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_108[38]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_108[37]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_108[36]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_108[35]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_108[34]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_108[33]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_108[32]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_108[31]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_108[30]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_108[29]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_108[28]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_108[27]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_108[26]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_108[25]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_108[24]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_108[23]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_108[22]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_108[21]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_108[20]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_108[19]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_108[18]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_108[17]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_108[16]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_108[15]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_108[14]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_108[13]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_108[12]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_108[11]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_108[10]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_108[9]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_108[8]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_108[7]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_108[6]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_108[5]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_108[4]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_108[3]))) | (return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_108[2])));
  assign return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm[0])
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm, return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1,
      and_dcpl_469);
  assign return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_51_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm, return_add_generic_AC_RND_CONV_false_20_mux_27_cse,
      and_dcpl_469);
  assign return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_49_0,
      return_extract_21_mux_cse, and_dcpl_469);
  assign return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_469);
  assign return_add_generic_AC_RND_CONV_false_21_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_107[54]))) | (return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (z_out_107[53]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_107[52]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_107[51]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_107[50]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_107[49]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_107[48]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_107[47]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_107[46]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_107[45]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_107[44]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_107[43]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_107[42]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_107[41]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_107[40]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_107[39]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_107[38]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_107[37]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_107[36]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_107[35]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_107[34]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_107[33]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_107[32]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_107[31]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_107[30]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_107[29]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_107[28]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_107[27]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_107[26]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_107[25]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_107[24]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_107[23]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_107[22]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_107[21]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_107[20]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_107[19]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_107[18]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_107[17]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_107[16]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_107[15]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_107[14]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_107[13]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_107[12]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_107[11]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_107[10]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_107[9]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_107[8]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_107[7]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_107[6]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_107[5]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_107[4]))) | ((return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_107[3]))) | (return_add_generic_AC_RND_CONV_false_21_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_107[2])));
  assign return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_4_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva, operator_14_false_1_acc_psp_sva_12_10[2]);
  assign return_mult_generic_AC_RND_CONV_false_5_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_4_nl
      & (~ (z_out_106[105]));
  assign return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_1_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_20_exception_sva_1);
  assign and_328_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_20_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign or_443_nl = and_328_cse | operator_11_true_return_1_sva | or_dcpl_285;
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_6_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs, or_443_nl);
  assign return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_1_mux_30
      & (~ return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_6_nl)) | return_add_generic_AC_RND_CONV_false_20_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_20_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1
      & return_mult_generic_AC_RND_CONV_false_1_op1_zero_sva_1 & return_add_generic_AC_RND_CONV_false_20_do_sub_sva);
  assign and_615_nl = and_dcpl_259 & and_dcpl_503;
  assign return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_20_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1[51]), and_615_nl);
  assign return_add_generic_AC_RND_CONV_false_20_if_7_return_add_generic_AC_RND_CONV_false_20_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_20_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1[50:0]),
      return_add_generic_AC_RND_CONV_false_20_if_7_return_add_generic_AC_RND_CONV_false_20_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_96,
      (z_out_98[11:0]), z_out_96[11]);
  assign return_extract_57_return_extract_57_or_2_nl = (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_extract_57_return_extract_57_or_2_nl,
      return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1[50]), return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0 = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1[50:1]),
      (return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1[49:0]), return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1[0])
      & (~ return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0, and_dcpl_340);
  assign return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49:0]),
      return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_340);
  assign return_add_generic_AC_RND_CONV_false_22_e1_eq_e2_equal_tmp = (stage_PE_1_x_re_d_sva[62:52])
      == ({return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1});
  assign return_add_generic_AC_RND_CONV_false_22_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_110[54]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx4
      & (~ (z_out_110[53]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_110[52]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_110[51]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_110[50]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_110[49]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_110[48]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_110[47]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_110[46]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_110[45]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_110[44]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_110[43]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_110[42]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_110[41]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_110[40]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_110[39]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_110[38]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_110[37]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_110[36]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_110[35]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_110[34]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_110[33]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_110[32]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_110[31]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_110[30]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_110[29]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_110[28]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_110[27]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_110[26]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_110[25]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_110[24]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_110[23]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_110[22]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_110[21]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_110[20]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_110[19]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_110[18]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_110[17]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_110[16]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_110[15]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_110[14]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_110[13]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_110[12]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_110[11]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_110[10]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_110[9]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_110[8]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_110[7]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_110[6]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_110[5]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_110[4]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_110[3]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx3
      & (~ (z_out_110[2])));
  assign return_add_generic_AC_RND_CONV_false_24_e_dif_qr_lpi_3_dfm_mx0_10_0 = MUX_v_11_2_2((z_out_96[10:0]),
      (z_out_98[10:0]), z_out_96[11]);
  assign return_add_generic_AC_RND_CONV_false_22_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_22_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_22_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_22_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp
      = ~((return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_20_if_5_or_nl = and_328_cse | return_add_generic_AC_RND_CONV_false_if_5_return_add_generic_AC_RND_CONV_false_if_5_and_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_20_mux_18_nl = MUX_s_1_2_2(and_328_cse,
      return_add_generic_AC_RND_CONV_false_20_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_20_exception_sva_1 = return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1
      | return_mult_generic_AC_RND_CONV_false_1_op1_zero_sva_1 | return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_20_mux_18_nl;
  assign return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_8_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_21_exception_sva_1);
  assign and_332_cse = ((operator_33_true_12_acc_psp_sva[11]) | (~ return_add_generic_AC_RND_CONV_false_21_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign or_447_nl = and_332_cse | operator_11_true_return_22_sva | or_dcpl_337;
  assign return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs, or_447_nl);
  assign return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_1_mux_30
      & (~ return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_1_nl)) | return_add_generic_AC_RND_CONV_false_21_exception_sva_1;
  assign and_616_nl = and_dcpl_263 & and_dcpl_541;
  assign return_add_generic_AC_RND_CONV_false_21_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_r_nan_or_mx0w0,
      (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1[51]), and_616_nl);
  assign return_add_generic_AC_RND_CONV_false_21_if_7_return_add_generic_AC_RND_CONV_false_21_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_21_exception_sva_1 | return_add_generic_AC_RND_CONV_false_12_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1[50:0]),
      return_add_generic_AC_RND_CONV_false_21_if_7_return_add_generic_AC_RND_CONV_false_21_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_70,
      z_out_69, z_out_70[11]);
  assign return_extract_59_return_extract_59_or_2_nl = (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_extract_59_return_extract_59_or_2_nl,
      return_add_generic_AC_RND_CONV_false_21_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_m_r_51_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1[50]), return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0 = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1[50:1]),
      (return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1[49:0]), return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1[0])
      & (~ return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_23_op1_mu_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0,
      and_dcpl_447);
  assign return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_51_lpi_3_dfm_mx0 =
      MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[50]),
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0, and_dcpl_447);
  assign return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[49:0]),
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_447);
  assign return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1,
      and_dcpl_447);
  assign return_add_generic_AC_RND_CONV_false_23_e1_eq_e2_equal_tmp = (stage_PE_1_tmp_re_d_sva[62:52])
      == ({return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1});
  assign return_add_generic_AC_RND_CONV_false_23_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_110[54]))) | (return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (z_out_110[53]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_110[52]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_110[51]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_110[50]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_110[49]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_110[48]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_110[47]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_110[46]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_110[45]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_110[44]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_110[43]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_110[42]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_110[41]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_110[40]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_110[39]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_110[38]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_110[37]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_110[36]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_110[35]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_110[34]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_110[33]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_110[32]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_110[31]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_110[30]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_110[29]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_110[28]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_110[27]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_110[26]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_110[25]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_110[24]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_110[23]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_110[22]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_110[21]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_110[20]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_110[19]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_110[18]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_110[17]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_110[16]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_110[15]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_110[14]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_110[13]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_110[12]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_110[11]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_110[10]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_110[9]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_110[8]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_110[7]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_110[6]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_110[5]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_110[4]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_110[3]))) | (return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_110[2])));
  assign return_add_generic_AC_RND_CONV_false_25_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_107[54]))) | (return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (z_out_107[53]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_107[52]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_107[51]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_107[50]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_107[49]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_107[48]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_107[47]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_107[46]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_107[45]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_107[44]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_107[43]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_107[42]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_107[41]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_107[40]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_107[39]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_107[38]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_107[37]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_107[36]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_107[35]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_107[34]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_107[33]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_107[32]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_107[31]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_107[30]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_107[29]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_107[28]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_107[27]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_107[26]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_107[25]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_107[24]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_107[23]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_107[22]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_107[21]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_107[20]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_107[19]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_107[18]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_107[17]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_107[16]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_107[15]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_107[14]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_107[13]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_107[12]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_107[11]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_107[10]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_107[9]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_107[8]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_107[7]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_107[6]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_107[5]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_107[4]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_107[3]))) | (return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_107[2])));
  assign return_add_generic_AC_RND_CONV_false_23_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_23_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_23_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp
      = ~((return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_21_if_5_or_nl = and_332_cse | return_add_generic_AC_RND_CONV_false_if_5_return_add_generic_AC_RND_CONV_false_if_5_and_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_21_mux_14_nl = MUX_s_1_2_2(and_332_cse,
      return_add_generic_AC_RND_CONV_false_21_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_21_exception_sva_1 = return_add_generic_AC_RND_CONV_false_21_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_21_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_21_mux_14_nl;
  assign return_add_generic_AC_RND_CONV_false_22_if_5_or_nl = and_368_cse | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_22_mux_17_nl = MUX_s_1_2_2(and_368_cse,
      return_add_generic_AC_RND_CONV_false_22_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_22_exception_sva_1 = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_22_mux_17_nl;
  assign return_add_generic_AC_RND_CONV_false_22_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_22_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_23_if_5_or_nl = and_374_cse | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_23_mux_17_nl = MUX_s_1_2_2(and_374_cse,
      return_add_generic_AC_RND_CONV_false_23_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_23_exception_sva_1 = operator_11_true_return_22_sva
      | return_mult_generic_AC_RND_CONV_false_1_op1_zero_sva_1 | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_23_mux_17_nl;
  assign return_add_generic_AC_RND_CONV_false_23_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_23_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_12_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_24_if_5_or_nl = and_382_cse | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_24_mux_10_nl = MUX_s_1_2_2(and_382_cse,
      return_add_generic_AC_RND_CONV_false_24_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_24_exception_sva_1 = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_24_mux_10_nl;
  assign return_add_generic_AC_RND_CONV_false_24_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_24_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_25_if_5_or_nl = and_389_cse | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_25_mux_10_nl = MUX_s_1_2_2(and_389_cse,
      return_add_generic_AC_RND_CONV_false_25_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_25_exception_sva_1 = operator_11_true_return_22_sva
      | operator_11_true_return_26_sva | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_unequal_tmp | return_add_generic_AC_RND_CONV_false_25_mux_10_nl;
  assign return_add_generic_AC_RND_CONV_false_25_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_25_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva;
  assign return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1) | (z_out_106[105]);
  assign return_mult_generic_AC_RND_CONV_false_6_if_if_not_nl = ~ (operator_6_false_58_acc_psp_sva_1[11]);
  assign return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3 = MUX_v_11_2_2(11'b00000000000,
      (operator_6_false_58_acc_psp_sva_1[10:0]), return_mult_generic_AC_RND_CONV_false_6_if_if_not_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp = conv_u2s_11_12(out_f_d_rsci_q_d[62:52])
      + conv_s2s_5_12({4'b1011 , (~ return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp)})
      + 12'b000000000001;
  assign return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp = nl_return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp[11:0];
  assign nl_operator_6_false_58_acc_psp_sva_1 = return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp
      + conv_s2s_7_12({1'b1 , (~ leading_sign_53_0_6_out_1)}) + 12'b000000000001;
  assign operator_6_false_58_acc_psp_sva_1 = nl_operator_6_false_58_acc_psp_sva_1[11:0];
  assign return_mult_generic_AC_RND_CONV_false_6_e_incr_lpi_2_dfm_2 = ~((~(((z_out_106[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((z_out_106[51]) | return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_or_2))
      | (z_out_106[105]))) | (return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp[11]));
  assign return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1
      = ~((out_f_d_rsci_q_d[62:52]==11'b00000000000) & return_extract_3_m_zero_sva_mx1w0);
  assign return_mult_generic_AC_RND_CONV_false_6_lor_lpi_2_dfm_1 = (operator_11_true_3_operator_11_true_3_and_tmp
      & return_extract_3_m_zero_sva_mx1w0) | ((return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3==11'b11111111110)
      & return_mult_generic_AC_RND_CONV_false_6_e_incr_lpi_2_dfm_2) | return_mult_generic_AC_RND_CONV_false_6_op1_nan_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_6_op1_nan_sva_1 = operator_11_true_3_operator_11_true_3_and_tmp
      & (~ return_extract_3_m_zero_sva_mx1w0);
  assign return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1 = (~ return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_6_lor_lpi_2_dfm_1;
  assign return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_6_if_1_and_1_tmp_1 | (return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp[11]));
  assign return_mult_generic_AC_RND_CONV_false_6_and_2_nl = return_mult_generic_AC_RND_CONV_false_6_if_1_and_1_tmp_1
      & (~ (return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp[11]));
  assign return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1 =
      MUX1HOT_v_53_3_2((z_out_106[104:52]), (z_out_106[103:51]), (return_mult_generic_AC_RND_CONV_false_6_else_1_rshift_itm[53:1]),
      {return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_nor_nl
      , return_mult_generic_AC_RND_CONV_false_6_and_2_nl , (return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp[11])});
  assign return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_mux_1_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1,
      return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva, return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp[11]);
  assign return_mult_generic_AC_RND_CONV_false_6_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_mux_1_nl
      & (~ (z_out_106[105]));
  assign nl_stage_monty_mul_acc_2_psp_sva_1 = operator_32_false_2_acc_psp_1_sva_1
      + conv_u2s_14_15(signext_14_13({(operator_32_false_2_acc_psp_1_sva_1[14]) ,
      11'b00000000000 , (operator_32_false_2_acc_psp_1_sva_1[14])}));
  assign stage_monty_mul_acc_2_psp_sva_1 = nl_stage_monty_mul_acc_2_psp_sva_1[14:0];
  assign nl_operator_32_false_2_acc_2_nl = conv_s2u_23_24({z_out_113 , (in_u_rsci_q_d[11:0])})
      + ({z_out_101 , 4'b0000 , z_out_101});
  assign operator_32_false_2_acc_2_nl = nl_operator_32_false_2_acc_2_nl[23:0];
  assign nl_operator_32_false_2_acc_psp_1_sva_1 = conv_u2s_14_15(readslicef_24_14_10(operator_32_false_2_acc_2_nl))
      + 15'b100111111111111;
  assign operator_32_false_2_acc_psp_1_sva_1 = nl_operator_32_false_2_acc_psp_1_sva_1[14:0];
  assign return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_9
      = (operator_33_true_12_acc_psp_sva[0]) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_11
      = MUX_v_10_2_2(10'b0000000000, (operator_33_true_12_acc_psp_sva[10:1]), return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva);
  assign return_add_generic_AC_RND_CONV_false_1_if_5_or_3 = return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva
      | (~((operator_33_true_12_acc_psp_sva!=13'b0000000000000)));
  assign return_add_generic_AC_RND_CONV_false_1_mux_28 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva,
      return_add_generic_AC_RND_CONV_false_1_if_5_or_3, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_1_mux_30 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_9,
      return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_2_cse,
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_if_5_return_add_generic_AC_RND_CONV_false_if_5_and_1_tmp
      = (return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_5_cse[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_2_cse
      & (return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_5_cse[11:10]==2'b00);
  assign nl_return_mult_generic_AC_RND_CONV_false_1_if_acc_2_nl = -(z_out_111[12:0]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_acc_2_nl = nl_return_mult_generic_AC_RND_CONV_false_1_if_acc_2_nl[12:0];
  assign return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1 = readslicef_13_1_12(return_mult_generic_AC_RND_CONV_false_1_if_acc_2_nl);
  assign return_mult_generic_AC_RND_CONV_false_1_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_1_exp_ovf_oif_aelse_and_1_tmp
      = (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1==12'b011111111110)
      & return_mult_generic_AC_RND_CONV_false_1_e_incr_lpi_3_dfm_2;
  assign return_mult_generic_AC_RND_CONV_false_else_2_else_else_mux_2 = MUX_v_11_2_2((return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[10:0]),
      (return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_acc_tmp[10:0]), return_mult_generic_AC_RND_CONV_false_1_e_incr_lpi_3_dfm_2);
  assign nl_return_add_generic_AC_RND_CONV_false_17_acc_3_nl = -(z_out_102[10:0]);
  assign return_add_generic_AC_RND_CONV_false_17_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_17_acc_3_nl[10:0];
  assign return_add_generic_AC_RND_CONV_false_17_acc_3_itm_10 = readslicef_11_1_10(return_add_generic_AC_RND_CONV_false_17_acc_3_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_8_acc_3_nl = -(z_out_85[11:0]);
  assign return_add_generic_AC_RND_CONV_false_8_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_8_acc_3_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_8_acc_3_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_15_acc_3_nl = -(z_out_85[11:0]);
  assign return_add_generic_AC_RND_CONV_false_15_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_15_acc_3_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_15_acc_3_nl);
  assign return_add_generic_AC_RND_CONV_false_4_sticky_bit_and_158 = return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm
      & (~ (z_out_109[2]));
  assign return_add_generic_AC_RND_CONV_false_6_mux_36 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_9,
      operator_6_false_17_acc_itm_0, z_out_89[53]);
  assign nl_return_add_generic_AC_RND_CONV_false_16_acc_3_nl = -(operator_33_true_32_acc_tmp[11:0]);
  assign return_add_generic_AC_RND_CONV_false_16_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_16_acc_3_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_16_acc_3_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_16_acc_3_nl);
  assign return_add_generic_AC_RND_CONV_false_3_return_add_generic_AC_RND_CONV_false_3_and_9
      = (operator_33_true_32_acc_tmp[0]) & return_add_generic_AC_RND_CONV_false_16_acc_3_itm_11_1;
  assign nl_return_add_generic_AC_RND_CONV_false_18_acc_3_nl = -(z_out_102[10:0]);
  assign return_add_generic_AC_RND_CONV_false_18_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_18_acc_3_nl[10:0];
  assign return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1 = readslicef_11_1_10(return_add_generic_AC_RND_CONV_false_18_acc_3_nl);
  assign return_add_generic_AC_RND_CONV_false_18_if_5_return_add_generic_AC_RND_CONV_false_18_if_5_nor_2
      = ~((operator_33_true_36_acc_psp_1_sva!=12'b000000000000));
  assign return_add_generic_AC_RND_CONV_false_17_if_5_return_add_generic_AC_RND_CONV_false_17_if_5_nor_2
      = ~((operator_32_false_1_acc_psp_sva_11_0!=12'b000000000000));
  assign return_add_generic_AC_RND_CONV_false_2_aif_equal_tmp = ({return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1
      , return_extract_2_mux_4_cse , return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1})
      == ({drf_qr_lval_13_smx_0_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_13_op2_mu_0_lpi_3_dfm_1});
  assign return_add_generic_AC_RND_CONV_false_15_aif_equal_tmp = ({return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_1
      , return_extract_33_mux_3_cse , return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1})
      == ({drf_qr_lval_13_smx_0_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_13_op2_mu_0_lpi_3_dfm_1});
  assign and_dcpl_18 = mode_lpi_1_dfm & (~ inverse_lpi_1_dfm_1);
  assign or_tmp_21 = (~ (z_out_86[12])) | operator_11_true_47_operator_11_true_47_and_tmp
      | return_mult_generic_AC_RND_CONV_false_3_op2_zero_sva_1 | operator_11_true_return_1_sva;
  assign or_tmp_26 = (~ (z_out_86[12])) | operator_11_true_15_operator_11_true_15_and_tmp
      | return_mult_generic_AC_RND_CONV_false_op2_zero_sva_1 | operator_11_true_return_1_sva;
  assign or_tmp_30 = (((~ (z_out_86[12])) | operator_11_true_47_operator_11_true_47_and_tmp
      | return_extract_47_return_extract_47_nor_tmp) & return_extract_15_return_extract_15_nor_tmp
      & return_extract_47_m_zero_return_extract_47_m_zero_nor_tmp) | operator_11_true_return_1_sva;
  assign or_82_cse = (~ (z_out_86[12])) | operator_11_true_15_operator_11_true_15_and_tmp;
  assign mux_tmp_12 = MUX_s_1_2_2(or_tmp_30, or_tmp_21, or_82_cse);
  assign or_87_cse = (~ (z_out_86[12])) | operator_11_true_49_operator_11_true_49_and_tmp;
  assign mux_14_nl = MUX_s_1_2_2(operator_11_true_return_1_sva, or_tmp_30, or_87_cse);
  assign mux_13_nl = MUX_s_1_2_2(operator_11_true_return_1_sva, or_tmp_21, or_87_cse);
  assign mux_tmp_15 = MUX_s_1_2_2(mux_14_nl, mux_13_nl, or_82_cse);
  assign or_81_cse = (~ (z_out_86[12])) | operator_11_true_17_operator_11_true_17_and_tmp;
  assign mux_17_nl = MUX_s_1_2_2(mux_tmp_15, mux_tmp_12, return_extract_49_return_extract_49_nor_tmp);
  assign mux_18_nl = MUX_s_1_2_2(operator_11_true_return_1_sva, mux_17_nl, return_mult_generic_AC_RND_CONV_false_1_op2_zero_sva_1);
  assign mux_16_nl = MUX_s_1_2_2(mux_tmp_15, mux_tmp_12, return_mult_generic_AC_RND_CONV_false_4_op2_zero_sva_1);
  assign mux_tmp_19 = MUX_s_1_2_2(mux_18_nl, mux_16_nl, or_81_cse);
  assign mux_10_nl = MUX_s_1_2_2(operator_11_true_return_1_sva, or_tmp_26, return_mult_generic_AC_RND_CONV_false_1_op2_zero_sva_1);
  assign mux_11_nl = MUX_s_1_2_2(mux_10_nl, or_tmp_26, or_81_cse);
  assign mux_20_nl = MUX_s_1_2_2(mux_tmp_19, mux_11_nl, return_extract_21_m_zero_sva);
  assign or_72_nl = return_mult_generic_AC_RND_CONV_false_4_op2_zero_sva_1 | (~ (z_out_86[12]))
      | operator_11_true_49_operator_11_true_49_and_tmp;
  assign mux_9_nl = MUX_s_1_2_2(operator_11_true_return_1_sva, or_tmp_21, or_72_nl);
  assign or_76_nl = return_extract_21_m_zero_sva | mux_9_nl;
  assign mux_21_nl = MUX_s_1_2_2(mux_20_nl, or_76_nl, return_extract_12_m_zero_sva);
  assign mux_tmp_22 = MUX_s_1_2_2(mux_tmp_19, mux_21_nl, operator_11_true_return_21_sva);
  assign and_tmp_1 = (return_extract_51_and_cse | (~ (z_out_68[12])) | operator_11_true_51_operator_11_true_51_and_tmp
      | return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1) & mux_tmp_22;
  assign and_dcpl_57 = ~(return_add_generic_AC_RND_CONV_false_14_op1_nan_sva | return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva);
  assign and_dcpl_64 = ~(return_add_generic_AC_RND_CONV_false_10_op1_nan_sva | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign or_dcpl_93 = operator_11_true_return_26_sva | return_add_generic_AC_RND_CONV_false_10_unequal_tmp;
  assign and_dcpl_75 = ~(operator_11_true_return_26_sva | return_add_generic_AC_RND_CONV_false_10_unequal_tmp);
  assign nor_34_cse = ~((fsm_output[52]) | (fsm_output[27]));
  assign nor_35_cse = ~((fsm_output[54:53]!=2'b00));
  assign and_225_cse = mode_lpi_1_dfm & BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm;
  assign nl_for_acc_nl = conv_u2s_3_4(for_i_3_0_sva_2[3:1]) + 4'b1011;
  assign for_acc_nl = nl_for_acc_nl[3:0];
  assign and_dcpl_159 = or_2748_cse & (~((~(t_in_10_0_lpi_1_dfm_1_1 & (~(t_in_10_0_lpi_1_dfm_1_10
      | t_in_10_0_lpi_1_dfm_1_9 | t_in_10_0_lpi_1_dfm_1_8 | t_in_10_0_lpi_1_dfm_1_7
      | t_in_10_0_lpi_1_dfm_1_6 | t_in_10_0_lpi_1_dfm_1_5 | t_in_10_0_lpi_1_dfm_1_4
      | t_in_10_0_lpi_1_dfm_1_3 | t_in_10_0_lpi_1_dfm_1_2)))) & (readslicef_4_1_3(for_acc_nl))));
  assign and_dcpl_160 = ~(and_225_cse | (z_out_101[9]));
  assign and_dcpl_166 = (operator_16_false_io_read_mode1_rsc_cse_sva[14:11]==4'b0000);
  assign and_dcpl_172 = ~((operator_16_false_io_read_mode1_rsc_cse_sva[3:2]!=2'b00));
  assign and_dcpl_175 = and_dcpl_172 & (operator_16_false_io_read_mode1_rsc_cse_sva[10:4]==7'b0000000);
  assign or_dcpl_179 = (operator_16_false_io_read_mode1_rsc_cse_sva[1:0]!=2'b01);
  assign or_dcpl_180 = (operator_16_false_io_read_mode1_rsc_cse_sva[15:14]!=2'b00);
  assign or_dcpl_184 = (operator_16_false_io_read_mode1_rsc_cse_sva[13:10]!=4'b0000);
  assign or_dcpl_190 = (operator_16_false_io_read_mode1_rsc_cse_sva[3:2]!=2'b00);
  assign or_dcpl_192 = or_dcpl_190 | (operator_16_false_io_read_mode1_rsc_cse_sva[9:4]!=6'b000000);
  assign and_dcpl_177 = ~((~(or_dcpl_192 | or_dcpl_184 | or_dcpl_180 | or_dcpl_179))
      | operator_16_false_operator_16_false_nor_cse_sva);
  assign and_dcpl_183 = ~((~(or_dcpl_192 | or_dcpl_184 | or_dcpl_180 | (~((operator_16_false_io_read_mode1_rsc_cse_sva[1])
      ^ (operator_16_false_io_read_mode1_rsc_cse_sva[0]))))) | operator_16_false_operator_16_false_nor_cse_sva);
  assign or_dcpl_198 = (fsm_output[3]) | (fsm_output[28]);
  assign or_dcpl_200 = (fsm_output[5:4]!=2'b00);
  assign or_dcpl_201 = (fsm_output[30:29]!=2'b00);
  assign or_dcpl_204 = (fsm_output[4:3]!=2'b00);
  assign or_dcpl_207 = (fsm_output[54:53]!=2'b00);
  assign and_dcpl_185 = ~(mode_lpi_1_dfm | inverse_lpi_1_dfm_1);
  assign or_dcpl_208 = (fsm_output[11:10]!=2'b00);
  assign or_dcpl_209 = (fsm_output[46]) | (fsm_output[48]);
  assign or_dcpl_221 = (fsm_output[35:34]!=2'b00);
  assign or_dcpl_223 = (fsm_output[43]) | (fsm_output[41]);
  assign or_dcpl_224 = (fsm_output[42]) | (fsm_output[44]);
  assign or_dcpl_227 = (and_dcpl_172 & (~((operator_16_false_io_read_mode1_rsc_cse_sva[5:4]!=2'b00)))
      & (~((operator_16_false_io_read_mode1_rsc_cse_sva[7:6]!=2'b00))) & (~((operator_16_false_io_read_mode1_rsc_cse_sva[9:8]!=2'b00)))
      & (~((operator_16_false_io_read_mode1_rsc_cse_sva[11:10]!=2'b00))) & (~((operator_16_false_io_read_mode1_rsc_cse_sva[13:12]!=2'b00)))
      & (~((operator_16_false_io_read_mode1_rsc_cse_sva[15:14]!=2'b00))) & (~ (operator_16_false_io_read_mode1_rsc_cse_sva[1]))
      & (operator_16_false_io_read_mode1_rsc_cse_sva[0])) | operator_16_false_operator_16_false_nor_cse_sva;
  assign or_dcpl_228 = (fsm_output[30]) | (fsm_output[8]);
  assign or_dcpl_230 = (fsm_output[29:28]!=2'b00);
  assign or_dcpl_233 = (fsm_output[32:31]!=2'b00);
  assign or_dcpl_235 = (fsm_output[36:35]!=2'b00);
  assign or_dcpl_236 = (fsm_output[21:20]!=2'b00);
  assign or_dcpl_239 = (fsm_output[22]) | (fsm_output[25]);
  assign or_dcpl_240 = or_dcpl_239 | (fsm_output[24]);
  assign or_dcpl_245 = (fsm_output[10:9]!=2'b00);
  assign or_dcpl_248 = (fsm_output[19:18]!=2'b00);
  assign and_dcpl_202 = ~((fsm_output[0]) | (fsm_output[56]));
  assign or_dcpl_253 = (fsm_output[47]) | (fsm_output[49]);
  assign or_dcpl_269 = (fsm_output[9:8]!=2'b00);
  assign or_dcpl_272 = (fsm_output[24]) | (fsm_output[20]);
  assign or_dcpl_273 = (fsm_output[26]) | (fsm_output[22]);
  assign or_dcpl_283 = ~(reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd
      & return_add_generic_AC_RND_CONV_false_if_5_return_add_generic_AC_RND_CONV_false_if_5_and_1_tmp);
  assign and_dcpl_203 = stage_PE_1_and_1_tmp & or_dcpl_283;
  assign and_dcpl_204 = ~(operator_11_true_return_1_sva | operator_11_true_return_21_sva);
  assign or_dcpl_284 = ~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_1_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva);
  assign and_275_cse = reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd
      & return_add_generic_AC_RND_CONV_false_if_5_return_add_generic_AC_RND_CONV_false_if_5_and_1_tmp;
  assign or_dcpl_285 = and_275_cse | operator_11_true_return_21_sva;
  assign or_dcpl_289 = ~(mode_lpi_1_dfm & inverse_lpi_1_dfm_1);
  assign and_dcpl_210 = mode_lpi_1_dfm & (~ (operator_14_false_1_acc_psp_sva_12_10[2]));
  assign or_dcpl_296 = (~ inverse_lpi_1_dfm_1) | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva;
  assign and_dcpl_216 = return_add_generic_AC_RND_CONV_false_2_if_5_return_add_generic_AC_RND_CONV_false_2_if_5_and_tmp
      & (z_out_89[53]);
  assign or_dcpl_301 = or_dcpl_93 | return_add_generic_AC_RND_CONV_false_22_op1_inf_sva;
  assign and_dcpl_217 = (z_out_89[53]) & return_add_generic_AC_RND_CONV_false_3_if_5_return_add_generic_AC_RND_CONV_false_3_if_5_and_tmp;
  assign or_dcpl_308 = or_dcpl_289 | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva;
  assign or_dcpl_311 = operator_11_true_return_22_sva | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva;
  assign or_dcpl_312 = or_dcpl_311 | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva;
  assign and_dcpl_219 = mode_lpi_1_dfm & (~ return_add_generic_AC_RND_CONV_false_10_op1_nan_sva);
  assign or_dcpl_320 = ~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva);
  assign and_dcpl_222 = ~(operator_11_true_return_22_sva | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva);
  assign and_dcpl_223 = and_dcpl_222 & (~ return_add_generic_AC_RND_CONV_false_10_op2_nan_sva);
  assign and_dcpl_224 = and_dcpl_223 & (~(return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm
      & (z_out_89[53])));
  assign or_dcpl_324 = or_dcpl_312 | (return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm
      & (z_out_89[53]));
  assign and_dcpl_229 = (~ operator_11_true_return_21_sva) & mode_lpi_1_dfm & or_dcpl_283;
  assign and_dcpl_231 = ~(((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_7_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva)
      | operator_11_true_return_1_sva);
  assign and_dcpl_235 = (~ return_add_generic_AC_RND_CONV_false_10_op2_nan_sva) &
      mode_lpi_1_dfm & or_dcpl_283;
  assign and_dcpl_237 = (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_8_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
      & and_dcpl_222;
  assign or_dcpl_337 = return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva
      | and_275_cse;
  assign or_dcpl_342 = ~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_14_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva);
  assign and_dcpl_251 = (z_out_89[53]) & return_add_generic_AC_RND_CONV_false_15_if_5_return_add_generic_AC_RND_CONV_false_15_if_5_and_tmp;
  assign or_dcpl_359 = return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva;
  assign and_dcpl_253 = (z_out_89[53]) & return_add_generic_AC_RND_CONV_false_16_if_5_return_add_generic_AC_RND_CONV_false_16_if_5_and_tmp;
  assign or_dcpl_367 = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva;
  assign or_dcpl_371 = ~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva);
  assign and_dcpl_259 = ~(((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_20_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva)
      | operator_11_true_return_1_sva);
  assign and_dcpl_263 = (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_21_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
      & and_dcpl_222;
  assign and_dcpl_266 = and_dcpl_18 & (~ return_add_generic_AC_RND_CONV_false_14_op1_nan_sva);
  assign and_dcpl_268 = ~(operator_11_true_return_1_sva | return_add_generic_AC_RND_CONV_false_22_op1_inf_sva);
  assign and_dcpl_274 = and_dcpl_18 & (~ return_add_generic_AC_RND_CONV_false_10_op1_nan_sva);
  assign and_dcpl_276 = ~(operator_11_true_return_21_sva | operator_11_true_return_22_sva);
  assign and_dcpl_285 = and_dcpl_75 & (~ return_add_generic_AC_RND_CONV_false_22_op1_inf_sva);
  assign or_dcpl_438 = operator_11_true_return_22_sva | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva;
  assign and_dcpl_323 = and_dcpl_202 & (~ (fsm_output[1]));
  assign and_dcpl_327 = ~((fsm_output[55:53]!=3'b000));
  assign and_dcpl_329 = ~((fsm_output[2:1]!=2'b00));
  assign and_dcpl_330 = and_dcpl_202 & and_dcpl_329;
  assign and_dcpl_333 = ~((fsm_output[2]) | (fsm_output[55]));
  assign or_dcpl_466 = (fsm_output[33:32]!=2'b00);
  assign or_dcpl_470 = (fsm_output[18:17]!=2'b00);
  assign or_dcpl_473 = (fsm_output[21]) | (fsm_output[43]);
  assign or_dcpl_476 = (fsm_output[19]) | (fsm_output[23]);
  assign and_dcpl_340 = ~(and_435_cse | (z_out_96[11]));
  assign and_dcpl_341 = ~(and_528_cse | (z_out_69[11]));
  assign and_dcpl_344 = ~((fsm_output[53]) | (fsm_output[8]));
  assign and_dcpl_354 = ~((fsm_output[18:17]!=2'b00));
  assign and_dcpl_360 = ~((fsm_output[44]) | (fsm_output[19]));
  assign and_dcpl_369 = ~((fsm_output[4]) | (fsm_output[29]));
  assign and_dcpl_382 = ~((fsm_output[25:24]!=2'b00));
  assign and_dcpl_389 = ~((fsm_output[2]) | (fsm_output[47]));
  assign and_dcpl_393 = ~((fsm_output[51:50]!=2'b00));
  assign or_dcpl_484 = (fsm_output[12]) | (fsm_output[37]);
  assign and_dcpl_402 = ~((fsm_output[28]) | (fsm_output[0]));
  assign and_dcpl_403 = ~((fsm_output[3]) | (fsm_output[26]));
  assign and_dcpl_405 = and_dcpl_393 & nor_34_cse;
  assign and_dcpl_420 = and_dcpl_403 & (~ (fsm_output[28]));
  assign and_dcpl_421 = and_dcpl_405 & and_dcpl_420;
  assign or_dcpl_485 = (fsm_output[42]) | (fsm_output[17]);
  assign or_dcpl_492 = (fsm_output[8]) | (fsm_output[12]);
  assign or_dcpl_493 = (fsm_output[15]) | (fsm_output[40]);
  assign or_dcpl_497 = operator_6_false_17_or_cse | return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse;
  assign or_dcpl_502 = (fsm_output[39]) | (fsm_output[17]);
  assign or_dcpl_503 = (fsm_output[42]) | (fsm_output[14]);
  assign or_dcpl_504 = or_dcpl_503 | or_dcpl_502;
  assign or_dcpl_509 = (fsm_output[11]) | (fsm_output[8]);
  assign or_dcpl_511 = (fsm_output[38]) | (fsm_output[15]);
  assign or_dcpl_515 = (fsm_output[16]) | (fsm_output[7]);
  assign or_dcpl_516 = (fsm_output[21]) | (fsm_output[14]);
  assign or_dcpl_519 = (fsm_output[20:19]!=2'b00);
  assign or_dcpl_520 = (fsm_output[46:45]!=2'b00);
  assign or_dcpl_521 = or_dcpl_520 | (fsm_output[44]);
  assign or_dcpl_522 = or_dcpl_521 | or_dcpl_519;
  assign and_dcpl_446 = ~(return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_and_cse
      | (z_out_95[11]));
  assign and_dcpl_447 = ~(and_606_cse | (z_out_70[11]));
  assign or_dcpl_528 = (fsm_output[30]) | (fsm_output[40]) | (fsm_output[5]);
  assign or_dcpl_529 = (fsm_output[7]) | (fsm_output[13]);
  assign or_dcpl_532 = (fsm_output[14]) | (fsm_output[18]);
  assign or_dcpl_534 = (fsm_output[44]) | (fsm_output[19]);
  assign or_dcpl_535 = or_dcpl_520 | or_dcpl_534;
  assign or_dcpl_545 = (fsm_output[25:24]!=2'b00);
  assign or_dcpl_553 = (fsm_output[8]) | (fsm_output[33]);
  assign or_dcpl_554 = or_dcpl_553 | or_dcpl_484;
  assign or_dcpl_555 = (fsm_output[40]) | (fsm_output[11]);
  assign or_dcpl_559 = (fsm_output[10]) | (fsm_output[13]);
  assign or_dcpl_560 = (fsm_output[9]) | (fsm_output[35]);
  assign or_dcpl_562 = (fsm_output[16]) | (fsm_output[34]);
  assign and_dcpl_448 = ~(return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_and_1_cse
      | (z_out_70[11]));
  assign and_dcpl_452 = ~(return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_and_1_cse
      | (z_out_95[11]));
  assign or_dcpl_573 = ~(return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp
      & return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_itm_52);
  assign or_dcpl_575 = (fsm_output[32]) | (fsm_output[12]);
  assign or_dcpl_576 = or_dcpl_575 | (fsm_output[37]);
  assign or_dcpl_579 = (fsm_output[36]) | (fsm_output[40]);
  assign or_dcpl_580 = or_dcpl_579 | (fsm_output[11]);
  assign or_dcpl_584 = operator_6_false_17_or_cse | (fsm_output[13]);
  assign or_dcpl_585 = (fsm_output[34]) | (fsm_output[7]);
  assign or_dcpl_586 = or_dcpl_585 | (fsm_output[9]);
  assign or_dcpl_588 = (fsm_output[17]) | (fsm_output[41]);
  assign or_dcpl_590 = or_dcpl_503 | (fsm_output[39]);
  assign and_dcpl_460 = ~(and_526_cse | (return_add_generic_AC_RND_CONV_false_17_e_dif_acc_tmp[10]));
  assign or_dcpl_596 = (fsm_output[33]) | (fsm_output[6]);
  assign or_dcpl_597 = or_dcpl_596 | or_dcpl_233;
  assign or_dcpl_598 = (fsm_output[8:7]!=2'b00);
  assign or_dcpl_602 = (fsm_output[48]) | (fsm_output[44]);
  assign or_dcpl_604 = (fsm_output[46]) | (fsm_output[42]);
  assign or_dcpl_605 = (fsm_output[45]) | (fsm_output[47]);
  assign or_dcpl_606 = or_dcpl_605 | or_dcpl_604;
  assign or_dcpl_618 = (fsm_output[49]) | (fsm_output[46]);
  assign or_dcpl_619 = (fsm_output[50]) | (fsm_output[45]);
  assign or_dcpl_620 = or_dcpl_619 | (fsm_output[47]);
  assign or_dcpl_621 = or_dcpl_620 | or_dcpl_618;
  assign or_dcpl_625 = (fsm_output[43]) | (fsm_output[18]);
  assign or_dcpl_626 = or_dcpl_625 | (fsm_output[17]);
  assign or_dcpl_627 = or_dcpl_224 | (fsm_output[19]);
  assign or_dcpl_628 = or_dcpl_627 | or_dcpl_626;
  assign and_dcpl_466 = ~(return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_and_1_cse
      | (z_out_69[11]));
  assign and_dcpl_467 = ~(return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_20_e_dif1_acc_2_tmp[11]));
  assign and_dcpl_468 = or_dcpl_573 & (~ (z_out_70[11]));
  assign and_dcpl_469 = ~(return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_21_op1_smaller_oelse_and_cse
      | (return_add_generic_AC_RND_CONV_false_21_e_dif1_acc_2_tmp[11]));
  assign or_dcpl_632 = (fsm_output[6]) | (fsm_output[32]);
  assign or_dcpl_633 = or_dcpl_632 | (fsm_output[31]);
  assign or_dcpl_634 = or_dcpl_598 | (fsm_output[33]);
  assign or_dcpl_635 = or_dcpl_634 | or_dcpl_633;
  assign or_dcpl_640 = or_dcpl_484 | (fsm_output[31]);
  assign or_dcpl_645 = or_dcpl_585 | or_dcpl_560;
  assign or_dcpl_654 = (fsm_output[17]) | (fsm_output[34]);
  assign or_dcpl_664 = or_dcpl_534 | (fsm_output[43]);
  assign and_dcpl_474 = ~(return_add_generic_AC_RND_CONV_false_11_do_sub_sva | return_mult_generic_AC_RND_CONV_false_1_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_1_exp_ovf_oif_aelse_and_1_tmp);
  assign and_dcpl_475 = and_dcpl_474 & (~((return_mult_generic_AC_RND_CONV_false_1_exp_plus_1_acc_tmp[11])
      | return_add_generic_AC_RND_CONV_false_17_mux_6_itm));
  assign and_dcpl_478 = ~(operator_11_true_return_22_sva | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign and_dcpl_479 = ~(return_add_generic_AC_RND_CONV_false_11_do_sub_sva | return_mult_generic_AC_RND_CONV_false_1_exp_ovf_return_mult_generic_AC_RND_CONV_false_1_exp_ovf_or_tmp);
  assign or_dcpl_671 = or_dcpl_545 | (fsm_output[20]);
  assign or_dcpl_673 = or_dcpl_476 | (fsm_output[22]);
  assign or_dcpl_678 = or_dcpl_553 | (fsm_output[6]);
  assign or_dcpl_679 = or_dcpl_678 | or_dcpl_233;
  assign or_dcpl_680 = (fsm_output[36]) | (fsm_output[11]);
  assign or_dcpl_684 = ~(return_add_generic_AC_RND_CONV_false_17_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_4_op1_mu_52_lpi_3_dfm_1 , stage_PE_gm_re_d_mux_cse
      , return_add_generic_AC_RND_CONV_false_4_op1_mu_0_lpi_3_dfm_1}) == ({stage_PE_gm_im_d_mux_cse
      , stage_PE_gm_im_d_mux_2_cse , return_add_generic_AC_RND_CONV_false_4_op2_mu_0_lpi_3_dfm_1})));
  assign or_dcpl_685 = (fsm_output[40]) | (fsm_output[8]);
  assign or_dcpl_686 = (fsm_output[10]) | (fsm_output[15]);
  assign or_dcpl_698 = (fsm_output[7]) | (fsm_output[9]);
  assign or_dcpl_699 = or_dcpl_698 | (fsm_output[35]);
  assign or_dcpl_702 = or_dcpl_470 | (fsm_output[41]);
  assign or_dcpl_708 = ~((({return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm
      , return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1 , return_extract_2_mux_4_cse
      , return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1})) & return_add_generic_AC_RND_CONV_false_1_e1_eq_e2_equal_tmp);
  assign or_dcpl_709 = ~((({drf_qr_lval_13_smx_0_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_10_op2_mu_1_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_10_op2_mu_1_50_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1})) & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_equal_tmp);
  assign and_dcpl_501 = (~(return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp
      & return_add_generic_AC_RND_CONV_false_15_aif_equal_tmp)) & inverse_lpi_1_dfm_1;
  assign or_dcpl_711 = ~((({return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1}))
      & return_add_generic_AC_RND_CONV_false_22_e1_eq_e2_equal_tmp);
  assign or_dcpl_719 = or_dcpl_685 | (fsm_output[33]);
  assign or_dcpl_725 = (fsm_output[23:22]!=2'b00);
  assign or_dcpl_726 = or_dcpl_725 | (fsm_output[20]);
  assign or_dcpl_728 = or_dcpl_602 | (fsm_output[19]);
  assign or_dcpl_740 = or_dcpl_605 | (fsm_output[46]);
  assign or_dcpl_744 = (fsm_output[37]) | (fsm_output[31]);
  assign or_dcpl_750 = (fsm_output[9]) | (fsm_output[13]);
  assign or_dcpl_762 = (fsm_output[42]) | (fsm_output[48]);
  assign or_dcpl_763 = (fsm_output[47:46]!=2'b00);
  assign or_dcpl_776 = (fsm_output[40]) | (fsm_output[32]);
  assign or_dcpl_788 = or_dcpl_236 | (fsm_output[43]);
  assign or_dcpl_789 = or_dcpl_627 | or_dcpl_788;
  assign or_dcpl_800 = or_dcpl_619 | or_dcpl_253;
  assign or_dcpl_809 = or_dcpl_763 | (fsm_output[42]);
  assign and_dcpl_503 = (~(operator_11_true_return_21_sva | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva))
      & or_dcpl_283;
  assign or_dcpl_845 = or_dcpl_598 | or_dcpl_466;
  assign or_dcpl_848 = or_dcpl_534 | or_dcpl_725;
  assign or_dcpl_849 = or_dcpl_740 | or_dcpl_762 | or_dcpl_848;
  assign or_dcpl_854 = ~((~((~ (operator_33_true_32_acc_tmp[11])) & return_add_generic_AC_RND_CONV_false_16_else_4_return_add_generic_AC_RND_CONV_false_16_else_4_nand_tmp))
      & return_add_generic_AC_RND_CONV_false_16_acc_3_itm_11_1);
  assign or_dcpl_866 = or_dcpl_620 | or_dcpl_618 | (fsm_output[48]);
  assign or_dcpl_870 = or_dcpl_553 | (fsm_output[32]);
  assign or_dcpl_874 = or_dcpl_654 | (fsm_output[7]);
  assign or_dcpl_876 = (fsm_output[42]) | (fsm_output[43]) | (fsm_output[18]);
  assign or_dcpl_890 = or_dcpl_698 | (fsm_output[8]) | or_dcpl_466;
  assign or_dcpl_906 = (fsm_output[11]) | (fsm_output[33]);
  assign or_dcpl_928 = or_dcpl_520 | or_dcpl_224;
  assign or_dcpl_933 = (fsm_output[41]) | (fsm_output[34]);
  assign or_dcpl_943 = (fsm_output[16]) | (fsm_output[35]);
  assign or_dcpl_967 = ~(return_add_generic_AC_RND_CONV_false_e1_eq_e2_equal_tmp
      & return_add_generic_AC_RND_CONV_false_2_aif_equal_tmp);
  assign or_dcpl_970 = (fsm_output[15]) | (fsm_output[36]);
  assign or_dcpl_980 = ~(return_add_generic_AC_RND_CONV_false_9_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_23_op1_mu_52_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1})));
  assign or_dcpl_981 = ~(return_add_generic_AC_RND_CONV_false_14_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm
      , return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_1 , return_extract_33_mux_3_cse
      , return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1})));
  assign or_dcpl_982 = ~((({return_add_generic_AC_RND_CONV_false_23_op1_mu_52_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1}))
      & return_add_generic_AC_RND_CONV_false_23_e1_eq_e2_equal_tmp);
  assign and_dcpl_531 = ~(return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_6_op1_smaller_oelse_and_cse
      | (z_out_95[11]));
  assign and_dcpl_534 = (~ return_add_generic_AC_RND_CONV_false_14_op1_nan_sva) &
      return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1;
  assign and_dcpl_541 = (~(return_add_generic_AC_RND_CONV_false_10_op2_nan_sva |
      return_add_generic_AC_RND_CONV_false_12_r_zero_1_sva)) & or_dcpl_283;
  assign and_dcpl_543 = ~(return_add_generic_AC_RND_CONV_false_19_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_19_op1_smaller_oelse_and_cse
      | (z_out_69[11]));
  assign or_tmp_64 = operator_16_false_operator_16_false_nor_cse_sva & (fsm_output[54]);
  assign and_630_cse = and_dcpl_183 & (fsm_output[54]);
  assign and_647_cse = and_6_cse & (fsm_output[31]);
  assign and_660_cse = and_dcpl_177 & or_dcpl_207;
  assign and_662_cse = and_6_cse & (fsm_output[6]);
  assign and_680_cse = inverse_lpi_1_dfm_1 & (fsm_output[32]);
  assign and_741_cse = and_dcpl_177 & (fsm_output[53]);
  assign and_746_cse = inverse_lpi_1_dfm_1 & (fsm_output[7]);
  assign and_836_cse = ~(return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1 &
      mode_lpi_1_dfm);
  assign and_840_cse = ~(mode_lpi_1_dfm & return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1);
  assign or_tmp_231 = (~ inverse_lpi_1_dfm_1) & (fsm_output[2]);
  assign or_tmp_334 = (fsm_output[29]) | (fsm_output[32]);
  assign or_tmp_450 = (fsm_output[46]) | (fsm_output[21]);
  assign or_tmp_759 = (fsm_output[22]) | (fsm_output[16]) | or_dcpl_596;
  assign or_tmp_762 = (fsm_output[45]) | (fsm_output[37]);
  assign and_2185_cse = return_add_generic_AC_RND_CONV_false_8_op1_smaller_return_add_generic_AC_RND_CONV_false_8_op1_smaller_or_cse
      & (fsm_output[14]);
  assign and_2184_cse = return_add_generic_AC_RND_CONV_false_21_op1_smaller_return_add_generic_AC_RND_CONV_false_21_op1_smaller_or_cse
      & (fsm_output[39]);
  assign or_tmp_946 = return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse
      & (fsm_output[18]);
  assign out1_rsci_idat_63_0_mx0c1 = and_dcpl_175 & and_dcpl_166 & (~((operator_16_false_io_read_mode1_rsc_cse_sva[15])
      | (operator_16_false_io_read_mode1_rsc_cse_sva[1]))) & (operator_16_false_io_read_mode1_rsc_cse_sva[0])
      & (~ operator_16_false_operator_16_false_nor_cse_sva) & (fsm_output[54]);
  assign out1_rsci_idat_63_0_mx0c2 = and_dcpl_177 & (fsm_output[54]);
  assign out1_rsci_idat_79_64_mx0c1 = and_dcpl_175 & and_dcpl_166 & (~ (operator_16_false_io_read_mode1_rsc_cse_sva[15]))
      & (operator_16_false_io_read_mode1_rsc_cse_sva[1]) & (~((operator_16_false_io_read_mode1_rsc_cse_sva[0])
      | operator_16_false_operator_16_false_nor_cse_sva)) & (fsm_output[54]);
  assign BUTTERFLY_1_i_9_0_sva_mx0c3 = (fsm_output[50]) | (fsm_output[46]) | (fsm_output[25])
      | (fsm_output[21]);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx8c1 = ~(return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp
      | inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx8c2 = or_dcpl_573
      & (~ (z_out_70[11])) & inverse_lpi_1_dfm_1;
  assign BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx0c8 = (fsm_output[50])
      | (fsm_output[25]);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_mx1c2 = or_dcpl_627
      | (fsm_output[43]) | (fsm_output[14]) | (fsm_output[18]) | or_dcpl_502 | (fsm_output[41])
      | (fsm_output[16]) | (fsm_output[13]) | (fsm_output[38]);
  assign return_add_generic_AC_RND_CONV_false_18_mux_1_itm_mx1c2 = or_dcpl_224 |
      return_add_generic_AC_RND_CONV_false_12_r_zero_or_1_cse | or_dcpl_702 | or_dcpl_943
      | or_dcpl_559 | (fsm_output[38]) | (fsm_output[12]) | (fsm_output[37]);
  assign not_tmp_376 = stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0 ^ stage_PE_1_tmp_re_d_1_lpi_3_dfm_63;
  assign not_tmp_395 = stage_PE_1_tmp_im_d_1_lpi_3_dfm_63_mx0 ^ stage_PE_1_tmp_re_d_1_lpi_3_dfm_63;
  assign BUTTERFLY_1_i_mux1h_1_nl = MUX1HOT_s_1_7_2(reg_BUTTERFLY_1_i_9_0_ftd, (~
      reg_BUTTERFLY_1_i_9_0_ftd), (BUTTERFLY_1_fry_9_0_sva[9]), (~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm),
      (~ (BUTTERFLY_i_9_0_sva_1[9])), (~ (BUTTERFLY_1_fry_9_0_sva[9])), (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[9]),
      {or_1174_ssc , (fsm_output[9]) , or_1176_ssc , or_1177_ssc , (fsm_output[28])
      , or_1179_ssc , (fsm_output[53])});
  assign or_2033_nl = or_1174_ssc | (fsm_output[9]) | or_1177_ssc;
  assign or_2009_nl = or_1179_ssc | or_1176_ssc;
  assign mux1h_6_nl = MUX1HOT_v_9_4_2(reg_BUTTERFLY_1_i_9_0_ftd_1, (BUTTERFLY_i_9_0_sva_1[8:0]),
      (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[8:0]),
      (BUTTERFLY_1_fry_9_0_sva[8:0]), {or_2033_nl , (fsm_output[28]) , (fsm_output[53])
      , or_2009_nl});
  assign in_f_d_rsci_adr_d = {BUTTERFLY_1_i_mux1h_1_nl , mux1h_6_nl};
  assign nor_175_m1c = ~(or_tmp_958 | or_tmp_959 | or_tmp_960);
  assign BUTTERFLY_if_1_if_and_7_cse = return_add_generic_AC_RND_CONV_false_10_or_1_svs_1
      & (fsm_output[22]);
  assign BUTTERFLY_if_1_if_and_9_cse = return_add_generic_AC_RND_CONV_false_12_or_1_svs_1
      & (fsm_output[26]);
  assign BUTTERFLY_if_1_if_and_6_cse = return_add_generic_AC_RND_CONV_false_9_or_1_svs_1
      & (fsm_output[20]);
  assign BUTTERFLY_if_1_if_and_8_cse = return_add_generic_AC_RND_CONV_false_11_or_1_svs_1
      & (fsm_output[24]);
  assign BUTTERFLY_if_1_if_and_5_cse = return_add_generic_AC_RND_CONV_false_or_1_svs_1
      & (fsm_output[8]);
  assign BUTTERFLY_if_1_if_or_2_cse = ((~ return_add_generic_AC_RND_CONV_false_or_1_svs_1)
      & (fsm_output[8])) | ((~ return_add_generic_AC_RND_CONV_false_9_or_1_svs_1)
      & (fsm_output[20])) | ((~ return_add_generic_AC_RND_CONV_false_10_or_1_svs_1)
      & (fsm_output[22])) | ((~ return_add_generic_AC_RND_CONV_false_11_or_1_svs_1)
      & (fsm_output[24])) | ((~ return_add_generic_AC_RND_CONV_false_12_or_1_svs_1)
      & (fsm_output[26]));
  assign and_339_cse = reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd
      & return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign BUTTERFLY_if_1_if_or_1_nl = (fsm_output[9]) | (fsm_output[22]);
  assign BUTTERFLY_if_1_if_mux1h_nl = MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_16_mux_itm,
      operator_11_true_return_24_sva, return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_17_mux_6_itm, return_add_generic_AC_RND_CONV_false_11_mux_itm,
      return_add_generic_AC_RND_CONV_false_12_mux_itm, {BUTTERFLY_if_1_if_or_cse
      , BUTTERFLY_if_1_if_or_1_nl , (fsm_output[16]) , (fsm_output[18]) , (fsm_output[24])
      , (fsm_output[26])});
  assign and_2629_nl = (fsm_output[8]) & nor_175_m1c;
  assign or_2745_nl = ((fsm_output[20]) & nor_175_m1c) | ((fsm_output[22]) & nor_175_m1c)
      | ((fsm_output[24]) & nor_175_m1c) | ((fsm_output[26]) & nor_175_m1c);
  assign mux1h_1_nl = MUX1HOT_v_10_6_2(return_add_generic_AC_RND_CONV_false_1_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0, return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1, (return_add_generic_AC_RND_CONV_false_9_exp_plus_1_12_1_lpi_3_dfm_1[9:0]),
      return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_11,
      {and_2629_nl , (fsm_output[9]) , (fsm_output[16]) , (fsm_output[18]) , or_2745_nl
      , or_tmp_959});
  assign not_1022_nl = ~ or_tmp_960;
  assign and_2637_nl = MUX_v_10_2_2(10'b0000000000, mux1h_1_nl, not_1022_nl);
  assign or_2027_nl = MUX_v_10_2_2(and_2637_nl, 10'b1111111111, or_tmp_958);
  assign or_358_nl = and_281_cse | operator_11_true_return_1_sva | or_dcpl_285;
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_2_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs, or_358_nl);
  assign return_add_generic_AC_RND_CONV_false_e_r_return_add_generic_AC_RND_CONV_false_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_30 & (~ return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_2_nl))
      | return_add_generic_AC_RND_CONV_false_exception_sva_1;
  assign or_467_nl = and_340_cse | operator_11_true_return_1_sva | or_dcpl_367 |
      and_339_cse;
  assign return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs, or_467_nl);
  assign return_add_generic_AC_RND_CONV_false_9_e_r_return_add_generic_AC_RND_CONV_false_9_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_30 & (~ return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_nl))
      | return_add_generic_AC_RND_CONV_false_9_exception_sva_1;
  assign or_476_nl = and_348_cse | operator_11_true_return_21_sva | operator_11_true_return_22_sva
      | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva | and_339_cse;
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_7_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs, or_476_nl);
  assign return_add_generic_AC_RND_CONV_false_10_e_r_return_add_generic_AC_RND_CONV_false_10_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_30 & (~ return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_7_nl))
      | return_add_generic_AC_RND_CONV_false_10_exception_sva_1;
  assign or_483_nl = and_356_cse | or_dcpl_93 | or_dcpl_367 | and_339_cse;
  assign return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_2_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs, or_483_nl);
  assign return_add_generic_AC_RND_CONV_false_11_e_r_return_add_generic_AC_RND_CONV_false_11_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_30 & (~ return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_2_nl))
      | return_add_generic_AC_RND_CONV_false_11_exception_sva_1;
  assign or_490_nl = and_362_cse | or_dcpl_311 | or_dcpl_359 | and_339_cse;
  assign return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_3_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs, or_490_nl);
  assign return_add_generic_AC_RND_CONV_false_12_e_r_return_add_generic_AC_RND_CONV_false_12_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_30 & (~ return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_3_nl))
      | return_add_generic_AC_RND_CONV_false_12_exception_sva_1;
  assign BUTTERFLY_if_1_if_mux1h_2_nl = MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_e_r_return_add_generic_AC_RND_CONV_false_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm,
      return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_9_e_r_return_add_generic_AC_RND_CONV_false_9_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_10_e_r_return_add_generic_AC_RND_CONV_false_10_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_11_e_r_return_add_generic_AC_RND_CONV_false_11_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_12_e_r_return_add_generic_AC_RND_CONV_false_12_e_r_or_1_nl,
      {(fsm_output[8]) , (fsm_output[9]) , (fsm_output[16]) , (fsm_output[18]) ,
      (fsm_output[20]) , (fsm_output[22]) , (fsm_output[24]) , (fsm_output[26])});
  assign return_add_generic_AC_RND_CONV_false_9_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0 | (return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0 & return_add_generic_AC_RND_CONV_false_18_mux_itm);
  assign return_add_generic_AC_RND_CONV_false_10_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_mx2w0 | (operator_11_true_return_22_sva
      & return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0 & return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_11_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_unequal_tmp | return_add_generic_AC_RND_CONV_false_11_do_sub_sva;
  assign return_add_generic_AC_RND_CONV_false_12_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | operator_11_true_return_1_sva;
  assign BUTTERFLY_if_1_if_or_3_nl = BUTTERFLY_if_1_if_and_5_cse | ((~ and_2472_tmp)
      & (fsm_output[16]));
  assign BUTTERFLY_if_1_if_and_11_nl = and_2472_tmp & (fsm_output[16]);
  assign BUTTERFLY_if_1_if_mux1h_3_nl = MUX1HOT_s_1_9_2(return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_r_nan_or_cse, drf_qr_lval_14_smx_0_lpi_3_dfm,
      (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1[51]), return_add_generic_AC_RND_CONV_false_8_m_r_51_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_9_r_nan_or_nl, return_add_generic_AC_RND_CONV_false_10_r_nan_or_nl,
      return_add_generic_AC_RND_CONV_false_11_r_nan_or_nl, return_add_generic_AC_RND_CONV_false_12_r_nan_or_nl,
      {BUTTERFLY_if_1_if_or_2_cse , BUTTERFLY_if_1_if_or_3_nl , (fsm_output[9]) ,
      BUTTERFLY_if_1_if_and_11_nl , (fsm_output[18]) , BUTTERFLY_if_1_if_and_6_cse
      , BUTTERFLY_if_1_if_and_7_cse , BUTTERFLY_if_1_if_and_8_cse , BUTTERFLY_if_1_if_and_9_cse});
  assign mux1h_2_nl = MUX1HOT_v_51_4_2(return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm,
      return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm,
      {(fsm_output[9]) , (fsm_output[16]) , (fsm_output[18]) , BUTTERFLY_if_1_if_or_2_cse});
  assign nor_246_nl = ~(BUTTERFLY_if_1_if_and_7_cse | BUTTERFLY_if_1_if_and_9_cse
      | BUTTERFLY_if_1_if_and_6_cse | BUTTERFLY_if_1_if_and_8_cse | BUTTERFLY_if_1_if_and_5_cse);
  assign and_3934_nl = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      mux1h_2_nl, nor_246_nl);
  assign in_f_d_rsci_d_d = {BUTTERFLY_if_1_if_mux1h_nl , or_2027_nl , BUTTERFLY_if_1_if_mux1h_2_nl
      , BUTTERFLY_if_1_if_mux1h_3_nl , and_3934_nl};
  assign in_f_d_rsci_we_d_pff = (stage_PE_1_and_1_tmp & ((fsm_output[18]) | (fsm_output[16])
      | or_dcpl_269)) | (and_dcpl_18 & (or_dcpl_273 | or_dcpl_272));
  assign in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = (mode_lpi_1_dfm & ((fsm_output[28])
      | (fsm_output[31]))) | (and_dcpl_18 & or_dcpl_221) | (stage_PE_1_and_1_tmp
      & or_dcpl_201) | and_741_cse;
  assign BUTTERFLY_1_i_or_3_cse = (inverse_lpi_1_dfm_1 & (fsm_output[28])) | ((~
      inverse_lpi_1_dfm_1) & (fsm_output[28]));
  assign BUTTERFLY_1_i_mux1h_nl = MUX1HOT_s_1_4_2(reg_BUTTERFLY_1_i_9_0_ftd, (BUTTERFLY_1_fry_9_0_sva[9]),
      (z_out_67[9]), (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[9]),
      {or_1159_ssc , or_1160_ssc , BUTTERFLY_1_i_or_3_cse , or_dcpl_207});
  assign BUTTERFLY_1_i_mux1h_6_nl = MUX1HOT_v_9_4_2(reg_BUTTERFLY_1_i_9_0_ftd_1,
      (BUTTERFLY_1_fry_9_0_sva[8:0]), (z_out_67[8:0]), (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[8:0]),
      {or_1159_ssc , or_1160_ssc , BUTTERFLY_1_i_or_3_cse , or_dcpl_207});
  assign in_u_rsci_adr_d = {BUTTERFLY_1_i_mux1h_nl , BUTTERFLY_1_i_mux1h_6_nl};
  assign BUTTERFLY_else_1_if_or_nl = (fsm_output[6]) | return_add_generic_AC_RND_CONV_false_11_and_10_cse;
  assign in_u_rsci_d_d = MUX1HOT_v_16_4_2(z_out_59, (z_out_111[15:0]), ({BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0
      , BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0 , BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1}),
      ({{1{stage_monty_mul_acc_2_psp_sva_1[14]}}, stage_monty_mul_acc_2_psp_sva_1}),
      {BUTTERFLY_else_1_if_or_nl , and_746_cse , (fsm_output[8]) , (fsm_output[54])});
  assign in_u_rsci_we_d_pff = ((~ mode_lpi_1_dfm) & (fsm_output[7])) | and_630_cse
      | and_662_cse | (and_dcpl_185 & (fsm_output[8]));
  assign in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = and_741_cse | (~(mode_lpi_1_dfm
      | (~((fsm_output[28]) | (fsm_output[30])))));
  assign BUTTERFLY_if_1_mux1h_2_nl = MUX1HOT_s_1_7_2((~ (BUTTERFLY_i_9_0_sva_1[9])),
      (~ (BUTTERFLY_1_fry_9_0_sva[9])), (BUTTERFLY_1_fry_9_0_sva[9]), reg_BUTTERFLY_1_i_9_0_ftd,
      (~ reg_BUTTERFLY_1_i_9_0_ftd), (~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm),
      (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[9]),
      {(fsm_output[3]) , or_1146_ssc , or_1147_ssc , or_1148_ssc , (fsm_output[34])
      , or_1150_ssc , (fsm_output[53])});
  assign or_2034_nl = or_1148_ssc | (fsm_output[34]) | or_1150_ssc;
  assign or_2010_nl = or_1147_ssc | or_1146_ssc;
  assign mux1h_7_nl = MUX1HOT_v_9_4_2((BUTTERFLY_i_9_0_sva_1[8:0]), reg_BUTTERFLY_1_i_9_0_ftd_1,
      (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[8:0]),
      (BUTTERFLY_1_fry_9_0_sva[8:0]), {(fsm_output[3]) , or_2034_nl , (fsm_output[53])
      , or_2010_nl});
  assign out_f_d_rsci_adr_d = {BUTTERFLY_if_1_mux1h_2_nl , mux1h_7_nl};
  assign nor_177_m1c = ~(or_tmp_963 | or_tmp_964 | or_tmp_965);
  assign BUTTERFLY_if_1_and_9_cse = return_add_generic_AC_RND_CONV_false_23_or_1_svs_1
      & (fsm_output[47]);
  assign BUTTERFLY_if_1_and_11_cse = return_add_generic_AC_RND_CONV_false_25_or_1_svs_1
      & (fsm_output[51]);
  assign BUTTERFLY_if_1_and_8_cse = return_add_generic_AC_RND_CONV_false_22_or_1_svs_1
      & (fsm_output[45]);
  assign BUTTERFLY_if_1_and_10_cse = return_add_generic_AC_RND_CONV_false_24_or_1_svs_1
      & (fsm_output[49]);
  assign BUTTERFLY_if_1_and_7_cse = return_add_generic_AC_RND_CONV_false_13_or_1_svs_1
      & (fsm_output[33]);
  assign BUTTERFLY_if_1_or_2_cse = ((~ return_add_generic_AC_RND_CONV_false_13_or_1_svs_1)
      & (fsm_output[33])) | ((~ return_add_generic_AC_RND_CONV_false_22_or_1_svs_1)
      & (fsm_output[45])) | ((~ return_add_generic_AC_RND_CONV_false_23_or_1_svs_1)
      & (fsm_output[47])) | ((~ return_add_generic_AC_RND_CONV_false_24_or_1_svs_1)
      & (fsm_output[49])) | ((~ return_add_generic_AC_RND_CONV_false_25_or_1_svs_1)
      & (fsm_output[51]));
  assign BUTTERFLY_if_1_or_nl = (fsm_output[33]) | (fsm_output[45]);
  assign BUTTERFLY_if_1_or_1_nl = (fsm_output[34]) | (fsm_output[47]);
  assign BUTTERFLY_if_1_mux1h_1_nl = MUX1HOT_s_1_6_2(operator_11_true_return_24_sva,
      return_add_generic_AC_RND_CONV_false_11_mux_itm, return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_17_mux_6_itm, return_add_generic_AC_RND_CONV_false_12_mux_itm,
      return_add_generic_AC_RND_CONV_false_16_mux_itm, {BUTTERFLY_if_1_or_nl , BUTTERFLY_if_1_or_1_nl
      , (fsm_output[41]) , (fsm_output[43]) , (fsm_output[49]) , (fsm_output[51])});
  assign or_2746_nl = ((fsm_output[33]) & nor_177_m1c) | ((fsm_output[45]) & nor_177_m1c)
      | ((fsm_output[47]) & nor_177_m1c) | ((fsm_output[49]) & nor_177_m1c) | ((fsm_output[51])
      & nor_177_m1c);
  assign mux1h_3_nl = MUX1HOT_v_10_5_2((return_add_generic_AC_RND_CONV_false_9_exp_plus_1_12_1_lpi_3_dfm_1[9:0]),
      return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0, return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_11,
      {or_2746_nl , (fsm_output[34]) , (fsm_output[41]) , (fsm_output[43]) , or_tmp_963});
  assign not_1025_nl = ~ or_tmp_964;
  assign and_2654_nl = MUX_v_10_2_2(10'b0000000000, mux1h_3_nl, not_1025_nl);
  assign or_2028_nl = MUX_v_10_2_2(and_2654_nl, 10'b1111111111, or_tmp_965);
  assign or_416_nl = and_317_cse | operator_11_true_return_1_sva | and_339_cse |
      operator_11_true_return_21_sva;
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_5_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs, or_416_nl);
  assign return_add_generic_AC_RND_CONV_false_13_e_r_return_add_generic_AC_RND_CONV_false_13_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_30 & (~ return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_5_nl))
      | return_add_generic_AC_RND_CONV_false_13_exception_sva_1;
  assign or_498_nl = and_368_cse | operator_11_true_return_1_sva | return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva | and_339_cse;
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_8_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs, or_498_nl);
  assign return_add_generic_AC_RND_CONV_false_22_e_r_return_add_generic_AC_RND_CONV_false_22_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_30 & (~ return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_8_nl))
      | return_add_generic_AC_RND_CONV_false_22_exception_sva_1;
  assign or_506_nl = and_374_cse | operator_11_true_return_21_sva | or_dcpl_438 |
      and_339_cse;
  assign return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_4_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs, or_506_nl);
  assign return_add_generic_AC_RND_CONV_false_23_e_r_return_add_generic_AC_RND_CONV_false_23_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_30 & (~ return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_4_nl))
      | return_add_generic_AC_RND_CONV_false_23_exception_sva_1;
  assign or_514_nl = and_382_cse | return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | or_dcpl_359 | and_339_cse;
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_9_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs, or_514_nl);
  assign return_add_generic_AC_RND_CONV_false_24_e_r_return_add_generic_AC_RND_CONV_false_24_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_30 & (~ return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_9_nl))
      | return_add_generic_AC_RND_CONV_false_24_exception_sva_1;
  assign or_521_nl = and_389_cse | or_dcpl_93 | or_dcpl_438 | and_339_cse;
  assign return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_3_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs, or_521_nl);
  assign return_add_generic_AC_RND_CONV_false_25_e_r_return_add_generic_AC_RND_CONV_false_25_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_30 & (~ return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_3_nl))
      | return_add_generic_AC_RND_CONV_false_25_exception_sva_1;
  assign BUTTERFLY_if_1_mux1h_6_nl = MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_13_e_r_return_add_generic_AC_RND_CONV_false_13_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm,
      return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_22_e_r_return_add_generic_AC_RND_CONV_false_22_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_23_e_r_return_add_generic_AC_RND_CONV_false_23_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_24_e_r_return_add_generic_AC_RND_CONV_false_24_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_25_e_r_return_add_generic_AC_RND_CONV_false_25_e_r_or_1_nl,
      {(fsm_output[33]) , (fsm_output[34]) , (fsm_output[41]) , (fsm_output[43])
      , (fsm_output[45]) , (fsm_output[47]) , (fsm_output[49]) , (fsm_output[51])});
  assign return_add_generic_AC_RND_CONV_false_22_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_23_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | (operator_11_true_return_22_sva
      & return_mult_generic_AC_RND_CONV_false_1_op1_zero_sva_1 & return_add_generic_AC_RND_CONV_false_18_mux_itm);
  assign return_add_generic_AC_RND_CONV_false_24_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_11_do_sub_sva;
  assign return_add_generic_AC_RND_CONV_false_25_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_unequal_tmp | operator_11_true_return_1_sva;
  assign BUTTERFLY_if_1_mux1h_7_nl = MUX1HOT_s_1_9_2(return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_r_nan_or_cse, drf_qr_lval_14_smx_0_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_21_m_r_51_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_22_r_nan_or_nl, return_add_generic_AC_RND_CONV_false_23_r_nan_or_nl,
      return_add_generic_AC_RND_CONV_false_24_r_nan_or_nl, return_add_generic_AC_RND_CONV_false_25_r_nan_or_nl,
      {BUTTERFLY_if_1_or_2_cse , BUTTERFLY_if_1_and_7_cse , (fsm_output[34]) , (fsm_output[41])
      , (fsm_output[43]) , BUTTERFLY_if_1_and_8_cse , BUTTERFLY_if_1_and_9_cse ,
      BUTTERFLY_if_1_and_10_cse , BUTTERFLY_if_1_and_11_cse});
  assign mux1h_4_nl = MUX1HOT_v_51_4_2(return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm,
      return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm,
      {(fsm_output[34]) , (fsm_output[41]) , (fsm_output[43]) , BUTTERFLY_if_1_or_2_cse});
  assign nor_247_nl = ~(BUTTERFLY_if_1_and_9_cse | BUTTERFLY_if_1_and_11_cse | BUTTERFLY_if_1_and_8_cse
      | BUTTERFLY_if_1_and_10_cse | BUTTERFLY_if_1_and_7_cse);
  assign and_3935_nl = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      mux1h_4_nl, nor_247_nl);
  assign out_f_d_rsci_d_d = {BUTTERFLY_if_1_mux1h_1_nl , or_2028_nl , BUTTERFLY_if_1_mux1h_6_nl
      , BUTTERFLY_if_1_mux1h_7_nl , and_3935_nl};
  assign out_f_d_rsci_we_d_pff = (and_dcpl_18 & ((fsm_output[51]) | (fsm_output[45])
      | or_dcpl_253)) | (stage_PE_1_and_1_tmp & (or_dcpl_223 | (fsm_output[34:33]!=2'b00)));
  assign out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = (mode_lpi_1_dfm & ((fsm_output[3])
      | (fsm_output[6]))) | (or_dcpl_227 & (fsm_output[53])) | (stage_PE_1_and_1_tmp
      & or_dcpl_200) | (and_dcpl_18 & or_dcpl_245);
  assign BUTTERFLY_else_1_or_cse = (inverse_lpi_1_dfm_1 & (fsm_output[3])) | ((~
      inverse_lpi_1_dfm_1) & (fsm_output[3]));
  assign BUTTERFLY_else_1_mux1h_nl = MUX1HOT_s_1_4_2((z_out_67[9]), reg_BUTTERFLY_1_i_9_0_ftd,
      (BUTTERFLY_1_fry_9_0_sva[9]), (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[9]),
      {BUTTERFLY_else_1_or_cse , or_1132_ssc , or_1133_ssc , (fsm_output[53])});
  assign BUTTERFLY_else_1_mux1h_1_nl = MUX1HOT_v_9_4_2((z_out_67[8:0]), reg_BUTTERFLY_1_i_9_0_ftd_1,
      (BUTTERFLY_1_fry_9_0_sva[8:0]), (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[8:0]),
      {BUTTERFLY_else_1_or_cse , or_1132_ssc , or_1133_ssc , (fsm_output[53])});
  assign out_u_rsci_adr_d = {BUTTERFLY_else_1_mux1h_nl , BUTTERFLY_else_1_mux1h_1_nl};
  assign BUTTERFLY_else_1_if_or_1_nl = (fsm_output[31]) | return_add_generic_AC_RND_CONV_false_12_and_112_cse;
  assign out_u_rsci_d_d = MUX1HOT_v_16_3_2(z_out_59, (z_out_111[15:0]), ({BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0
      , BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0 , BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1}),
      {BUTTERFLY_else_1_if_or_1_nl , and_680_cse , (fsm_output[33])});
  assign out_u_rsci_we_d_pff = and_647_cse | (and_dcpl_185 & (fsm_output[33])) |
      ((~ mode_lpi_1_dfm) & (fsm_output[32]));
  assign out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = (~(mode_lpi_1_dfm | (~((fsm_output[3])
      | (fsm_output[5]))))) | (operator_16_false_operator_16_false_nor_cse_sva &
      (fsm_output[53]));
  assign BUTTERFLY_1_else_nand_tmp = ~((~((fsm_output[3]) | (fsm_output[28]))) &
      (~((fsm_output[55]) | (fsm_output[42]))) & and_dcpl_360 & (~ (fsm_output[23]))
      & (~((fsm_output[22]) | (fsm_output[20]))) & (~((fsm_output[21]) | (fsm_output[43])))
      & and_dcpl_354 & (~ (fsm_output[41])) & (~((fsm_output[16]) | (fsm_output[34])))
      & (~((fsm_output[7]) | (fsm_output[9]))) & (~((fsm_output[35]) | (fsm_output[10])
      | (fsm_output[54]))) & and_dcpl_344 & (~ (fsm_output[33])) & (~((fsm_output[6])
      | (fsm_output[32]) | (fsm_output[31]))));
  assign and_dcpl_564 = BUTTERFLY_1_else_nand_tmp & (~ return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs_mx0w0);
  assign or_tmp = ((~ return_add_generic_AC_RND_CONV_false_14_exception_sva_1) &
      (fsm_output[31])) | ((~ return_add_generic_AC_RND_CONV_false_1_exception_sva_1)
      & (fsm_output[6]));
  assign or_tmp_954 = (return_add_generic_AC_RND_CONV_false_14_exception_sva_1 &
      (fsm_output[31])) | (return_add_generic_AC_RND_CONV_false_16_exception_sva_1
      & (fsm_output[35])) | (return_add_generic_AC_RND_CONV_false_2_exception_sva_1
      & (fsm_output[9])) | (return_add_generic_AC_RND_CONV_false_1_exception_sva_1
      & (fsm_output[6])) | (return_add_generic_AC_RND_CONV_false_3_exception_sva_1
      & (fsm_output[10])) | (return_add_generic_AC_RND_CONV_false_15_exception_sva_1
      & (fsm_output[34]));
  assign or_tmp_955 = ~(BUTTERFLY_1_else_nand_tmp & (~(return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs_mx0w0
      & (~ return_add_generic_AC_RND_CONV_false_16_exception_sva_1) & (fsm_output[35])))
      & (~((~((~ return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0) |
      return_add_generic_AC_RND_CONV_false_2_exception_sva_1)) & (fsm_output[9])))
      & (~(return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs_mx0w0 & (~ return_add_generic_AC_RND_CONV_false_3_exception_sva_1)
      & (fsm_output[10]))) & (~((~((~ return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs_mx0w0)
      | return_add_generic_AC_RND_CONV_false_15_exception_sva_1)) & (fsm_output[34]))));
  assign or_tmp_956 = (and_dcpl_564 & (~((z_out_89[53]) | return_add_generic_AC_RND_CONV_false_16_exception_sva_1))
      & (fsm_output[35])) | (and_dcpl_564 & (~((z_out_89[53]) | return_add_generic_AC_RND_CONV_false_3_exception_sva_1))
      & (fsm_output[10]));
  assign or_tmp_958 = (return_add_generic_AC_RND_CONV_false_10_exception_sva_1 &
      (fsm_output[22])) | (return_add_generic_AC_RND_CONV_false_12_exception_sva_1
      & (fsm_output[26])) | (return_add_generic_AC_RND_CONV_false_9_exception_sva_1
      & (fsm_output[20])) | (return_add_generic_AC_RND_CONV_false_11_exception_sva_1
      & (fsm_output[24])) | (return_add_generic_AC_RND_CONV_false_exception_sva_1
      & (fsm_output[8]));
  assign or_tmp_959 = ((~(return_add_generic_AC_RND_CONV_false_10_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1))
      & (fsm_output[22])) | ((~(return_add_generic_AC_RND_CONV_false_12_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1))
      & (fsm_output[26])) | ((~(return_add_generic_AC_RND_CONV_false_9_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w1))
      & (fsm_output[20])) | ((~(return_add_generic_AC_RND_CONV_false_11_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w1))
      & (fsm_output[24]));
  assign or_tmp_960 = ((~ return_add_generic_AC_RND_CONV_false_10_exception_sva_1)
      & return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1 & (fsm_output[22]))
      | ((~ return_add_generic_AC_RND_CONV_false_12_exception_sva_1) & return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1
      & (fsm_output[26])) | ((~ return_add_generic_AC_RND_CONV_false_9_exception_sva_1)
      & return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w1 & (fsm_output[20]))
      | ((~ return_add_generic_AC_RND_CONV_false_11_exception_sva_1) & return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w1
      & (fsm_output[24]));
  assign or_tmp_963 = ((~(return_add_generic_AC_RND_CONV_false_23_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1))
      & (fsm_output[47])) | ((~(return_add_generic_AC_RND_CONV_false_25_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w1))
      & (fsm_output[51])) | ((~(return_add_generic_AC_RND_CONV_false_22_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1))
      & (fsm_output[45])) | ((~(return_add_generic_AC_RND_CONV_false_24_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1))
      & (fsm_output[49])) | ((~(return_add_generic_AC_RND_CONV_false_13_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1))
      & (fsm_output[33]));
  assign or_tmp_964 = ((~ return_add_generic_AC_RND_CONV_false_23_exception_sva_1)
      & return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1 & (fsm_output[47]))
      | ((~ return_add_generic_AC_RND_CONV_false_25_exception_sva_1) & return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w1
      & (fsm_output[51])) | ((~ return_add_generic_AC_RND_CONV_false_22_exception_sva_1)
      & return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1 & (fsm_output[45]))
      | ((~ return_add_generic_AC_RND_CONV_false_24_exception_sva_1) & return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1
      & (fsm_output[49])) | ((~ return_add_generic_AC_RND_CONV_false_13_exception_sva_1)
      & return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1 & (fsm_output[33]));
  assign or_tmp_965 = (return_add_generic_AC_RND_CONV_false_23_exception_sva_1 &
      (fsm_output[47])) | (return_add_generic_AC_RND_CONV_false_25_exception_sva_1
      & (fsm_output[51])) | (return_add_generic_AC_RND_CONV_false_22_exception_sva_1
      & (fsm_output[45])) | (return_add_generic_AC_RND_CONV_false_24_exception_sva_1
      & (fsm_output[49])) | (return_add_generic_AC_RND_CONV_false_13_exception_sva_1
      & (fsm_output[33]));
  assign and_3379_cse = inverse_lpi_1_dfm_1 & or_dcpl_198;
  assign or_2455_cse = (fsm_output[38]) | (fsm_output[11]) | (fsm_output[36]) | (fsm_output[13]);
  assign or_tmp_1400 = (fsm_output[45]) | (fsm_output[20]);
  assign or_tmp_1439 = (fsm_output[40]) | (fsm_output[15]) | (fsm_output[34]);
  assign or_tmp_1440 = (fsm_output[42]) | (fsm_output[17]) | (fsm_output[9]);
  assign or_tmp_1491 = (fsm_output[41]) | (fsm_output[31]) | (fsm_output[8]) | (fsm_output[16])
      | (fsm_output[6]) | (fsm_output[34]);
  assign or_tmp_1492 = (fsm_output[33]) | (fsm_output[9]);
  assign or_1342_itm = or_dcpl_504 | return_add_generic_AC_RND_CONV_false_11_or_4_cse
      | return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse | or_dcpl_497 |
      or_dcpl_493 | or_dcpl_492;
  assign return_add_generic_AC_RND_CONV_false_7_exp_and_ssc = run_wen & ((~(and_dcpl_467
      | or_dcpl_511 | (fsm_output[40]) | (fsm_output[33]))) | (fsm_output[5]) | (fsm_output[7])
      | or_dcpl_208 | (fsm_output[14:13]!=2'b00) | or_dcpl_521 | or_dcpl_673 | or_dcpl_671
      | or_dcpl_473 | (fsm_output[18]) | (fsm_output[30]) | (fsm_output[32]) | or_dcpl_235
      | (fsm_output[37]));
  assign return_add_generic_AC_RND_CONV_false_12_res_mant_and_1_ssc = return_add_generic_AC_RND_CONV_false_12_res_mant_and_ssc
      & (~ or_dcpl_845);
  assign return_add_generic_AC_RND_CONV_false_9_mux_28_cse = MUX_v_56_2_2((z_out_74[56:1]),
      (~ (z_out_74[56:1])), return_add_generic_AC_RND_CONV_false_18_mux_itm);
  assign return_add_generic_AC_RND_CONV_false_6_res_mant_conc_2_itm_56_1 = MUX_v_56_2_2((~
      (z_out_73[56:1])), (z_out_73[56:1]), not_tmp_376);
  assign return_add_generic_AC_RND_CONV_false_7_mux_31_cse = MUX_v_56_2_2((z_out_75[56:1]),
      (~ (z_out_75[56:1])), return_add_generic_AC_RND_CONV_false_20_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_10_mux_28_cse = MUX_v_56_2_2((z_out_74[56:1]),
      (~ (z_out_74[56:1])), return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_19_res_mant_conc_2_itm_56_1 = MUX_v_56_2_2((~
      (z_out_74[56:1])), (z_out_74[56:1]), not_tmp_395);
  assign return_mult_generic_AC_RND_CONV_false_return_mult_generic_AC_RND_CONV_false_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_if_1_and_1_tmp_1 | (operator_14_false_1_acc_psp_sva_12_10[2]));
  assign return_mult_generic_AC_RND_CONV_false_1_return_mult_generic_AC_RND_CONV_false_1_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_tmp_1 | (operator_14_false_1_acc_psp_sva_12_10[2]));
  assign return_mult_generic_AC_RND_CONV_false_2_return_mult_generic_AC_RND_CONV_false_2_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_2_if_1_and_1_tmp_1 | (operator_14_false_1_acc_psp_sva_12_10[2]));
  assign return_mult_generic_AC_RND_CONV_false_3_return_mult_generic_AC_RND_CONV_false_3_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_3_if_1_and_1_tmp_1 | (operator_14_false_1_acc_psp_sva_12_10[2]));
  assign return_mult_generic_AC_RND_CONV_false_4_return_mult_generic_AC_RND_CONV_false_4_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_4_if_1_and_1_tmp_1 | (operator_14_false_1_acc_psp_sva_12_10[2]));
  assign return_mult_generic_AC_RND_CONV_false_5_return_mult_generic_AC_RND_CONV_false_5_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_5_if_1_and_1_tmp_1 | (operator_14_false_1_acc_psp_sva_12_10[2]));
  assign return_mult_generic_AC_RND_CONV_false_mux1h_cse = MUX1HOT_s_1_6_2(return_mult_generic_AC_RND_CONV_false_return_mult_generic_AC_RND_CONV_false_nor_nl,
      return_mult_generic_AC_RND_CONV_false_1_return_mult_generic_AC_RND_CONV_false_1_nor_nl,
      return_mult_generic_AC_RND_CONV_false_2_return_mult_generic_AC_RND_CONV_false_2_nor_nl,
      return_mult_generic_AC_RND_CONV_false_3_return_mult_generic_AC_RND_CONV_false_3_nor_nl,
      return_mult_generic_AC_RND_CONV_false_4_return_mult_generic_AC_RND_CONV_false_4_nor_nl,
      return_mult_generic_AC_RND_CONV_false_5_return_mult_generic_AC_RND_CONV_false_5_nor_nl,
      {(fsm_output[12]) , (fsm_output[13]) , (fsm_output[14]) , (fsm_output[37])
      , (fsm_output[38]) , (fsm_output[39])});
  assign return_mult_generic_AC_RND_CONV_false_and_2_nl = return_mult_generic_AC_RND_CONV_false_if_1_and_1_tmp_1
      & (~ (operator_14_false_1_acc_psp_sva_12_10[2]));
  assign return_mult_generic_AC_RND_CONV_false_1_and_2_nl = return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_tmp_1
      & (~ (operator_14_false_1_acc_psp_sva_12_10[2]));
  assign return_mult_generic_AC_RND_CONV_false_2_and_2_nl = return_mult_generic_AC_RND_CONV_false_2_if_1_and_1_tmp_1
      & (~ (operator_14_false_1_acc_psp_sva_12_10[2]));
  assign return_mult_generic_AC_RND_CONV_false_3_and_2_nl = return_mult_generic_AC_RND_CONV_false_3_if_1_and_1_tmp_1
      & (~ (operator_14_false_1_acc_psp_sva_12_10[2]));
  assign return_mult_generic_AC_RND_CONV_false_4_and_2_nl = return_mult_generic_AC_RND_CONV_false_4_if_1_and_1_tmp_1
      & (~ (operator_14_false_1_acc_psp_sva_12_10[2]));
  assign return_mult_generic_AC_RND_CONV_false_5_and_2_nl = return_mult_generic_AC_RND_CONV_false_5_if_1_and_1_tmp_1
      & (~ (operator_14_false_1_acc_psp_sva_12_10[2]));
  assign return_mult_generic_AC_RND_CONV_false_mux1h_1_cse = MUX1HOT_s_1_6_2(return_mult_generic_AC_RND_CONV_false_and_2_nl,
      return_mult_generic_AC_RND_CONV_false_1_and_2_nl, return_mult_generic_AC_RND_CONV_false_2_and_2_nl,
      return_mult_generic_AC_RND_CONV_false_3_and_2_nl, return_mult_generic_AC_RND_CONV_false_4_and_2_nl,
      return_mult_generic_AC_RND_CONV_false_5_and_2_nl, {(fsm_output[12]) , (fsm_output[13])
      , (fsm_output[14]) , (fsm_output[37]) , (fsm_output[38]) , (fsm_output[39])});
  assign return_add_generic_AC_RND_CONV_false_e_dif1_or_1_cse = return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse
      | (fsm_output[32]) | (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_12_or_9_cse = BUTTERFLY_else_or_cse
      | or_tmp_1400 | or_dcpl_553 | or_dcpl_493;
  assign return_add_generic_AC_RND_CONV_false_12_or_11_cse_1 = (fsm_output[16]) |
      (fsm_output[43]);
  assign operator_6_false_33_or_5_cse = (fsm_output[19]) | (fsm_output[48]);
  assign operator_6_false_33_or_7_cse = (fsm_output[21]) | (fsm_output[50]);
  assign operator_6_false_33_or_1_cse = (fsm_output[23]) | (fsm_output[44]);
  assign operator_6_false_33_or_3_cse = (fsm_output[25]) | (fsm_output[46]);
  assign operator_6_false_3_or_1_ssc = or_tmp_1492 | or_dcpl_625;
  assign operator_6_false_3_or_6_cse = (fsm_output[20]) | (fsm_output[49]);
  assign operator_6_false_3_or_8_cse = (fsm_output[22]) | (fsm_output[51]);
  assign operator_6_false_3_or_2_cse = (fsm_output[24]) | (fsm_output[45]);
  assign operator_6_false_3_or_4_cse = (fsm_output[26]) | (fsm_output[47]);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif1_or_1_cse = (fsm_output[18])
      | return_add_generic_AC_RND_CONV_false_11_or_5_cse;
  assign return_add_generic_AC_RND_CONV_false_1_res_rounded_or_2_cse = (fsm_output[15])
      | (fsm_output[17]) | (fsm_output[19]) | (fsm_output[40]) | (fsm_output[42]);
  assign return_add_generic_AC_RND_CONV_false_7_res_rounded_and_cse = (z_out_79[3])
      & ((z_out_79[0]) | (z_out_79[1]) | (z_out_79[2]) | (z_out_79[4]));
  assign return_add_generic_AC_RND_CONV_false_7_mux_33_cse = MUX_v_6_2_2(return_add_generic_AC_RND_CONV_false_7_e_dif_sat_sva_1,
      return_add_generic_AC_RND_CONV_false_8_e_dif_sat_sva_1, fsm_output[39]);
  assign BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_4_cse = MUX_s_1_2_2((operator_32_false_3_acc_psp_sva_1[17]),
      (z_out_98[17]), BUTTERFLY_else_or_cse);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_or_cse = return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse
      | (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_12_or_22_cse = or_dcpl_534 | operator_6_false_17_or_cse;
  assign operator_6_false_33_or_12_cse = or_tmp_1439 | or_tmp_1440;
  assign operator_6_false_33_or_14_cse = (fsm_output[21]) | (fsm_output[48]);
  assign operator_6_false_33_or_15_cse = (fsm_output[23]) | (fsm_output[46]);
  assign operator_6_false_3_or_12_cse = (fsm_output[26]) | (fsm_output[51]);
  assign return_add_generic_AC_RND_CONV_false_12_or_41_cse = or_dcpl_534 | return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse;
  assign return_add_generic_AC_RND_CONV_false_3_or_4_cse = (fsm_output[5]) | (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_2_and_cse = (~ return_add_generic_AC_RND_CONV_false_9_acc_2_itm_11_1)
      & (fsm_output[19]);
  assign return_add_generic_AC_RND_CONV_false_2_and_6_cse = (~ return_add_generic_AC_RND_CONV_false_22_acc_2_itm_11_1)
      & (fsm_output[44]);
  assign return_add_generic_AC_RND_CONV_false_2_and_1_cse = return_add_generic_AC_RND_CONV_false_9_acc_2_itm_11_1
      & (fsm_output[19]);
  assign return_add_generic_AC_RND_CONV_false_2_and_2_cse = (~ return_add_generic_AC_RND_CONV_false_10_acc_2_itm_11_1)
      & (fsm_output[21]);
  assign return_add_generic_AC_RND_CONV_false_2_and_8_cse = (~ return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1)
      & (fsm_output[46]);
  assign return_add_generic_AC_RND_CONV_false_2_or_5_cse = (return_add_generic_AC_RND_CONV_false_10_acc_2_itm_11_1
      & (fsm_output[21])) | (return_add_generic_AC_RND_CONV_false_22_acc_2_itm_11_1
      & (fsm_output[44])) | (return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11_1
      & (fsm_output[48]));
  assign return_add_generic_AC_RND_CONV_false_2_and_4_cse = (~ return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1)
      & (fsm_output[23]);
  assign return_add_generic_AC_RND_CONV_false_2_and_10_cse = (~ return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11_1)
      & (fsm_output[48]);
  assign return_add_generic_AC_RND_CONV_false_2_or_7_cse = (return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1
      & (fsm_output[23])) | (return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1
      & (fsm_output[46]));
  assign return_add_generic_AC_RND_CONV_false_1_and_16_cse = (~ return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse)
      & (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_1_and_20_cse = (~ return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse)
      & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_1_or_7_cse = (return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse
      & (fsm_output[5])) | ((~ return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse)
      & (fsm_output[7]));
  assign return_add_generic_AC_RND_CONV_false_1_or_9_cse = (return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse
      & (fsm_output[30])) | ((~ return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse)
      & (fsm_output[32]));
  assign return_add_generic_AC_RND_CONV_false_12_and_33_cse = (~ return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse)
      & (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_12_and_39_cse = (~ or_547_cse) & (fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_12_and_25_cse = (~ or_673_cse) & (fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_12_and_27_cse = (~ or_1102_cse) & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_12_or_24_cse = return_add_generic_AC_RND_CONV_false_12_and_25_cse
      | return_add_generic_AC_RND_CONV_false_12_and_27_cse;
  assign return_add_generic_AC_RND_CONV_false_12_and_29_cse = (~ return_add_generic_AC_RND_CONV_false_6_op1_smaller_lor_lpi_3_dfm_2)
      & (fsm_output[11]);
  assign return_add_generic_AC_RND_CONV_false_12_and_31_cse = (~ return_add_generic_AC_RND_CONV_false_21_op1_smaller_return_add_generic_AC_RND_CONV_false_21_op1_smaller_or_cse)
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_12_and_35_cse = (~ return_add_generic_AC_RND_CONV_false_19_op1_smaller_lor_lpi_3_dfm_2)
      & (fsm_output[36]);
  assign return_add_generic_AC_RND_CONV_false_12_and_37_cse = (~ return_add_generic_AC_RND_CONV_false_8_op1_smaller_return_add_generic_AC_RND_CONV_false_8_op1_smaller_or_cse)
      & (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_12_and_30_cse = return_add_generic_AC_RND_CONV_false_6_op1_smaller_lor_lpi_3_dfm_2
      & (fsm_output[11]);
  assign return_add_generic_AC_RND_CONV_false_12_and_32_cse = return_add_generic_AC_RND_CONV_false_21_op1_smaller_return_add_generic_AC_RND_CONV_false_21_op1_smaller_or_cse
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_12_and_36_cse = return_add_generic_AC_RND_CONV_false_19_op1_smaller_lor_lpi_3_dfm_2
      & (fsm_output[36]);
  assign return_add_generic_AC_RND_CONV_false_12_and_38_cse = return_add_generic_AC_RND_CONV_false_8_op1_smaller_return_add_generic_AC_RND_CONV_false_8_op1_smaller_or_cse
      & (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_1_or_6_cse = return_add_generic_AC_RND_CONV_false_1_and_16_cse
      | return_add_generic_AC_RND_CONV_false_1_and_20_cse;
  assign return_add_generic_AC_RND_CONV_false_12_or_27_cse = BUTTERFLY_else_or_cse
      | or_dcpl_553 | return_add_generic_AC_RND_CONV_false_12_and_33_cse | return_add_generic_AC_RND_CONV_false_12_and_39_cse;
  assign return_add_generic_AC_RND_CONV_false_12_or_29_cse = return_add_generic_AC_RND_CONV_false_12_and_29_cse
      | return_add_generic_AC_RND_CONV_false_12_and_31_cse | return_add_generic_AC_RND_CONV_false_12_and_35_cse
      | return_add_generic_AC_RND_CONV_false_12_and_37_cse;
  assign return_add_generic_AC_RND_CONV_false_12_or_44_cse = return_add_generic_AC_RND_CONV_false_12_and_32_cse
      | return_add_generic_AC_RND_CONV_false_12_and_38_cse;
  assign or_2707_itm = (fsm_output[45]) | (fsm_output[20]) | (fsm_output[31]) | (fsm_output[6]);
  assign nl_operator_32_false_2_acc_5_itm = conv_u2u_10_11(~ z_out_101) + conv_u2u_4_11(in_u_rsci_q_d[15:12]);
  assign operator_32_false_2_acc_5_itm = nl_operator_32_false_2_acc_5_itm[10:0];
  assign and_3925_ssc = (and_2184_cse | (fsm_output[29]) | (fsm_output[31]) | (fsm_output[6])
      | (fsm_output[4]) | (fsm_output[32]) | (fsm_output[7]) | (fsm_output[9]) |
      (fsm_output[34]) | (fsm_output[12]) | (fsm_output[14]) | (fsm_output[38]))
      & run_wen;
  assign BUTTERFLY_1_else_1_if_and_1_rgt = (~ inverse_lpi_1_dfm_1) & or_1341_cse;
  assign BUTTERFLY_1_else_1_if_or_rgt = (inverse_lpi_1_dfm_1 & or_1341_cse) | or_1342_itm;
  assign return_add_generic_AC_RND_CONV_false_7_exp_and_2_ssc = return_add_generic_AC_RND_CONV_false_7_exp_and_ssc
      & (~(or_dcpl_521 | or_dcpl_476 | or_dcpl_240 | or_dcpl_236));
  assign return_add_generic_AC_RND_CONV_false_12_return_add_generic_AC_RND_CONV_false_12_nor_1_ssc
      = ~(return_add_generic_AC_RND_CONV_false_12_acc_2_itm_11_1 | (fsm_output[50]));
  assign return_add_generic_AC_RND_CONV_false_12_or_16_ssc = (return_add_generic_AC_RND_CONV_false_12_acc_2_itm_11_1
      & (~ (fsm_output[50]))) | (return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11_1
      & (fsm_output[50]));
  assign return_add_generic_AC_RND_CONV_false_12_and_6_ssc = (~ return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11_1)
      & (fsm_output[50]);
  assign return_add_generic_AC_RND_CONV_false_2_or_4_ssc = return_add_generic_AC_RND_CONV_false_2_and_cse
      | return_add_generic_AC_RND_CONV_false_2_and_10_cse;
  assign return_add_generic_AC_RND_CONV_false_2_or_6_ssc = return_add_generic_AC_RND_CONV_false_2_and_4_cse
      | return_add_generic_AC_RND_CONV_false_2_and_6_cse;
  assign return_add_generic_AC_RND_CONV_false_3_or_2_seb = (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[14]) | (fsm_output[18]) | (fsm_output[30]) | (fsm_output[32])
      | (fsm_output[39]) | (fsm_output[43]) | BUTTERFLY_else_or_cse;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      out1_rsci_idat_63 <= 1'b0;
      out1_rsci_idat_62_52 <= 11'b00000000000;
      out1_rsci_idat_51 <= 1'b0;
      out1_rsci_idat_50_0 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      out1_rsci_idat_63 <= 1'b0;
      out1_rsci_idat_62_52 <= 11'b00000000000;
      out1_rsci_idat_51 <= 1'b0;
      out1_rsci_idat_50_0 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( for_1_if_and_ssc ) begin
      out1_rsci_idat_63 <= MUX_s_1_2_2((out_f_d_rsci_q_d[63]), (in_f_d_rsci_q_d[63]),
          out1_rsci_idat_63_0_mx0c2);
      out1_rsci_idat_62_52 <= MUX1HOT_v_11_3_2((out_f_d_rsci_q_d[62:52]), return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_or_nl,
          (in_f_d_rsci_q_d[62:52]), {or_tmp_64 , out1_rsci_idat_63_0_mx0c1 , out1_rsci_idat_63_0_mx0c2});
      out1_rsci_idat_51 <= MUX1HOT_s_1_4_2((out_f_d_rsci_q_d[51]), (z_out_88[51]),
          return_mult_generic_AC_RND_CONV_false_6_op1_nan_sva_1, (in_f_d_rsci_q_d[51]),
          {or_tmp_64 , BUTTERFLY_if_1_and_nl , BUTTERFLY_if_1_and_1_nl , out1_rsci_idat_63_0_mx0c2});
      out1_rsci_idat_50_0 <= MUX1HOT_v_51_3_2((out_f_d_rsci_q_d[50:0]), return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_and_1_nl,
          (in_f_d_rsci_q_d[50:0]), {or_tmp_64 , out1_rsci_idat_63_0_mx0c1 , out1_rsci_idat_63_0_mx0c2});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      out1_rsci_idat_79_64 <= 16'b0000000000000000;
    end
    else if ( rst ) begin
      out1_rsci_idat_79_64 <= 16'b0000000000000000;
    end
    else if ( run_wen & (or_tmp_64 | out1_rsci_idat_79_64_mx0c1 | and_630_cse) )
        begin
      out1_rsci_idat_79_64 <= MUX1HOT_v_16_3_2(out_u_rsci_q_d, in_u_rsci_q_d, ({{1{stage_monty_mul_acc_2_psp_sva_1[14]}},
          stage_monty_mul_acc_2_psp_sva_1}), {or_tmp_64 , out1_rsci_idat_79_64_mx0c1
          , and_630_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_cgo_cse <= 1'b0;
      BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo <= 1'b0;
      BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo <= 1'b0;
      BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo <= 1'b0;
      BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo <= 1'b0;
      reg_out_u_triosy_obj_iswt0_cse <= 1'b0;
      reg_out1_rsci_iswt0_cse <= 1'b0;
      reg_out_u_rsci_cgo_ir_cse <= 1'b0;
      reg_out_f_d_rsci_cgo_ir_cse <= 1'b0;
      reg_in_u_rsci_cgo_ir_cse <= 1'b0;
      reg_in_f_d_rsci_cgo_ir_cse <= 1'b0;
      reg_ap_start_rsci_iswt0_cse <= 1'b0;
      reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_addr_cse <= 10'b0000000000;
      reg_BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_addr_cse <= 10'b0000000000;
      return_add_generic_AC_RND_CONV_false_12_mux_2_itm <= 1'b0;
      operator_32_false_1_acc_psp_sva_16_12 <= 5'b00000;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd <= 1'b0;
      operator_14_false_1_acc_psp_sva_12_10 <= 3'b000;
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_51 <= 1'b0;
    end
    else if ( rst ) begin
      reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_cgo_cse <= 1'b0;
      BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo <= 1'b0;
      BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo <= 1'b0;
      BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo <= 1'b0;
      BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo <= 1'b0;
      reg_out_u_triosy_obj_iswt0_cse <= 1'b0;
      reg_out1_rsci_iswt0_cse <= 1'b0;
      reg_out_u_rsci_cgo_ir_cse <= 1'b0;
      reg_out_f_d_rsci_cgo_ir_cse <= 1'b0;
      reg_in_u_rsci_cgo_ir_cse <= 1'b0;
      reg_in_f_d_rsci_cgo_ir_cse <= 1'b0;
      reg_ap_start_rsci_iswt0_cse <= 1'b0;
      reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_addr_cse <= 10'b0000000000;
      reg_BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_addr_cse <= 10'b0000000000;
      return_add_generic_AC_RND_CONV_false_12_mux_2_itm <= 1'b0;
      operator_32_false_1_acc_psp_sva_16_12 <= 5'b00000;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd <= 1'b0;
      operator_14_false_1_acc_psp_sva_12_10 <= 3'b000;
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_51 <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_cgo_cse <= or_dcpl_198
          | (fsm_output[4]) | (fsm_output[29]);
      BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_cgo <= inverse_lpi_1_dfm_1 & or_dcpl_200;
      BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_cgo <= (~ inverse_lpi_1_dfm_1) &
          or_dcpl_200;
      BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_cgo <= inverse_lpi_1_dfm_1 & or_dcpl_201;
      BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_cgo <= (~ inverse_lpi_1_dfm_1)
          & or_dcpl_201;
      reg_out_u_triosy_obj_iswt0_cse <= (z_out_113[10]) & (fsm_output[55]);
      reg_out1_rsci_iswt0_cse <= fsm_output[54];
      reg_out_u_rsci_cgo_ir_cse <= or_1119_rmff;
      reg_out_f_d_rsci_cgo_ir_cse <= or_1120_rmff;
      reg_in_u_rsci_cgo_ir_cse <= or_1121_rmff;
      reg_in_f_d_rsci_cgo_ir_cse <= or_1122_rmff;
      reg_ap_start_rsci_iswt0_cse <= ~ and_dcpl_202;
      reg_BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_addr_cse <= z_out_66;
      reg_BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_addr_cse <= return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0;
      return_add_generic_AC_RND_CONV_false_12_mux_2_itm <= MUX1HOT_s_1_16_2((~ return_add_generic_AC_RND_CONV_false_3_res_mant_3_0_sva_1),
          return_add_generic_AC_RND_CONV_false_3_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_2_res_mant_3_0_sva_1),
          return_add_generic_AC_RND_CONV_false_2_res_mant_3_0_sva_1, return_add_generic_AC_RND_CONV_false_8_res_mant_3_0_sva_1,
          (~ return_add_generic_AC_RND_CONV_false_8_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_12_res_mant_3_0_sva_1,
          (~ return_add_generic_AC_RND_CONV_false_12_res_mant_3_0_sva_1), (~ return_add_generic_AC_RND_CONV_false_16_res_mant_3_0_sva_1),
          return_add_generic_AC_RND_CONV_false_16_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_15_res_mant_3_0_sva_1),
          return_add_generic_AC_RND_CONV_false_15_res_mant_3_0_sva_1, return_add_generic_AC_RND_CONV_false_21_res_mant_3_0_sva_1,
          (~ return_add_generic_AC_RND_CONV_false_21_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_25_res_mant_3_0_sva_1,
          (~ return_add_generic_AC_RND_CONV_false_25_res_mant_3_0_sva_1), {return_add_generic_AC_RND_CONV_false_12_and_89_cse
          , return_add_generic_AC_RND_CONV_false_12_and_90_cse , return_add_generic_AC_RND_CONV_false_12_and_91_cse
          , return_add_generic_AC_RND_CONV_false_12_and_92_cse , return_add_generic_AC_RND_CONV_false_12_and_93_nl
          , return_add_generic_AC_RND_CONV_false_12_and_94_nl , return_add_generic_AC_RND_CONV_false_12_and_95_cse
          , return_add_generic_AC_RND_CONV_false_12_and_96_cse , return_add_generic_AC_RND_CONV_false_12_and_97_cse
          , return_add_generic_AC_RND_CONV_false_12_and_98_cse , return_add_generic_AC_RND_CONV_false_12_and_99_cse
          , return_add_generic_AC_RND_CONV_false_12_and_100_cse , return_add_generic_AC_RND_CONV_false_12_and_101_nl
          , return_add_generic_AC_RND_CONV_false_12_and_102_nl , return_add_generic_AC_RND_CONV_false_12_and_103_cse
          , return_add_generic_AC_RND_CONV_false_12_and_104_cse});
      operator_32_false_1_acc_psp_sva_16_12 <= MUX_v_5_2_2((stage_u_add_acc_1_itm_1[16:12]),
          (z_out_64[16:12]), BUTTERFLY_else_or_cse);
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd <= MUX_s_1_2_2((z_out_88[53]),
          (z_out_89[53]), return_add_generic_AC_RND_CONV_false_13_or_3_cse);
      operator_14_false_1_acc_psp_sva_12_10 <= MUX_v_3_2_2((z_out_86[12:10]), (z_out_68[12:10]),
          return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse);
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_51 <= MUX_s_1_2_2(stage_PE_tmp_re_d_1_lpi_3_dfm_51_mx0,
          stage_PE_1_tmp_im_d_1_lpi_3_dfm_51_mx1, or_dcpl_235);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & or_dcpl_284 & and_dcpl_204 & and_dcpl_203 & (fsm_output[6])
        ) begin
      return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_1_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_1_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[5])) | or_dcpl_289 | (~ return_add_generic_AC_RND_CONV_false_1_acc_2_itm_11_1)))
        ) begin
      return_add_generic_AC_RND_CONV_false_1_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & and_dcpl_210 & (fsm_output[14]) ) begin
      return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_else_4_unequal_tmp))
        & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
        & and_dcpl_204 & and_dcpl_203 & (fsm_output[8]) ) begin
      return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[7])) | or_dcpl_289 | (~ return_add_generic_AC_RND_CONV_false_acc_2_itm_11_1)))
        ) begin
      return_add_generic_AC_RND_CONV_false_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[9])) | or_dcpl_301 | and_dcpl_216 | (~
        mode_lpi_1_dfm) | return_add_generic_AC_RND_CONV_false_2_r_inf_lpi_3_dfm_2
        | or_dcpl_296)) ) begin
      return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & and_dcpl_210 & (fsm_output[12]) ) begin
      return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[10])) | or_dcpl_312 | return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2
        | or_dcpl_308 | and_dcpl_217)) ) begin
      return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & and_dcpl_224 & or_dcpl_320 & and_dcpl_219 & (fsm_output[13])
        ) begin
      return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (fsm_output[11]) & mode_lpi_1_dfm & return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1
        ) begin
      return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp <= ~((operator_33_true_12_acc_tmp[11:0]==12'b011111111111));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & and_dcpl_210 & (fsm_output[13]) ) begin
      return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & and_dcpl_231 & and_dcpl_229 & (fsm_output[16]) ) begin
      return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_7_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_7_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[15])) | and_836_cse)) ) begin
      return_add_generic_AC_RND_CONV_false_7_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & and_dcpl_237 & and_dcpl_235 & (fsm_output[18]) ) begin
      return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_8_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_8_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[17])) | and_840_cse)) ) begin
      return_add_generic_AC_RND_CONV_false_8_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & or_dcpl_342 & and_dcpl_204 & and_dcpl_203 & (fsm_output[31])
        ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_14_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_14_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[30])) | or_dcpl_289 | (~ return_add_generic_AC_RND_CONV_false_14_acc_2_itm_11_1)))
        ) begin
      return_add_generic_AC_RND_CONV_false_14_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & and_dcpl_210 & (fsm_output[39]) ) begin
      return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_13_else_4_unequal_tmp))
        & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
        & and_dcpl_204 & stage_PE_1_and_1_tmp & nand_102_cse & (fsm_output[33]) )
        begin
      return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_13_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_13_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[32])) | or_dcpl_289 | (~ return_add_generic_AC_RND_CONV_false_13_acc_2_itm_11_1)))
        ) begin
      return_add_generic_AC_RND_CONV_false_13_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[34])) | return_add_generic_AC_RND_CONV_false_15_r_inf_lpi_3_dfm_2
        | or_dcpl_312 | and_dcpl_251 | (~ mode_lpi_1_dfm) | or_dcpl_296)) ) begin
      return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & and_dcpl_210 & (fsm_output[37]) ) begin
      return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[35])) | or_dcpl_301 | return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2
        | or_dcpl_308 | and_dcpl_253)) ) begin
      return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & and_dcpl_224 & or_dcpl_371 & and_dcpl_219 & (fsm_output[38])
        ) begin
      return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (fsm_output[36]) & mode_lpi_1_dfm & return_add_generic_AC_RND_CONV_false_19_acc_2_itm_11_1
        ) begin
      return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp <= ~((operator_33_true_38_acc_tmp[11:0]==12'b011111111111));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & and_dcpl_210 & (fsm_output[38]) ) begin
      return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_1_if_acc_2_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & and_dcpl_259 & and_dcpl_229 & (fsm_output[41]) ) begin
      return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_20_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_20_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[40])) | and_836_cse)) ) begin
      return_add_generic_AC_RND_CONV_false_20_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & and_dcpl_263 & and_dcpl_235 & (fsm_output[43]) ) begin
      return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_21_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_21_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[42])) | and_840_cse)) ) begin
      return_add_generic_AC_RND_CONV_false_21_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[54])) | or_dcpl_190 | (operator_16_false_io_read_mode1_rsc_cse_sva[13:4]!=10'b0000000000)
        | or_dcpl_180 | or_dcpl_179 | operator_16_false_operator_16_false_nor_cse_sva
        | (return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp[11]))) ) begin
      return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_9_else_4_unequal_tmp))
        & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
        & and_dcpl_268 & and_dcpl_266 & nand_102_cse & (fsm_output[20]) ) begin
      return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_9_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_9_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[19])) | or_32_cse | (~ return_add_generic_AC_RND_CONV_false_9_acc_2_itm_11_1)))
        ) begin
      return_add_generic_AC_RND_CONV_false_9_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_10_else_4_unequal_tmp))
        & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
        & and_dcpl_276 & and_dcpl_274 & nand_102_cse & (fsm_output[22]) ) begin
      return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[21])) | or_32_cse | (~ return_add_generic_AC_RND_CONV_false_10_acc_2_itm_11_1)))
        ) begin
      return_add_generic_AC_RND_CONV_false_10_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & and_dcpl_285 & (~((~((~ (operator_33_true_12_acc_psp_sva[11]))
        & return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
        & and_dcpl_266 & nand_102_cse & (fsm_output[24]) ) begin
      return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[23])) | or_32_cse | (~ return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1)))
        ) begin
      return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & and_dcpl_223 & (~((~((~ (operator_33_true_12_acc_psp_sva[11]))
        & return_add_generic_AC_RND_CONV_false_12_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
        & and_dcpl_274 & nand_102_cse & (fsm_output[26]) ) begin
      return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[25])) | or_32_cse | (~ return_add_generic_AC_RND_CONV_false_12_acc_2_itm_11_1)))
        ) begin
      return_add_generic_AC_RND_CONV_false_12_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_22_else_4_unequal_tmp))
        & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
        & and_dcpl_268 & and_dcpl_274 & nand_102_cse & (fsm_output[45]) ) begin
      return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_22_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_22_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[44])) | or_32_cse | (~ return_add_generic_AC_RND_CONV_false_22_acc_2_itm_11_1)))
        ) begin
      return_add_generic_AC_RND_CONV_false_22_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_23_else_4_unequal_tmp))
        & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
        & and_dcpl_276 & and_dcpl_266 & nand_102_cse & (fsm_output[47]) ) begin
      return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_23_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_23_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[46])) | or_32_cse | (~ return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1)))
        ) begin
      return_add_generic_AC_RND_CONV_false_23_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_22_op1_inf_sva |
        return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva))
        & (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_24_else_4_unequal_tmp))
        & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
        & and_dcpl_274 & nand_102_cse & (fsm_output[49]) ) begin
      return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_24_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_24_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[48])) | or_32_cse | (~ return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11_1)))
        ) begin
      return_add_generic_AC_RND_CONV_false_24_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & and_dcpl_75 & (~ operator_11_true_return_22_sva) & (~((~((~
        (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_25_else_4_unequal_tmp))
        & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
        & and_dcpl_266 & nand_102_cse & (fsm_output[51]) ) begin
      return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_25_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_25_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ (fsm_output[50])) | or_32_cse | (~ return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11_1)))
        ) begin
      return_add_generic_AC_RND_CONV_false_25_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_8_else_4_return_add_generic_AC_RND_CONV_false_8_else_4_nand_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_16_false_io_read_mode1_rsc_cse_sva <= 16'b0000000000000000;
    end
    else if ( rst ) begin
      operator_16_false_io_read_mode1_rsc_cse_sva <= 16'b0000000000000000;
    end
    else if ( operator_16_false_and_cse & (~ operator_16_false_operator_16_false_nor_tmp)
        ) begin
      operator_16_false_io_read_mode1_rsc_cse_sva <= mode1_rsci_idat;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_16_false_operator_16_false_nor_cse_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_16_false_operator_16_false_nor_cse_sva <= 1'b0;
    end
    else if ( operator_16_false_and_cse ) begin
      operator_16_false_operator_16_false_nor_cse_sva <= operator_16_false_operator_16_false_nor_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      t_in_10_0_lpi_1_dfm_1_8 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_7 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_6 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_5 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_4 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_3 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_2 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_1 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_0 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_10 <= 1'b0;
      m_in_0_lpi_1_dfm <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_14 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_13 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_12 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_11 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_10 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_9 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_8 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_7 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_6 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_5 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_4 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_3 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_2 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_1 <= 1'b0;
    end
    else if ( rst ) begin
      t_in_10_0_lpi_1_dfm_1_8 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_7 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_6 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_5 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_4 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_3 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_2 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_1 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_0 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_10 <= 1'b0;
      m_in_0_lpi_1_dfm <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_14 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_13 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_12 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_11 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_10 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_9 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_8 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_7 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_6 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_5 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_4 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_3 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_2 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_1 <= 1'b0;
    end
    else if ( t_in_and_cse ) begin
      t_in_10_0_lpi_1_dfm_1_8 <= t_in_mux_nl & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_7 <= t_in_mux_2_nl & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_6 <= t_in_mux_3_nl & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_5 <= t_in_mux_4_nl & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_4 <= t_in_mux_5_nl & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_3 <= t_in_mux_6_nl & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_2 <= t_in_mux_7_nl & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_1 <= t_in_mux_8_nl & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_0 <= t_in_mux_9_nl & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_10 <= MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_10_mx0w0, need_ovf_1_need_ovf_1_and_nl,
          t_in_or_3_cse);
      m_in_0_lpi_1_dfm <= MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_10_mx0w0, need_ovf_1_need_ovf_1_and_1_nl,
          t_in_or_3_cse);
      m_in_15_1_lpi_1_dfm_1_14 <= m_in_mux_nl & t_in_or_3_cse;
      m_in_15_1_lpi_1_dfm_1_13 <= m_in_mux_14_nl & t_in_or_3_cse;
      m_in_15_1_lpi_1_dfm_1_12 <= m_in_mux_13_nl & t_in_or_3_cse;
      m_in_15_1_lpi_1_dfm_1_11 <= m_in_mux_12_nl & t_in_or_3_cse;
      m_in_15_1_lpi_1_dfm_1_10 <= m_in_mux_11_nl & t_in_or_3_cse;
      m_in_15_1_lpi_1_dfm_1_9 <= m_in_mux_10_nl & t_in_or_3_cse;
      m_in_15_1_lpi_1_dfm_1_8 <= m_in_mux_9_nl & t_in_or_3_cse;
      m_in_15_1_lpi_1_dfm_1_7 <= m_in_mux_8_nl & t_in_or_3_cse;
      m_in_15_1_lpi_1_dfm_1_6 <= m_in_mux_7_nl & t_in_or_3_cse;
      m_in_15_1_lpi_1_dfm_1_5 <= m_in_mux_6_nl & t_in_or_3_cse;
      m_in_15_1_lpi_1_dfm_1_4 <= m_in_mux_5_nl & t_in_or_3_cse;
      m_in_15_1_lpi_1_dfm_1_3 <= m_in_mux_4_nl & t_in_or_3_cse;
      m_in_15_1_lpi_1_dfm_1_2 <= m_in_mux_3_nl & t_in_or_3_cse;
      m_in_15_1_lpi_1_dfm_1_1 <= m_in_mux_2_nl & t_in_or_3_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      t_in_10_0_lpi_1_dfm_1_9 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_0 <= 1'b0;
    end
    else if ( rst ) begin
      t_in_10_0_lpi_1_dfm_1_9 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_0 <= 1'b0;
    end
    else if ( t_in_and_3_cse ) begin
      t_in_10_0_lpi_1_dfm_1_9 <= MUX_s_1_2_2(mode_lpi_1_dfm_mx0w0, t_in_10_0_lpi_1_dfm_1_10,
          t_in_or_3_cse);
      m_in_15_1_lpi_1_dfm_1_0 <= MUX_s_1_2_2(mode_lpi_1_dfm_mx0w0, m_in_0_lpi_1_dfm,
          t_in_or_3_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      mode_lpi_1_dfm <= 1'b0;
      inverse_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( rst ) begin
      mode_lpi_1_dfm <= 1'b0;
      inverse_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( mode_and_cse ) begin
      mode_lpi_1_dfm <= mode_lpi_1_dfm_mx0w0;
      inverse_lpi_1_dfm_1 <= ~(((mode1_rsci_idat==16'b0000000000000010)) | operator_16_false_operator_16_false_nor_tmp);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_i_3_0_sva <= 4'b0000;
    end
    else if ( rst ) begin
      for_i_3_0_sva <= 4'b0000;
    end
    else if ( ((or_2748_cse & t_in_or_3_cse) | (fsm_output[1])) & run_wen ) begin
      for_i_3_0_sva <= MUX_v_4_2_2(4'b0000, for_i_3_0_sva_2, not_932_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_qr_1_10_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_qr_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_index_const_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_15_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_index_const_10_lpi_2_dfm <= 1'b0;
    end
    else if ( rst ) begin
      stage_PE_1_qr_1_10_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_qr_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_index_const_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_15_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_index_const_10_lpi_2_dfm <= 1'b0;
    end
    else if ( stage_PE_1_and_2_cse ) begin
      stage_PE_1_qr_1_10_1_lpi_2_dfm_8 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_8,
          t_in_10_0_lpi_1_dfm_1_9, t_in_10_0_lpi_1_dfm_1_8, {(~ inverse_lpi_1_dfm_1)
          , and_6_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_7 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_7,
          t_in_10_0_lpi_1_dfm_1_8, t_in_10_0_lpi_1_dfm_1_7, {(~ inverse_lpi_1_dfm_1)
          , and_6_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_6 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_6,
          t_in_10_0_lpi_1_dfm_1_7, t_in_10_0_lpi_1_dfm_1_6, {(~ inverse_lpi_1_dfm_1)
          , and_6_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_5 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_5,
          t_in_10_0_lpi_1_dfm_1_6, t_in_10_0_lpi_1_dfm_1_5, {(~ inverse_lpi_1_dfm_1)
          , and_6_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_4 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_4,
          t_in_10_0_lpi_1_dfm_1_5, t_in_10_0_lpi_1_dfm_1_4, {(~ inverse_lpi_1_dfm_1)
          , and_6_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_3 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_3,
          t_in_10_0_lpi_1_dfm_1_4, t_in_10_0_lpi_1_dfm_1_3, {(~ inverse_lpi_1_dfm_1)
          , and_6_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_2 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_2,
          t_in_10_0_lpi_1_dfm_1_3, t_in_10_0_lpi_1_dfm_1_2, {(~ inverse_lpi_1_dfm_1)
          , and_6_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_1 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_1,
          t_in_10_0_lpi_1_dfm_1_2, t_in_10_0_lpi_1_dfm_1_1, {(~ inverse_lpi_1_dfm_1)
          , and_6_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_0 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_0,
          t_in_10_0_lpi_1_dfm_1_1, t_in_10_0_lpi_1_dfm_1_0, {(~ inverse_lpi_1_dfm_1)
          , and_6_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_10_1_lpi_2_dfm_8 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_8,
          t_in_10_0_lpi_1_dfm_1_9, or_tmp_231);
      stage_PE_1_qr_10_1_lpi_2_dfm_7 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_7,
          t_in_10_0_lpi_1_dfm_1_8, or_tmp_231);
      stage_PE_1_qr_10_1_lpi_2_dfm_6 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_6,
          t_in_10_0_lpi_1_dfm_1_7, or_tmp_231);
      stage_PE_1_qr_10_1_lpi_2_dfm_5 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_5,
          t_in_10_0_lpi_1_dfm_1_6, or_tmp_231);
      stage_PE_1_qr_10_1_lpi_2_dfm_4 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_4,
          t_in_10_0_lpi_1_dfm_1_5, or_tmp_231);
      stage_PE_1_qr_10_1_lpi_2_dfm_3 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_3,
          t_in_10_0_lpi_1_dfm_1_4, or_tmp_231);
      stage_PE_1_qr_10_1_lpi_2_dfm_2 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_2,
          t_in_10_0_lpi_1_dfm_1_3, or_tmp_231);
      stage_PE_1_qr_10_1_lpi_2_dfm_1 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_1,
          t_in_10_0_lpi_1_dfm_1_2, or_tmp_231);
      stage_PE_1_qr_10_1_lpi_2_dfm_0 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_0,
          t_in_10_0_lpi_1_dfm_1_1, or_tmp_231);
      stage_PE_1_qr_0_lpi_2_dfm <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_0, m_in_0_lpi_1_dfm,
          t_in_10_0_lpi_1_dfm_1_10, {and_994_nl , and_996_nl , or_tmp_231});
      stage_PE_1_index_const_9_1_lpi_2_dfm_8 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_8,
          t_in_10_0_lpi_1_dfm_1_10, or_tmp_231);
      stage_PE_1_index_const_9_1_lpi_2_dfm_7 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_7,
          t_in_10_0_lpi_1_dfm_1_9, or_tmp_231);
      stage_PE_1_index_const_9_1_lpi_2_dfm_6 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_6,
          t_in_10_0_lpi_1_dfm_1_8, or_tmp_231);
      stage_PE_1_index_const_9_1_lpi_2_dfm_5 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_5,
          t_in_10_0_lpi_1_dfm_1_7, or_tmp_231);
      stage_PE_1_index_const_9_1_lpi_2_dfm_4 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_4,
          t_in_10_0_lpi_1_dfm_1_6, or_tmp_231);
      stage_PE_1_index_const_9_1_lpi_2_dfm_3 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_3,
          t_in_10_0_lpi_1_dfm_1_5, or_tmp_231);
      stage_PE_1_index_const_9_1_lpi_2_dfm_2 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_2,
          t_in_10_0_lpi_1_dfm_1_4, or_tmp_231);
      stage_PE_1_index_const_9_1_lpi_2_dfm_1 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_1,
          t_in_10_0_lpi_1_dfm_1_3, or_tmp_231);
      stage_PE_1_index_const_9_1_lpi_2_dfm_0 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_0,
          t_in_10_0_lpi_1_dfm_1_2, or_tmp_231);
      stage_PE_1_index_const_0_lpi_2_dfm <= MUX_s_1_2_2(stage_PE_qif_qelse_mux_nl,
          t_in_10_0_lpi_1_dfm_1_1, or_tmp_231);
      stage_PE_1_index_const_15_lpi_2_dfm <= m_in_15_1_lpi_1_dfm_1_14 & (~ mode_lpi_1_dfm)
          & inverse_lpi_1_dfm_1;
      stage_PE_1_index_const_14_11_lpi_2_dfm_3 <= stage_PE_qif_qelse_mux_1_nl & inverse_lpi_1_dfm_1;
      stage_PE_1_index_const_14_11_lpi_2_dfm_2 <= stage_PE_qif_qelse_mux_14_nl &
          inverse_lpi_1_dfm_1;
      stage_PE_1_index_const_14_11_lpi_2_dfm_1 <= stage_PE_qif_qelse_mux_13_nl &
          inverse_lpi_1_dfm_1;
      stage_PE_1_index_const_14_11_lpi_2_dfm_0 <= stage_PE_qif_qelse_mux_12_nl &
          inverse_lpi_1_dfm_1;
      stage_PE_1_index_const_10_lpi_2_dfm <= stage_PE_qif_qelse_mux_11_nl & inverse_lpi_1_dfm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_qr_1_0_lpi_2_dfm <= 1'b0;
    end
    else if ( rst ) begin
      stage_PE_1_qr_1_0_lpi_2_dfm <= 1'b0;
    end
    else if ( stage_PE_1_and_2_cse & (~ inverse_lpi_1_dfm_1) ) begin
      stage_PE_1_qr_1_0_lpi_2_dfm <= m_in_0_lpi_1_dfm;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_n_9_0_sva_8_0 <= 9'b000000000;
    end
    else if ( rst ) begin
      BUTTERFLY_1_n_9_0_sva_8_0 <= 9'b000000000;
    end
    else if ( run_wen & ((fsm_output[0]) | (fsm_output[56]) | (fsm_output[1]) | (fsm_output[2])
        | (fsm_output[55]) | (fsm_output[54]) | (fsm_output[53]) | t_in_or_3_cse)
        ) begin
      BUTTERFLY_1_n_9_0_sva_8_0 <= MUX_v_9_2_2(9'b000000000, (z_out_101[8:0]), t_in_or_3_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_26_m_zero_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_26_m_zero_sva <= 1'b0;
    end
    else if ( run_wen & ((~(inverse_lpi_1_dfm_1 | (and_dcpl_323 & and_dcpl_333 &
        and_dcpl_369 & nor_35_cse))) | (fsm_output[2])) ) begin
      return_extract_26_m_zero_sva <= MUX1HOT_s_1_3_2(stage_PE_1_and_1_tmp, return_extract_3_m_zero_sva_mx1w0,
          return_extract_56_m_zero_sva_mx2w0, {(fsm_output[2]) , (fsm_output[4])
          , (fsm_output[29])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0 <= 10'b0000000000;
      operator_33_true_12_acc_psp_sva <= 13'b0000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0 <= 10'b0000000000;
      operator_33_true_12_acc_psp_sva <= 13'b0000000000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_19_exp_plus_1_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0 <= MUX1HOT_v_10_3_2(or_2026_nl,
          (return_add_generic_AC_RND_CONV_false_6_exp_plus_1_12_1_lpi_3_dfm_1[9:0]),
          (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_2[9:0]),
          {and_1068_nl , (fsm_output[11]) , (fsm_output[36])});
      operator_33_true_12_acc_psp_sva <= MUX1HOT_v_13_4_2(z_out_84, operator_33_true_12_acc_tmp,
          z_out_85, operator_33_true_38_acc_tmp, {return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse
          , (fsm_output[11]) , operator_33_true_12_or_1_nl , (fsm_output[36])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_fry_9_0_sva <= 10'b0000000000;
    end
    else if ( rst ) begin
      BUTTERFLY_1_fry_9_0_sva <= 10'b0000000000;
    end
    else if ( run_wen & (~(and_dcpl_405 & and_dcpl_403 & and_dcpl_402 & (~((fsm_output[56])
        | (fsm_output[1]))) & and_dcpl_333 & (~((fsm_output[25]) | (fsm_output[54])
        | (fsm_output[53]))))) ) begin
      BUTTERFLY_1_fry_9_0_sva <= z_out_67;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_BUTTERFLY_1_i_9_0_ftd <= 1'b0;
    end
    else if ( rst ) begin
      reg_BUTTERFLY_1_i_9_0_ftd <= 1'b0;
    end
    else if ( BUTTERFLY_1_i_and_ssc ) begin
      reg_BUTTERFLY_1_i_9_0_ftd <= BUTTERFLY_i_9_0_sva_1[9];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_BUTTERFLY_1_i_9_0_ftd_1 <= 9'b000000000;
    end
    else if ( rst ) begin
      reg_BUTTERFLY_1_i_9_0_ftd_1 <= 9'b000000000;
    end
    else if ( BUTTERFLY_1_i_and_ssc & (~ or_tmp_450) ) begin
      reg_BUTTERFLY_1_i_9_0_ftd_1 <= MUX_v_9_2_2((BUTTERFLY_i_9_0_sva_1[8:0]), (BUTTERFLY_1_fry_9_0_sva[8:0]),
          BUTTERFLY_i_or_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm <= 1'b0;
    end
    else if ( rst ) begin
      BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm <= 1'b0;
    end
    else if ( run_wen & (~(nor_34_cse & (~ (fsm_output[3])) & and_dcpl_402 & (~ (fsm_output[56]))
        & and_dcpl_329 & (~ (fsm_output[55])) & nor_35_cse)) & mode_lpi_1_dfm ) begin
      BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm <= (BUTTERFLY_1_n_9_0_sva_8_0==9'b011111111);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_unequal_tmp <= 1'b0;
      operator_11_true_return_26_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_unequal_tmp <= 1'b0;
      operator_11_true_return_26_sva <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_10_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_10_unequal_tmp <= MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp,
          return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0, return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp,
          return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_mx2w0, return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1,
          {(fsm_output[4]) , BUTTERFLY_if_1_if_or_cse , (fsm_output[29]) , (fsm_output[31])
          , (fsm_output[47])});
      operator_11_true_return_26_sva <= MUX1HOT_s_1_5_2(operator_11_true_3_operator_11_true_3_and_tmp,
          return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0, operator_11_true_35_operator_11_true_35_and_tmp,
          return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0, return_mult_generic_AC_RND_CONV_false_1_op1_zero_sva_1,
          {(fsm_output[4]) , BUTTERFLY_if_1_if_or_cse , (fsm_output[29]) , (fsm_output[31])
          , (fsm_output[47])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm
          <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm
          <= 1'b0;
    end
    else if ( run_wen & (~ return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse)
        ) begin
      return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm
          <= MUX1HOT_s_1_9_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1,
          (return_add_generic_AC_RND_CONV_false_res_rounded_lpi_3_dfm_51_0_1[51]),
          return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm_mx1,
          (return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1[50]), drf_qr_lval_15_smx_0_lpi_3_dfm_mx2,
          (return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1[51]),
          return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm_mx3,
          BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx5, {(fsm_output[4])
          , return_add_generic_AC_RND_CONV_false_13_or_cse , (fsm_output[10]) , return_add_generic_AC_RND_CONV_false_13_or_4_cse
          , return_add_generic_AC_RND_CONV_false_13_and_2_cse , return_add_generic_AC_RND_CONV_false_13_or_3_cse
          , (fsm_output[29]) , (fsm_output[35]) , return_add_generic_AC_RND_CONV_false_13_and_4_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_13_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      drf_qr_lval_13_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & ((inverse_lpi_1_dfm_1 & (~(or_dcpl_522 | or_dcpl_516 | (fsm_output[17])
        | or_dcpl_515 | or_dcpl_245 | (fsm_output[13]) | or_dcpl_511 | or_dcpl_509
        | (fsm_output[5]) | (fsm_output[12])))) | (fsm_output[4]) | (fsm_output[18])
        | (fsm_output[31]) | (fsm_output[35]) | (fsm_output[37]) | (fsm_output[43]))
        ) begin
      drf_qr_lval_13_smx_0_lpi_3_dfm <= MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_10_exp_mux1h_3_cse, return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_1,
          drf_qr_lval_13_smx_0_lpi_3_dfm_mx3, return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_3_nl,
          return_add_generic_AC_RND_CONV_false_10_exp_mux1h_6_cse, {return_add_generic_AC_RND_CONV_false_13_or_2_cse
          , (fsm_output[18]) , (fsm_output[31]) , (fsm_output[35]) , (fsm_output[37])
          , (fsm_output[43])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_12_m_zero_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_12_m_zero_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_535 | or_dcpl_532 | (fsm_output[17]) | or_dcpl_529
        | (fsm_output[15]) | or_dcpl_528)) ) begin
      return_extract_12_m_zero_sva <= MUX1HOT_s_1_7_2(return_extract_3_m_zero_sva_mx1w0,
          return_extract_12_m_zero_return_extract_12_m_zero_nor_nl, return_extract_20_m_zero_return_extract_20_m_zero_nor_nl,
          return_extract_25_m_zero_return_extract_25_m_zero_nor_nl, return_extract_56_m_zero_sva_mx2w0,
          return_extract_53_m_zero_return_extract_53_m_zero_nor_nl, return_extract_59_m_zero_return_extract_59_m_zero_nor_nl,
          {return_add_generic_AC_RND_CONV_false_13_or_2_cse , or_dcpl_208 , (fsm_output[12])
          , (fsm_output[16]) , or_tmp_334 , (fsm_output[39]) , (fsm_output[43])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_1_sva <= 1'b0;
    end
    else if ( run_wen & (~((fsm_output[50]) | (fsm_output[49]) | (fsm_output[42])
        | or_dcpl_534 | or_dcpl_545 | (fsm_output[43]) | or_dcpl_532 | or_dcpl_502
        | (fsm_output[7]) | return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse
        | (fsm_output[15]) | (fsm_output[30]) | (fsm_output[40]) | (fsm_output[5])))
        ) begin
      operator_11_true_return_1_sva <= MUX1HOT_s_1_9_2(operator_11_true_3_operator_11_true_3_and_tmp,
          operator_11_true_12_operator_11_true_12_and_nl, operator_11_true_52_operator_11_true_52_and_nl,
          operator_11_true_25_operator_11_true_25_and_nl, return_add_generic_AC_RND_CONV_false_6_r_nan_and_2,
          operator_11_true_35_operator_11_true_35_and_tmp, operator_11_true_44_operator_11_true_44_and_nl,
          operator_11_true_57_operator_11_true_57_and_nl, return_add_generic_AC_RND_CONV_false_25_r_nan_and_nl,
          {return_add_generic_AC_RND_CONV_false_13_or_2_cse , or_dcpl_208 , or_dcpl_484
          , (fsm_output[16]) , (fsm_output[23]) , or_tmp_334 , or_dcpl_235 , (fsm_output[41])
          , (fsm_output[48])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & ((~(reg_return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_rgt_nl
        | return_add_generic_AC_RND_CONV_false_10_ls_or_2_cse | (fsm_output[17])
        | or_dcpl_562 | or_dcpl_560 | or_dcpl_559 | or_dcpl_511 | (fsm_output[36])
        | or_dcpl_555 | or_dcpl_554)) | (fsm_output[4]) | (fsm_output[29]) | (fsm_output[31]))
        ) begin
      return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm <= MUX1HOT_v_51_6_2(return_extract_2_mux_4_cse,
          (out_f_d_rsci_q_d[51:1]), (out_f_d_rsci_q_d[50:0]), return_extract_33_mux_3_cse,
          (in_f_d_rsci_q_d[51:1]), (in_f_d_rsci_q_d[50:0]), {return_add_generic_AC_RND_CONV_false_13_op2_mu_or_6_nl
          , return_add_generic_AC_RND_CONV_false_13_op2_mu_and_2_nl , return_add_generic_AC_RND_CONV_false_13_op2_mu_and_3_nl
          , return_add_generic_AC_RND_CONV_false_13_op2_mu_or_8_nl , return_add_generic_AC_RND_CONV_false_13_op2_mu_and_4_nl
          , return_add_generic_AC_RND_CONV_false_13_op2_mu_and_5_nl});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_tmp_re_d_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      stage_PE_1_tmp_re_d_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & ((inverse_lpi_1_dfm_1 & (~(or_dcpl_590 | or_dcpl_588 | (fsm_output[16])
        | or_dcpl_586 | or_dcpl_584 | or_dcpl_511 | (fsm_output[30]) | or_dcpl_580
        | or_dcpl_553 | (fsm_output[5]) | or_dcpl_576))) | (fsm_output[4]) | (fsm_output[29]))
        ) begin
      stage_PE_1_tmp_re_d_sva <= MUX_v_64_2_2(out_f_d_rsci_q_d, in_f_d_rsci_q_d,
          stage_PE_1_tmp_re_d_or_3_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_21_smx_9_0_lpi_3_dfm <= 10'b0000000000;
    end
    else if ( rst ) begin
      drf_qr_lval_21_smx_9_0_lpi_3_dfm <= 10'b0000000000;
    end
    else if ( run_wen & (~(or_dcpl_621 | or_dcpl_602 | or_dcpl_519 | (fsm_output[21])
        | (fsm_output[34]) | (fsm_output[7]) | or_dcpl_269 | or_dcpl_597)) ) begin
      drf_qr_lval_21_smx_9_0_lpi_3_dfm <= MUX1HOT_v_10_5_2((r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[61:52]),
          (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[61:52]), return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1,
          (stage_PE_1_tmp_re_d_sva[62:53]), return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1,
          {return_add_generic_AC_RND_CONV_false_18_exp_and_1_nl , return_add_generic_AC_RND_CONV_false_18_exp_and_2_itm
          , return_add_generic_AC_RND_CONV_false_18_exp_and_3_cse , return_add_generic_AC_RND_CONV_false_18_exp_or_cse
          , return_add_generic_AC_RND_CONV_false_18_exp_and_5_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_11_op_bigger_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm <= MUX1HOT_s_1_11_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
          drf_qr_lval_13_smx_0_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_2_nl,
          return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0,
          (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[50]), return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0,
          (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[50]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_7_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_8_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_9_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse , (fsm_output[14])
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_10_cse , (fsm_output[39])
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse , and_1046_cse});
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm <= MUX1HOT_s_1_11_2(return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_13_op2_mu_0_lpi_3_dfm_1,
          (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[50]), BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx2,
          return_add_generic_AC_RND_CONV_false_7_mux_27_cse, return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_20_mux_27_cse, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1,
          {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_7_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_8_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_9_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_21_nl
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_22_nl , (fsm_output[14])
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse , or_1302_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_10_cse , (fsm_output[39])
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_628 | or_dcpl_635)) ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm <= MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm_mx1w0,
          return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_23_op1_mu_52_lpi_3_dfm,
          return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm, {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_16_nl , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_32_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse
          , and_1046_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_50 <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_50 <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_12_op_bigger_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm <= MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm_mx1w0,
          return_add_generic_AC_RND_CONV_false_10_op2_mu_1_51_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[50]),
          return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[50]),
          {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse , return_add_generic_AC_RND_CONV_false_18_exp_and_3_cse
          , return_add_generic_AC_RND_CONV_false_18_exp_and_4_cse , return_add_generic_AC_RND_CONV_false_18_exp_and_5_cse
          , return_add_generic_AC_RND_CONV_false_18_exp_and_6_cse});
      return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_50 <= return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_mx1w0[50];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_18_op_bigger_mux_1_itm_50 <= 1'b0;
      return_add_generic_AC_RND_CONV_false_18_op_bigger_mux_1_itm_49_0 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_18_op_bigger_mux_1_itm_50 <= 1'b0;
      return_add_generic_AC_RND_CONV_false_18_op_bigger_mux_1_itm_49_0 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_12_op_bigger_and_1_cse ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm <= MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm_mx1w0,
          return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1, {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse
          , return_add_generic_AC_RND_CONV_false_18_exp_and_3_cse , return_add_generic_AC_RND_CONV_false_18_exp_or_cse
          , return_add_generic_AC_RND_CONV_false_18_exp_and_5_cse});
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_itm <= MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm_mx1w0,
          return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx0, drf_qr_lval_13_smx_0_lpi_3_dfm,
          return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_23_op1_mu_52_lpi_3_dfm,
          {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse , return_add_generic_AC_RND_CONV_false_18_exp_and_3_cse
          , return_add_generic_AC_RND_CONV_false_18_exp_and_4_cse , return_add_generic_AC_RND_CONV_false_18_exp_and_5_cse
          , return_add_generic_AC_RND_CONV_false_18_exp_and_6_cse});
      return_add_generic_AC_RND_CONV_false_18_op_bigger_mux_1_itm_50 <= return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_mx1w0[50];
      return_add_generic_AC_RND_CONV_false_18_op_bigger_mux_1_itm_49_0 <= MUX1HOT_v_50_5_2((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_mx1w0[49:0]),
          return_add_generic_AC_RND_CONV_false_10_op2_mu_1_50_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49:0]),
          return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[49:0]),
          {(~ or_dcpl_625) , or_tmp_946 , return_add_generic_AC_RND_CONV_false_18_exp_and_4_cse
          , or_1993_cse , return_add_generic_AC_RND_CONV_false_18_exp_and_6_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_41_return_extract_41_or_1_cse_sva <= 1'b0;
      stage_PE_1_gm_im_d_61_0_lpi_3_dfm <= 62'b00000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_extract_41_return_extract_41_or_1_cse_sva <= 1'b0;
      stage_PE_1_gm_im_d_61_0_lpi_3_dfm <= 62'b00000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( return_extract_41_and_1_cse ) begin
      return_extract_41_return_extract_41_or_1_cse_sva <= return_extract_41_return_extract_41_or_1_cse_sva_1;
      stage_PE_1_gm_im_d_61_0_lpi_3_dfm <= r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_11_mux_1_itm <= 56'b00000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_11_mux_1_itm <= 56'b00000000000000000000000000000000000000000000000000000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_11_op_smaller_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm <= MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx1w0,
          return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2,
          return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx3,
          {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse , (fsm_output[16])
          , (fsm_output[41])});
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm <= MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx1w0,
          return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx2,
          return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx4,
          {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse , (fsm_output[16])
          , (fsm_output[41])});
      return_add_generic_AC_RND_CONV_false_11_mux_1_itm <= MUX1HOT_v_56_4_2((~ (z_out_74[56:1])),
          (z_out_74[56:1]), (z_out_76[56:1]), (~ (z_out_76[56:1])), {return_add_generic_AC_RND_CONV_false_11_or_nl
          , return_add_generic_AC_RND_CONV_false_11_or_6_nl , return_add_generic_AC_RND_CONV_false_11_or_7_nl
          , return_add_generic_AC_RND_CONV_false_11_or_8_nl});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm <= 1'b0;
    end
    else if ( (((~(z_out_53_52 & return_add_generic_AC_RND_CONV_false_22_e1_eq_e2_equal_tmp))
        & (~ (z_out_96[11])) & (fsm_output[41])) | (fsm_output[16]) | (fsm_output[12])
        | (fsm_output[10]) | (fsm_output[30]) | (fsm_output[5]) | (fsm_output[32]))
        & run_wen ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm <= MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx1w0,
          return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx1,
          return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_3_nl,
          return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx2,
          return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx3,
          {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse , (fsm_output[10])
          , (fsm_output[12]) , (fsm_output[16]) , (fsm_output[32]) , (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm <= 1'b0;
    end
    else if ( rst ) begin
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm <= 1'b0;
    end
    else if ( run_wen & ((inverse_lpi_1_dfm_1 & (~(or_dcpl_664 | (fsm_output[18])
        | (fsm_output[7]) | (fsm_output[38]) | (fsm_output[8]) | or_dcpl_466))) |
        (fsm_output[5]) | BUTTERFLY_else_or_cse | or_dcpl_208 | (fsm_output[13])
        | (fsm_output[16]) | or_tmp_450 | BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx0c8
        | (fsm_output[30]) | or_dcpl_235 | (fsm_output[37]) | (fsm_output[41])) )
        begin
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm <= MUX1HOT_s_1_11_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx1w0,
          return_add_generic_AC_RND_CONV_false_4_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_4_res_mant_3_0_sva_1),
          return_extract_12_return_extract_12_or_1_cse_sva_1, BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx2,
          BUTTERFLY_1_fiy_mux1h_4_cse, (BUTTERFLY_1_fry_9_0_sva[9]), reg_BUTTERFLY_1_i_9_0_ftd,
          return_extract_44_return_extract_44_or_1_cse_sva_1, BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx5,
          BUTTERFLY_1_fiy_mux1h_10_cse, {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_3_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_4_cse
          , or_dcpl_208 , (fsm_output[13]) , (fsm_output[16]) , return_add_generic_AC_RND_CONV_false_11_op_smaller_or_nl
          , or_tmp_450 , or_dcpl_235 , (fsm_output[37]) , (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_19_smx_lpi_3_dfm <= 11'b00000000000;
    end
    else if ( rst ) begin
      drf_qr_lval_19_smx_lpi_3_dfm <= 11'b00000000000;
    end
    else if ( run_wen & (~(or_dcpl_586 | or_dcpl_680 | or_dcpl_679)) ) begin
      drf_qr_lval_19_smx_lpi_3_dfm <= MUX1HOT_v_11_3_2(drf_qr_lval_1_smx_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_and_2_nl,
          return_extract_32_mux_cse, {(fsm_output[5]) , operator_6_false_17_or_cse
          , (fsm_output[30])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva
          <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva
          <= 1'b0;
    end
    else if ( run_wen & (~(operator_6_false_17_or_cse | or_dcpl_484)) ) begin
      return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva
          <= MUX1HOT_s_1_20_2(return_add_generic_AC_RND_CONV_false_1_acc_2_itm_11_1,
          return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp,
          return_add_generic_AC_RND_CONV_false_acc_2_itm_11_1, return_add_generic_AC_RND_CONV_false_17_acc_3_itm_10,
          return_add_generic_AC_RND_CONV_false_6_acc_2_itm_11_1, return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp,
          return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1, return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1,
          return_add_generic_AC_RND_CONV_false_9_acc_2_itm_11_1, return_add_generic_AC_RND_CONV_false_10_acc_2_itm_11_1,
          return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1, return_add_generic_AC_RND_CONV_false_12_acc_2_itm_11_1,
          return_add_generic_AC_RND_CONV_false_14_acc_2_itm_11_1, return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp,
          return_add_generic_AC_RND_CONV_false_13_acc_2_itm_11_1, return_add_generic_AC_RND_CONV_false_19_acc_2_itm_11_1,
          return_add_generic_AC_RND_CONV_false_22_acc_2_itm_11_1, return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1,
          return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11_1, return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11_1,
          {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse
          , (fsm_output[11]) , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse
          , or_dcpl_493 , or_dcpl_485 , (fsm_output[19]) , (fsm_output[21]) , (fsm_output[23])
          , (fsm_output[25]) , (fsm_output[30]) , (fsm_output[31]) , (fsm_output[32])
          , (fsm_output[36]) , (fsm_output[44]) , (fsm_output[46]) , (fsm_output[48])
          , (fsm_output[50])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_17_mux_6_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_17_mux_6_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_485 | return_add_generic_AC_RND_CONV_false_11_or_4_cse
        | or_dcpl_645 | or_dcpl_686 | or_dcpl_685 | or_dcpl_597)) ) begin
      return_add_generic_AC_RND_CONV_false_17_mux_6_itm <= MUX1HOT_s_1_7_2(return_add_generic_AC_RND_CONV_false_4_if_2_return_add_generic_AC_RND_CONV_false_4_if_2_nor_1_nl,
          (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[63]), (~ inverse_lpi_1_dfm_1),
          return_mult_generic_AC_RND_CONV_false_1_op1_zero_sva_1, return_add_generic_AC_RND_CONV_false_17_mux_6_itm_mx2,
          return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0, return_add_generic_AC_RND_CONV_false_17_mux_6_itm_mx4,
          {return_add_generic_AC_RND_CONV_false_17_and_1_cse , return_add_generic_AC_RND_CONV_false_17_and_3_cse
          , return_add_generic_AC_RND_CONV_false_17_and_4_cse , or_756_nl , (fsm_output[14])
          , or_1538_nl , (fsm_output[39])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_520 | (fsm_output[42]) | or_dcpl_664 | or_dcpl_702
        | or_dcpl_562 | or_dcpl_699 | or_dcpl_686 | (fsm_output[40]) | or_dcpl_679))
        ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_itm <= MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_5_if_2_return_add_generic_AC_RND_CONV_false_5_if_2_and_2_nl,
          (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[63]), inverse_lpi_1_dfm_1,
          return_add_generic_AC_RND_CONV_false_9_do_sub_return_add_generic_AC_RND_CONV_false_9_do_sub_xor_nl,
          return_add_generic_AC_RND_CONV_false_23_do_sub_return_add_generic_AC_RND_CONV_false_23_do_sub_xor_nl,
          {return_add_generic_AC_RND_CONV_false_17_and_1_cse , return_add_generic_AC_RND_CONV_false_17_and_3_cse
          , return_add_generic_AC_RND_CONV_false_17_and_4_cse , (fsm_output[14])
          , (fsm_output[39])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_mux_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_mux_itm <= 1'b0;
    end
    else if ( run_wen & ((~(inverse_lpi_1_dfm_1 | (and_dcpl_421 & and_dcpl_323 &
        (~((fsm_output[2]) | (fsm_output[49]) | (fsm_output[55]))) & and_dcpl_369
        & and_dcpl_354 & (~((fsm_output[16]) | (fsm_output[7]))) & (~((fsm_output[30])
        | (fsm_output[54]) | (fsm_output[53]))) & (~ (fsm_output[31]))))) | (fsm_output[5])
        | (fsm_output[18]) | (fsm_output[32]) | (fsm_output[41])) ) begin
      return_add_generic_AC_RND_CONV_false_12_mux_itm <= MUX1HOT_s_1_13_2(return_add_generic_AC_RND_CONV_false_3_if_2_return_add_generic_AC_RND_CONV_false_3_if_2_nor_1_nl,
          (stage_PE_1_tmp_re_d_sva[63]), (~ (out_f_d_rsci_q_d[63])), return_extract_3_m_zero_sva_mx1w0,
          return_add_generic_AC_RND_CONV_false_12_if_2_return_add_generic_AC_RND_CONV_false_12_if_2_nor_mx3w0,
          (~ return_add_generic_AC_RND_CONV_false_17_mux_6_itm), return_add_generic_AC_RND_CONV_false_15_if_2_return_add_generic_AC_RND_CONV_false_15_if_2_nor_1_nl,
          (in_f_d_rsci_q_d[63]), (~ (stage_PE_1_tmp_re_d_sva[63])), return_extract_56_m_zero_sva_mx2w0,
          return_add_generic_AC_RND_CONV_false_11_if_2_return_add_generic_AC_RND_CONV_false_11_if_2_nor_mx5w0,
          (stage_PE_1_x_re_d_sva[63]), (~ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1),
          {return_add_generic_AC_RND_CONV_false_12_and_105_cse , return_add_generic_AC_RND_CONV_false_12_or_46_nl
          , return_add_generic_AC_RND_CONV_false_12_and_116_cse , (fsm_output[7])
          , return_add_generic_AC_RND_CONV_false_12_and_107_cse , return_add_generic_AC_RND_CONV_false_12_and_118_cse
          , return_add_generic_AC_RND_CONV_false_12_and_109_cse , return_add_generic_AC_RND_CONV_false_12_and_110_cse
          , return_add_generic_AC_RND_CONV_false_12_and_111_cse , return_add_generic_AC_RND_CONV_false_12_and_112_cse
          , return_add_generic_AC_RND_CONV_false_12_and_113_cse , return_add_generic_AC_RND_CONV_false_12_and_119_cse
          , return_add_generic_AC_RND_CONV_false_12_and_120_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_do_sub_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_do_sub_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_627 | or_dcpl_236 | or_dcpl_625 | or_dcpl_588
        | or_dcpl_515 | (fsm_output[15]) | or_dcpl_685 | or_dcpl_597)) ) begin
      return_add_generic_AC_RND_CONV_false_10_do_sub_sva <= MUX1HOT_s_1_7_2(return_add_generic_AC_RND_CONV_false_17_do_sub_return_add_generic_AC_RND_CONV_false_17_do_sub_return_add_generic_AC_RND_CONV_false_17_do_sub_xnor_nl,
          return_mult_generic_AC_RND_CONV_false_op2_zero_sva_1, return_mult_generic_AC_RND_CONV_false_1_op2_zero_sva_1,
          return_add_generic_AC_RND_CONV_false_10_do_sub_return_add_generic_AC_RND_CONV_false_10_do_sub_xor_nl,
          return_mult_generic_AC_RND_CONV_false_3_op2_zero_sva_1, return_mult_generic_AC_RND_CONV_false_4_op2_zero_sva_1,
          return_add_generic_AC_RND_CONV_false_22_do_sub_return_add_generic_AC_RND_CONV_false_22_do_sub_xor_nl,
          {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse , (fsm_output[11])
          , (fsm_output[12]) , (fsm_output[14]) , (fsm_output[36]) , (fsm_output[37])
          , (fsm_output[39])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_do_sub_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_do_sub_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_605 | (fsm_output[42]) | or_dcpl_728 | or_dcpl_726
        | or_dcpl_626 | return_add_generic_AC_RND_CONV_false_11_or_4_cse | (fsm_output[34])
        | or_dcpl_698 | (fsm_output[15]) | or_dcpl_719 | or_dcpl_633)) ) begin
      return_add_generic_AC_RND_CONV_false_11_do_sub_sva <= MUX1HOT_s_1_11_2(return_add_generic_AC_RND_CONV_false_18_do_sub_return_add_generic_AC_RND_CONV_false_18_do_sub_xor_nl,
          return_mult_generic_AC_RND_CONV_false_r_nan_or_nl, return_mult_generic_AC_RND_CONV_false_1_r_nan_or_nl,
          return_mult_generic_AC_RND_CONV_false_2_r_nan_or_nl, return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_xnor_nl,
          return_add_generic_AC_RND_CONV_false_11_r_nan_and_nl, return_mult_generic_AC_RND_CONV_false_3_r_nan_or_nl,
          return_mult_generic_AC_RND_CONV_false_4_r_nan_or_nl, return_mult_generic_AC_RND_CONV_false_5_r_nan_or_nl,
          return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_xnor_nl,
          return_add_generic_AC_RND_CONV_false_24_r_nan_and_nl, {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse
          , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13]) , (fsm_output[14])
          , (fsm_output[21]) , (fsm_output[36]) , (fsm_output[37]) , (fsm_output[38])
          , (fsm_output[39]) , (fsm_output[46])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_do_sub_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_do_sub_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_740 | or_dcpl_224 | (fsm_output[19]) | (fsm_output[22])
        | (fsm_output[20]) | or_dcpl_473 | or_dcpl_702 | (fsm_output[16:15]!=2'b00)
        | or_dcpl_719 | or_dcpl_484)) ) begin
      return_add_generic_AC_RND_CONV_false_12_do_sub_sva <= MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1,
          return_add_generic_AC_RND_CONV_false_12_do_sub_mux1h_1_cse, return_add_generic_AC_RND_CONV_false_6_do_sub_sva_1,
          return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_xnor_nl,
          return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_12_do_sub_mux1h_6_cse,
          return_add_generic_AC_RND_CONV_false_19_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_xnor_nl,
          {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[11]) , (fsm_output[14])
          , (fsm_output[30]) , (fsm_output[32]) , (fsm_output[36]) , (fsm_output[39])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_16_do_sub_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_16_do_sub_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_590 | or_dcpl_588 | or_dcpl_562 | (fsm_output[7])
        | or_dcpl_750 | or_dcpl_511 | (fsm_output[40]) | or_dcpl_553 | or_dcpl_632
        | (fsm_output[12]) | or_dcpl_744)) ) begin
      return_add_generic_AC_RND_CONV_false_16_do_sub_sva <= MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_12_do_sub_mux1h_1_cse,
          return_add_generic_AC_RND_CONV_false_8_do_sub_return_add_generic_AC_RND_CONV_false_8_do_sub_xor_nl,
          return_add_generic_AC_RND_CONV_false_12_do_sub_mux1h_6_cse, return_add_generic_AC_RND_CONV_false_21_do_sub_return_add_generic_AC_RND_CONV_false_21_do_sub_xor_nl,
          {(fsm_output[5]) , (fsm_output[11]) , (fsm_output[30]) , (fsm_output[36])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_763 | or_dcpl_762 | or_dcpl_534 | or_dcpl_236
        | (fsm_output[43]) | (fsm_output[35]) | or_dcpl_686 | (fsm_output[40]) |
        (fsm_output[12]) | (fsm_output[37]))) ) begin
      return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva <= MUX1HOT_s_1_3_2(all_same_out,
          all_same_out_1, leading_sign_57_0_1_0_19_out_2, {return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse
          , return_add_generic_AC_RND_CONV_false_10_r_zero_or_1_nl , (fsm_output[36])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_645 | or_dcpl_686 | or_dcpl_579 | or_dcpl_509
        | or_dcpl_596 | or_dcpl_575 | or_dcpl_744)) ) begin
      return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 <= MUX1HOT_s_1_5_2(return_extract_50_and_nl,
          return_mult_generic_AC_RND_CONV_false_2_zero_m_return_mult_generic_AC_RND_CONV_false_2_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_2_r_zero_return_mult_generic_AC_RND_CONV_false_2_r_zero_nor_nl,
          return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1, return_mult_generic_AC_RND_CONV_false_5_zero_m_return_mult_generic_AC_RND_CONV_false_5_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_5_r_zero_return_mult_generic_AC_RND_CONV_false_5_r_zero_nor_nl,
          return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2, {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse
          , (fsm_output[13]) , (fsm_output[14]) , (fsm_output[38]) , (fsm_output[39])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_21_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_21_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_522 | (fsm_output[21]) | (fsm_output[15]) | or_dcpl_776))
        ) begin
      operator_11_true_return_21_sva <= MUX1HOT_s_1_7_2(operator_11_true_3_operator_11_true_3_and_tmp,
          return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp,
          operator_11_true_53_operator_11_true_53_and_nl, operator_11_true_27_operator_11_true_27_and_nl,
          operator_11_true_35_operator_11_true_35_and_tmp, return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp,
          operator_11_true_59_operator_11_true_59_and_nl, {return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse
          , or_dcpl_208 , return_add_generic_AC_RND_CONV_false_10_ls_or_2_cse , (fsm_output[18])
          , return_add_generic_AC_RND_CONV_false_13_op2_mu_or_5_cse , or_dcpl_235
          , (fsm_output[43])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_24_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_24_sva <= 1'b0;
    end
    else if ( run_wen & ((~(inverse_lpi_1_dfm_1 | or_dcpl_789 | return_add_generic_AC_RND_CONV_false_10_ls_or_2_cse
        | (fsm_output[34]) | or_dcpl_560 | (fsm_output[10]) | return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse
        | (fsm_output[15]) | or_dcpl_580 | or_dcpl_678 | or_dcpl_484)) | (fsm_output[5])
        | (fsm_output[18]) | (fsm_output[32]) | (fsm_output[41])) ) begin
      operator_11_true_return_24_sva <= MUX1HOT_s_1_12_2(return_add_generic_AC_RND_CONV_false_1_if_2_return_add_generic_AC_RND_CONV_false_1_if_2_and_1_mx0w0,
          (stage_PE_1_tmp_re_d_sva[63]), (out_f_d_rsci_q_d[63]), operator_11_true_3_operator_11_true_3_and_tmp,
          return_add_generic_AC_RND_CONV_false_10_if_2_return_add_generic_AC_RND_CONV_false_10_if_2_and_1_mx3w0,
          return_add_generic_AC_RND_CONV_false_17_mux_6_itm, operator_11_true_35_operator_11_true_35_and_tmp,
          return_add_generic_AC_RND_CONV_false_13_if_2_return_add_generic_AC_RND_CONV_false_13_if_2_and_1_mx4w1,
          (in_f_d_rsci_q_d[63]), return_add_generic_AC_RND_CONV_false_9_if_2_return_add_generic_AC_RND_CONV_false_9_if_2_and_1_mx5w0,
          (stage_PE_1_x_re_d_sva[63]), return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1,
          {return_add_generic_AC_RND_CONV_false_12_and_105_cse , return_extract_24_exception_or_1_nl
          , return_add_generic_AC_RND_CONV_false_12_and_116_cse , (fsm_output[7])
          , return_add_generic_AC_RND_CONV_false_12_and_107_cse , return_add_generic_AC_RND_CONV_false_12_and_118_cse
          , return_add_generic_AC_RND_CONV_false_12_and_112_cse , return_add_generic_AC_RND_CONV_false_12_and_109_cse
          , return_add_generic_AC_RND_CONV_false_12_and_110_cse , return_add_generic_AC_RND_CONV_false_12_and_113_cse
          , return_add_generic_AC_RND_CONV_false_12_and_119_cse , return_add_generic_AC_RND_CONV_false_12_and_120_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_21_m_zero_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_21_m_zero_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_789 | (fsm_output[39]) | (fsm_output[38]) | (fsm_output[15])
        | or_dcpl_776)) ) begin
      return_extract_21_m_zero_sva <= MUX1HOT_s_1_7_2(return_extract_3_m_zero_sva_mx1w0,
          return_extract_21_m_zero_return_extract_21_m_zero_nor_nl, return_extract_27_m_zero_return_extract_27_m_zero_nor_nl,
          return_extract_56_m_zero_sva_mx2w0, return_extract_44_m_zero_return_extract_44_m_zero_nor_nl,
          return_extract_52_m_zero_return_extract_52_m_zero_nor_nl, return_extract_57_m_zero_return_extract_57_m_zero_nor_nl,
          {return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse , (fsm_output[14])
          , (fsm_output[18]) , return_add_generic_AC_RND_CONV_false_13_op2_mu_or_5_cse
          , or_dcpl_235 , (fsm_output[37]) , (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_6_false_17_acc_itm_6_1 <= 6'b000000;
    end
    else if ( rst ) begin
      operator_6_false_17_acc_itm_6_1 <= 6'b000000;
    end
    else if ( run_wen & (~(or_dcpl_800 | or_dcpl_209 | or_dcpl_725 | or_dcpl_545
        | or_dcpl_236 | return_add_generic_AC_RND_CONV_false_11_or_4_cse | or_dcpl_680))
        ) begin
      operator_6_false_17_acc_itm_6_1 <= MUX1HOT_v_6_4_2(operator_6_false_17_mux1h_cse_1,
          acc_18_cse_6_1, (drf_qr_lval_21_smx_9_0_lpi_3_dfm[5:0]), rtn_out_2, {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse
          , operator_6_false_17_or_8_cse , operator_6_false_17_and_2_nl , operator_6_false_17_or_9_nl});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_5_1 <= 5'b00000;
      return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_0 <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_5_1 <= 5'b00000;
      return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_0 <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_ssc ) begin
      return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_5_1 <= MUX1HOT_v_5_8_2((operator_6_false_17_mux1h_cse_1[5:1]),
          (operator_14_false_1_acc_psp_sva_9_0[5:1]), (rtn_out_2[5:1]), (drf_qr_lval_6_smx_lpi_3_dfm_mx0_9_1[4:0]),
          (return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1[5:1]), (drf_qr_lval_22_smx_lpi_3_dfm_mx0_9_1[4:0]),
          (leading_sign_57_0_1_0_19_out_3[5:1]), (return_add_generic_AC_RND_CONV_false_24_e_dif_sat_sva_1[5:1]),
          {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_1_cse
          , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_4_cse , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_4_cse
          , (fsm_output[16]) , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_5_cse
          , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_6_cse , (fsm_output[41])});
      return_add_generic_AC_RND_CONV_false_17_e_dif_sat_sva_0 <= MUX1HOT_s_1_8_2((operator_6_false_17_mux1h_cse_1[0]),
          (operator_14_false_1_acc_psp_sva_9_0[0]), (rtn_out_2[0]), drf_qr_lval_6_smx_lpi_3_dfm_mx0_0,
          (return_add_generic_AC_RND_CONV_false_11_e_dif_sat_sva_1[0]), drf_qr_lval_22_smx_lpi_3_dfm_mx0_0,
          (leading_sign_57_0_1_0_19_out_3[0]), (return_add_generic_AC_RND_CONV_false_24_e_dif_sat_sva_1[0]),
          {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_1_cse
          , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_4_cse , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_4_cse
          , (fsm_output[16]) , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_5_cse
          , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_and_6_cse , (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_ls_sva <= 6'b000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_ls_sva <= 6'b000000;
    end
    else if ( run_wen & (~(or_dcpl_809 | or_dcpl_728 | or_dcpl_788 | or_dcpl_493))
        ) begin
      return_add_generic_AC_RND_CONV_false_10_ls_sva <= MUX1HOT_v_6_3_2(rtn_out_1,
          rtn_out_2, rtn_out, {return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse
          , return_add_generic_AC_RND_CONV_false_10_ls_or_6_nl , return_add_generic_AC_RND_CONV_false_10_ls_or_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_32_false_1_acc_psp_sva_11_0 <= 12'b000000000000;
    end
    else if ( rst ) begin
      operator_32_false_1_acc_psp_sva_11_0 <= 12'b000000000000;
    end
    else if ( run_wen & (~(or_dcpl_699 | or_dcpl_509)) ) begin
      operator_32_false_1_acc_psp_sva_11_0 <= MUX1HOT_v_12_4_2((stage_u_add_acc_1_itm_1[11:0]),
          (z_out_64[11:0]), operator_6_false_7_acc_psp_sva_mx0w0, z_out_102, {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse
          , operator_32_false_1_or_1_nl , operator_32_false_1_operator_32_false_1_nor_nl
          , operator_6_false_7_or_rgt});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm
          <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm
          <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_529 | (fsm_output[8]) | or_dcpl_466)) ) begin
      return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm
          <= MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
          return_add_generic_AC_RND_CONV_false_14_mux1h_11_nl, nor_245_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_49_0 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_49_0 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_12_op_bigger_and_cse & (and_2393_rgt
        | and_2395_rgt | and_2185_cse | and_1251_cse | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse
        | and_2407_rgt | and_2409_rgt | and_2184_cse | and_1057_cse | and_1046_cse
        | (~ return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_mx1c2))
        ) begin
      return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_49_0 <= MUX1HOT_v_50_8_2((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_mx1w0[49:0]),
          (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[50:1]), (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[49:0]),
          return_extract_21_mux_cse, return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0,
          (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[49:0]),
          return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49:0]),
          {(~ return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_mx1c2)
          , return_extract_22_or_nl , return_extract_22_or_1_nl , return_extract_22_or_2_cse
          , and_1251_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse
          , and_1057_cse , and_1046_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm
          <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm
          <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~ (fsm_output[38])) ) begin
      return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm
          <= MUX1HOT_v_51_7_2(return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm_mx1w0,
          (return_add_generic_AC_RND_CONV_false_res_rounded_lpi_3_dfm_51_0_1[50:0]),
          return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx1,
          return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1, (return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1[50:0]),
          return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx2,
          return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1, {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse
          , return_add_generic_AC_RND_CONV_false_13_or_cse , or_dcpl_208 , (fsm_output[13])
          , return_add_generic_AC_RND_CONV_false_13_or_3_cse , or_dcpl_235 , (fsm_output[37])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_1 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_2 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_3 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_4 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_5 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_6 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_7 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_8 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_9 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_10 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_11 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_12 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_13 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_14 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_15 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_16 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_17 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_18 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_19 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_20 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_21 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_22 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_23 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_24 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_25 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_26 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_27 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_28 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_29 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_30 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_31 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_32 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_33 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_34 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_35 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_36 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_37 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_38 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_39 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_40 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_41 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_42 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_43 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_44 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_45 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_46 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_47 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_48 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_49 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_50 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_51 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_52 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_53 <= 1'b0;
    end
    else if ( rst ) begin
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_1 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_2 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_3 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_4 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_5 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_6 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_7 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_8 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_9 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_10 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_11 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_12 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_13 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_14 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_15 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_16 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_17 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_18 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_19 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_20 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_21 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_22 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_23 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_24 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_25 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_26 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_27 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_28 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_29 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_30 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_31 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_32 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_33 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_34 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_35 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_36 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_37 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_38 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_39 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_40 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_41 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_42 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_43 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_44 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_45 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_46 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_47 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_48 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_49 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_50 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_51 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_52 <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_53 <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_10_res_rounded_and_cse ) begin
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_1 <= z_out_65[53];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_2 <= z_out_65[52];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_3 <= z_out_65[51];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_4 <= z_out_65[50];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_5 <= z_out_65[49];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_6 <= z_out_65[48];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_7 <= z_out_65[47];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_8 <= z_out_65[46];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_9 <= z_out_65[45];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_10 <= z_out_65[44];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_11 <= z_out_65[43];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_12 <= z_out_65[42];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_13 <= z_out_65[41];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_14 <= z_out_65[40];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_15 <= z_out_65[39];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_16 <= z_out_65[38];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_17 <= z_out_65[37];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_18 <= z_out_65[36];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_19 <= z_out_65[35];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_20 <= z_out_65[34];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_21 <= z_out_65[33];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_22 <= z_out_65[32];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_23 <= z_out_65[31];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_24 <= z_out_65[30];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_25 <= z_out_65[29];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_26 <= z_out_65[28];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_27 <= z_out_65[27];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_28 <= z_out_65[26];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_29 <= z_out_65[25];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_30 <= z_out_65[24];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_31 <= z_out_65[23];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_32 <= z_out_65[22];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_33 <= z_out_65[21];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_34 <= z_out_65[20];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_35 <= z_out_65[19];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_36 <= z_out_65[18];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_37 <= z_out_65[17];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_38 <= z_out_65[16];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_39 <= z_out_65[15];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_40 <= z_out_65[14];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_41 <= z_out_65[13];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_42 <= z_out_65[12];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_43 <= z_out_65[11];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_44 <= z_out_65[10];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_45 <= z_out_65[9];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_46 <= z_out_65[8];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_47 <= z_out_65[7];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_48 <= z_out_65[6];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_49 <= z_out_65[5];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_50 <= z_out_65[4];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_51 <= z_out_65[3];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_52 <= z_out_65[2];
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_53 <= z_out_65[1];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_14_false_1_acc_psp_sva_9_0 <= 10'b0000000000;
    end
    else if ( rst ) begin
      operator_14_false_1_acc_psp_sva_9_0 <= 10'b0000000000;
    end
    else if ( run_wen & (~(or_dcpl_606 | or_dcpl_602 | return_add_generic_AC_RND_CONV_false_12_r_zero_or_1_cse
        | or_dcpl_470 | or_dcpl_598 | or_dcpl_597)) ) begin
      operator_14_false_1_acc_psp_sva_9_0 <= MUX1HOT_v_10_7_2((r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[61:52]),
          (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[61:52]), return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1,
          (stage_PE_1_x_re_d_sva[62:53]), return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1,
          (z_out_86[9:0]), (z_out_68[9:0]), {and_1245_nl , return_add_generic_AC_RND_CONV_false_18_exp_and_2_itm
          , and_1251_cse , or_1302_cse , and_1057_cse , operator_14_false_1_or_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_56 <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_56 <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_12_res_mant_and_ssc & and_dcpl_18
        ) begin
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_56 <= z_out_81[56];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_14_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      drf_qr_lval_14_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_849 | or_dcpl_788 | or_dcpl_470 | or_dcpl_845))
        ) begin
      drf_qr_lval_14_smx_0_lpi_3_dfm <= MUX1HOT_s_1_11_2(return_add_generic_AC_RND_CONV_false_1_r_nan_or_1_nl,
          (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1[51]),
          return_add_generic_AC_RND_CONV_false_2_r_nan_or_1_nl, (return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1[51]),
          return_add_generic_AC_RND_CONV_false_3_r_nan_or_1_nl, (return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1[51]),
          return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_or_nl,
          BUTTERFLY_1_fiy_mux1h_4_cse, return_add_generic_AC_RND_CONV_false_6_r_nan_or_mx6w0,
          return_add_generic_AC_RND_CONV_false_16_r_nan_or_1_nl, BUTTERFLY_1_fiy_mux1h_10_cse,
          {return_add_generic_AC_RND_CONV_false_11_exp_or_nl , return_add_generic_AC_RND_CONV_false_11_exp_or_2_nl
          , return_add_generic_AC_RND_CONV_false_11_exp_and_3_nl , return_add_generic_AC_RND_CONV_false_11_exp_or_3_nl
          , return_add_generic_AC_RND_CONV_false_11_exp_and_5_nl , return_add_generic_AC_RND_CONV_false_11_exp_or_4_nl
          , return_add_generic_AC_RND_CONV_false_10_ls_or_cse , (fsm_output[16])
          , return_add_generic_AC_RND_CONV_false_11_exp_and_9_nl , return_add_generic_AC_RND_CONV_false_11_exp_and_11_nl
          , (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_15_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      drf_qr_lval_15_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_866 | or_dcpl_534 | (fsm_output[23]) | or_dcpl_239
        | or_dcpl_272 | (fsm_output[21]) | or_dcpl_585 | or_dcpl_750 | (fsm_output[8])
        | or_dcpl_466)) ) begin
      drf_qr_lval_15_smx_0_lpi_3_dfm <= MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_5_res_mant_3_0_sva_1,
          (~ return_add_generic_AC_RND_CONV_false_5_res_mant_3_0_sva_1), drf_qr_lval_15_smx_0_lpi_3_dfm_mx2,
          return_add_generic_AC_RND_CONV_false_10_exp_mux1h_3_cse, BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx2,
          return_add_generic_AC_RND_CONV_false_10_exp_mux1h_6_cse, {return_add_generic_AC_RND_CONV_false_12_exp_and_1_nl
          , return_add_generic_AC_RND_CONV_false_12_exp_and_2_nl , (fsm_output[12])
          , (fsm_output[18]) , (fsm_output[38]) , (fsm_output[43])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm
          <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm
          <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_634 | or_dcpl_576)) ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_itm
          <= MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_1_e_r_return_add_generic_AC_RND_CONV_false_1_e_r_or_1_nl,
          return_add_generic_AC_RND_CONV_false_2_e_r_return_add_generic_AC_RND_CONV_false_2_e_r_or_1_nl,
          return_add_generic_AC_RND_CONV_false_3_e_r_return_add_generic_AC_RND_CONV_false_3_e_r_or_1_nl,
          return_add_generic_AC_RND_CONV_false_6_if_5_return_add_generic_AC_RND_CONV_false_6_if_5_and_nl,
          return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_nl,
          return_add_generic_AC_RND_CONV_false_15_e_r_return_add_generic_AC_RND_CONV_false_15_e_r_or_1_nl,
          return_add_generic_AC_RND_CONV_false_16_e_r_return_add_generic_AC_RND_CONV_false_16_e_r_or_1_nl,
          return_add_generic_AC_RND_CONV_false_19_if_5_return_add_generic_AC_RND_CONV_false_19_if_5_and_nl,
          {(fsm_output[6]) , (fsm_output[9]) , (fsm_output[10]) , (fsm_output[11])
          , (fsm_output[31]) , (fsm_output[34]) , (fsm_output[35]) , (fsm_output[36])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_6_false_21_acc_itm_0 <= 1'b0;
    end
    else if ( rst ) begin
      operator_6_false_21_acc_itm_0 <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_876 | or_dcpl_874 | (fsm_output[9]) | (fsm_output[36])
        | (fsm_output[11]) | or_dcpl_870)) ) begin
      operator_6_false_21_acc_itm_0 <= MUX_s_1_2_2((~ (rtn_out_2[0])), return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_or_nl,
          operator_6_false_17_or_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_op2_nan_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_op2_inf_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_op2_nan_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_op2_inf_sva <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_10_op2_nan_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_10_op2_nan_sva <= MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_mx2w0,
          return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0, return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1,
          return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1, {or_tmp_759 , (fsm_output[12])
          , or_tmp_762 , (fsm_output[41])});
      return_add_generic_AC_RND_CONV_false_10_op2_inf_sva <= MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0,
          return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0, return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1,
          return_mult_generic_AC_RND_CONV_false_1_op1_zero_sva_1, {or_tmp_759 , (fsm_output[12])
          , or_tmp_762 , (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_14_op1_nan_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_14_op1_nan_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_621 | or_dcpl_728 | or_dcpl_725 | or_dcpl_236
        | (fsm_output[18]) | or_dcpl_654 | or_dcpl_890)) ) begin
      return_add_generic_AC_RND_CONV_false_14_op1_nan_sva <= MUX1HOT_s_1_9_2(return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0,
          return_mult_generic_AC_RND_CONV_false_op2_inf_sva_1, return_mult_generic_AC_RND_CONV_false_1_op2_inf_sva_1,
          return_mult_generic_AC_RND_CONV_false_2_op2_inf_sva_1, return_add_generic_AC_RND_CONV_false_14_op1_nan_sva_mx0w5,
          return_mult_generic_AC_RND_CONV_false_3_op2_inf_sva_1, return_mult_generic_AC_RND_CONV_false_4_op2_inf_sva_1,
          return_mult_generic_AC_RND_CONV_false_5_op2_inf_sva_1, return_add_generic_AC_RND_CONV_false_10_op1_nan_sva_mx0w9,
          {BUTTERFLY_else_or_cse , (fsm_output[11]) , (fsm_output[12]) , (fsm_output[13])
          , (fsm_output[16]) , (fsm_output[36]) , (fsm_output[37]) , (fsm_output[38])
          , (fsm_output[43])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_866 | or_dcpl_673 | (fsm_output[21]) | (fsm_output[18])
        | or_dcpl_874 | or_dcpl_750 | (fsm_output[38]) | or_dcpl_680 | (fsm_output[8])
        | or_dcpl_466)) ) begin
      return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva <= MUX1HOT_s_1_3_2(all_same_out_1,
          return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1, return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp,
          {return_add_generic_AC_RND_CONV_false_16_r_zero_or_nl , operator_6_false_17_or_cse
          , or_dcpl_484});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_22_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_22_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_800 | or_dcpl_604 | (fsm_output[48]) | or_dcpl_848
        | or_dcpl_671 | or_dcpl_516 | or_dcpl_502 | return_add_generic_AC_RND_CONV_false_11_or_4_cse
        | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[15]) | (fsm_output[40])
        | or_dcpl_492 | (fsm_output[37]))) ) begin
      operator_11_true_return_22_sva <= MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0,
          operator_11_true_54_operator_11_true_54_and_nl, return_extract_58_and_1_nl,
          return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1, {or_1826_nl , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse
          , or_dcpl_625 , (fsm_output[36])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_6_false_21_acc_itm_6_1 <= 6'b000000;
    end
    else if ( rst ) begin
      operator_6_false_21_acc_itm_6_1 <= 6'b000000;
    end
    else if ( run_wen & (~(or_dcpl_876 | or_dcpl_654 | or_dcpl_890)) ) begin
      operator_6_false_21_acc_itm_6_1 <= acc_18_cse_6_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_ls_sva <= 6'b000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_ls_sva <= 6'b000000;
    end
    else if ( run_wen & (~(or_dcpl_928 | or_dcpl_725 | (fsm_output[21]) | (fsm_output[17])
        | return_add_generic_AC_RND_CONV_false_11_or_4_cse | or_dcpl_585 | or_dcpl_269
        | or_dcpl_466)) ) begin
      return_add_generic_AC_RND_CONV_false_11_ls_sva <= rtn_out_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_res_mant_4_sva <= 57'b000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_res_mant_4_sva <= 57'b000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~((fsm_output[45]) | (fsm_output[44]) | (fsm_output[22])
        | (fsm_output[21]) | or_dcpl_470 | or_dcpl_933 | or_dcpl_698 | or_dcpl_680
        | or_dcpl_870)) ) begin
      return_add_generic_AC_RND_CONV_false_11_res_mant_4_sva <= z_out_81;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_1_itm_55_50 <= 6'b000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_1_itm_55_50 <= 6'b000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_18_and_1_ssc & mode_lpi_1_dfm
        ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_1_itm_55_50 <= MUX_v_6_2_2((z_out_74[56:51]),
          (~ (z_out_74[56:51])), return_add_generic_AC_RND_CONV_false_11_do_sub_sva);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_18_and_1_ssc & (and_2325_rgt |
        and_2327_rgt | return_add_generic_AC_RND_CONV_false_13_and_2_cse | return_add_generic_AC_RND_CONV_false_13_and_1_cse
        | and_1251_cse | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse
        | and_2339_rgt | and_2341_rgt | return_add_generic_AC_RND_CONV_false_13_and_4_cse
        | return_add_generic_AC_RND_CONV_false_13_and_3_cse | and_1057_cse | and_1046_cse
        | (~ return_add_generic_AC_RND_CONV_false_18_mux_1_itm_mx1c2)) ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0 <= MUX1HOT_v_50_12_2((z_out_74[50:1]),
          (~ (z_out_74[50:1])), (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx1[49:0]),
          (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx1[50:1]),
          (return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1[50:1]), (return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1[49:0]),
          (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[49:0]),
          return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx2[49:0]),
          (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx2[50:1]),
          (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49:0]),
          return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0, {return_add_generic_AC_RND_CONV_false_18_return_add_generic_AC_RND_CONV_false_18_nor_nl
          , return_add_generic_AC_RND_CONV_false_18_and_9_nl , and_2325_rgt , and_2327_rgt
          , return_add_generic_AC_RND_CONV_false_6_or_nl , return_add_generic_AC_RND_CONV_false_13_or_4_cse
          , and_1251_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse
          , and_2339_rgt , and_2341_rgt , and_1057_cse , and_1046_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_23_op1_mu_52_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_23_op1_mu_52_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_23_op1_mu_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_23_op1_mu_52_lpi_3_dfm <= MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_1, fsm_output[29]);
      return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm <= MUX_v_51_2_2(return_extract_2_mux_4_cse,
          return_extract_33_mux_3_cse, fsm_output[29]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_mux_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_mux_itm <= 1'b0;
    end
    else if ( run_wen & ((~(inverse_lpi_1_dfm_1 | or_dcpl_535 | or_dcpl_726 | or_dcpl_516
        | (fsm_output[18]) | (fsm_output[39]) | or_dcpl_654 | (fsm_output[9]) | or_dcpl_497
        | or_dcpl_970 | (fsm_output[40]) | or_dcpl_509 | (fsm_output[33]) | or_dcpl_640))
        | (fsm_output[7]) | (fsm_output[16]) | (fsm_output[30]) | (fsm_output[43]))
        ) begin
      return_add_generic_AC_RND_CONV_false_11_mux_itm <= MUX1HOT_s_1_13_2(return_add_generic_AC_RND_CONV_false_2_if_2_return_add_generic_AC_RND_CONV_false_2_if_2_nor_1_nl,
          (out_f_d_rsci_q_d[63]), (~ (stage_PE_1_tmp_re_d_sva[63])), return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp,
          return_add_generic_AC_RND_CONV_false_11_if_2_return_add_generic_AC_RND_CONV_false_11_if_2_nor_mx5w0,
          (stage_PE_1_x_re_d_sva[63]), (~ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1),
          return_add_generic_AC_RND_CONV_false_13_if_2_return_add_generic_AC_RND_CONV_false_13_if_2_and_1_mx4w1,
          (stage_PE_1_tmp_re_d_sva[63]), (in_f_d_rsci_q_d[63]), return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp,
          return_add_generic_AC_RND_CONV_false_10_if_2_return_add_generic_AC_RND_CONV_false_10_if_2_and_1_mx3w0,
          return_add_generic_AC_RND_CONV_false_17_mux_6_itm, {and_596_nl , return_add_generic_AC_RND_CONV_false_2_if_2_and_nl
          , return_add_generic_AC_RND_CONV_false_2_if_2_and_1_nl , return_add_generic_AC_RND_CONV_false_11_and_10_cse
          , return_add_generic_AC_RND_CONV_false_11_and_11_cse , return_add_generic_AC_RND_CONV_false_11_and_17_cse
          , return_add_generic_AC_RND_CONV_false_11_and_18_cse , return_add_generic_AC_RND_CONV_false_11_and_13_cse
          , return_add_generic_AC_RND_CONV_false_11_or_9_nl , return_add_generic_AC_RND_CONV_false_11_and_20_cse
          , (fsm_output[32]) , return_add_generic_AC_RND_CONV_false_11_and_15_cse
          , return_add_generic_AC_RND_CONV_false_11_and_22_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_16_mux_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_16_mux_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_800 | or_dcpl_209 | or_dcpl_534 | or_dcpl_470
        | or_dcpl_221 | or_dcpl_466 | (fsm_output[31]))) ) begin
      return_add_generic_AC_RND_CONV_false_16_mux_itm <= MUX1HOT_s_1_10_2(return_add_generic_AC_RND_CONV_false_1_if_2_return_add_generic_AC_RND_CONV_false_1_if_2_and_1_mx0w0,
          (out_f_d_rsci_q_d[63]), (stage_PE_1_tmp_re_d_sva[63]), return_add_generic_AC_RND_CONV_false_9_if_2_return_add_generic_AC_RND_CONV_false_9_if_2_and_1_mx5w0,
          (stage_PE_1_x_re_d_sva[63]), return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_16_if_2_return_add_generic_AC_RND_CONV_false_16_if_2_nor_1_nl,
          (~ (in_f_d_rsci_q_d[63])), return_add_generic_AC_RND_CONV_false_12_if_2_return_add_generic_AC_RND_CONV_false_12_if_2_nor_mx3w0,
          (~ return_add_generic_AC_RND_CONV_false_17_mux_6_itm), {return_add_generic_AC_RND_CONV_false_16_and_1_nl
          , return_add_generic_AC_RND_CONV_false_16_and_9_nl , return_add_generic_AC_RND_CONV_false_16_or_nl
          , return_add_generic_AC_RND_CONV_false_11_and_11_cse , return_add_generic_AC_RND_CONV_false_11_and_17_cse
          , return_add_generic_AC_RND_CONV_false_11_and_18_cse , return_add_generic_AC_RND_CONV_false_11_and_13_cse
          , return_add_generic_AC_RND_CONV_false_11_and_20_cse , return_add_generic_AC_RND_CONV_false_11_and_15_cse
          , return_add_generic_AC_RND_CONV_false_11_and_22_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_20_do_sub_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_20_do_sub_sva <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_10_ls_or_2_cse |
        return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse | or_dcpl_493
        | or_dcpl_484)) ) begin
      return_add_generic_AC_RND_CONV_false_20_do_sub_sva <= MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1,
          return_add_generic_AC_RND_CONV_false_7_do_sub_return_add_generic_AC_RND_CONV_false_7_do_sub_xor_nl,
          return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_20_do_sub_return_add_generic_AC_RND_CONV_false_20_do_sub_xor_nl,
          {(fsm_output[7]) , (fsm_output[11]) , (fsm_output[32]) , (fsm_output[36])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_x_re_d_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      stage_PE_1_x_re_d_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_10_ls_or_2_cse |
        return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse | or_dcpl_497 |
        or_dcpl_970 | or_dcpl_555 | or_dcpl_554)) ) begin
      stage_PE_1_x_re_d_sva <= MUX_v_64_2_2(out_f_d_rsci_q_d, in_f_d_rsci_q_d, fsm_output[32]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_6_false_17_acc_itm_0 <= 1'b0;
    end
    else if ( rst ) begin
      operator_6_false_17_acc_itm_0 <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_11_or_4_cse | (fsm_output[35])
        | (fsm_output[10]) | (fsm_output[12]) | (fsm_output[37]))) ) begin
      operator_6_false_17_acc_itm_0 <= MUX1HOT_s_1_4_2((~ (rtn_out_2[0])), return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_or_1_nl,
          return_add_generic_AC_RND_CONV_false_6_exp_plus_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_19_exp_plus_1_0_lpi_3_dfm_1,
          {operator_6_false_17_or_8_cse , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse
          , (fsm_output[11]) , (fsm_output[36])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_op1_nan_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_op1_nan_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_606 | or_dcpl_602 | or_dcpl_476 | or_dcpl_239
        | or_dcpl_272 | or_dcpl_473 | or_dcpl_484)) ) begin
      return_add_generic_AC_RND_CONV_false_10_op1_nan_sva <= MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_mx2w0,
          return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0, return_add_generic_AC_RND_CONV_false_10_op1_nan_sva_mx0w9,
          return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1, return_add_generic_AC_RND_CONV_false_14_op1_nan_sva_mx0w5,
          {(fsm_output[8]) , or_dcpl_906 , (fsm_output[18]) , (fsm_output[36]) ,
          (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_22_op1_inf_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_22_op1_inf_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_849 | or_dcpl_236 | or_dcpl_625 | or_dcpl_654
        | or_dcpl_466)) ) begin
      return_add_generic_AC_RND_CONV_false_22_op1_inf_sva <= MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0,
          return_extract_56_and_1_nl, return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0,
          {(fsm_output[8]) , return_add_generic_AC_RND_CONV_false_11_or_4_cse , (fsm_output[31])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva <= 57'b000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva <= 57'b000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_809 | or_dcpl_519 | (fsm_output[43]) | or_dcpl_943
        | (fsm_output[10]) | or_dcpl_484)) ) begin
      return_add_generic_AC_RND_CONV_false_10_res_mant_4_sva <= z_out_81;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_33_true_36_acc_psp_1_sva <= 12'b000000000000;
    end
    else if ( rst ) begin
      operator_33_true_36_acc_psp_1_sva <= 12'b000000000000;
    end
    else if ( run_wen & (~((fsm_output[34]) | (fsm_output[10]) | (fsm_output[36])
        | or_dcpl_466)) ) begin
      operator_33_true_36_acc_psp_1_sva <= MUX_v_12_2_2(z_out_102, operator_6_false_7_acc_psp_sva_mx0w0,
          fsm_output[31]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_63 <= 1'b0;
      stage_d_mul_return_d_2_63_sva <= 1'b0;
      stage_d_mul_return_d_4_63_sva <= 1'b0;
    end
    else if ( rst ) begin
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_63 <= 1'b0;
      stage_d_mul_return_d_2_63_sva <= 1'b0;
      stage_d_mul_return_d_4_63_sva <= 1'b0;
    end
    else if ( stage_PE_1_tmp_re_d_and_1_cse ) begin
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_63 <= MUX1HOT_s_1_6_2((out_f_d_rsci_q_d[63]),
          return_add_generic_AC_RND_CONV_false_11_mux_itm, stage_d_mul_return_d_1_63_sva_1,
          (in_f_d_rsci_q_d[63]), return_add_generic_AC_RND_CONV_false_12_mux_itm,
          stage_d_mul_return_d_63_sva_1, {stage_PE_1_tmp_re_d_and_3_nl , stage_PE_1_tmp_re_d_and_4_nl
          , (fsm_output[11]) , stage_PE_1_tmp_re_d_and_5_nl , stage_PE_1_tmp_re_d_and_6_nl
          , (fsm_output[36])});
      stage_d_mul_return_d_2_63_sva <= MUX_s_1_2_2(stage_d_mul_return_d_2_63_sva_1,
          stage_d_mul_return_d_5_63_sva_1, fsm_output[36]);
      stage_d_mul_return_d_4_63_sva <= MUX_s_1_2_2(stage_d_mul_return_d_63_sva_1,
          stage_d_mul_return_d_4_63_sva_2, fsm_output[36]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_r_zero_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_r_zero_1_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_928 | or_dcpl_725 | or_dcpl_545 | or_dcpl_236
        | or_dcpl_588 | (fsm_output[16]) | (fsm_output[36]) | (fsm_output[11])))
        ) begin
      return_add_generic_AC_RND_CONV_false_12_r_zero_1_sva <= all_same_out_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_1_p_1_sva <= 106'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_1_p_1_sva <= 106'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & ((mode_lpi_1_dfm & (~ (z_out_86[12]))) | (mode_lpi_1_dfm
        & (~ (z_out_68[12])))) ) begin
      return_mult_generic_AC_RND_CONV_false_1_p_1_sva <= z_out_104;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_22_m_zero_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_22_m_zero_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_504 | return_add_generic_AC_RND_CONV_false_11_or_4_cse
        | or_dcpl_493)) & mode_lpi_1_dfm ) begin
      return_extract_22_m_zero_sva <= ~(BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx2
          | (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_9_ls_sva <= 6'b000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_9_ls_sva <= 6'b000000;
    end
    else if ( run_wen & (~(or_dcpl_248 | (fsm_output[17]))) ) begin
      return_add_generic_AC_RND_CONV_false_9_ls_sva <= rtn_out_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0 <= 5'b00000;
    end
    else if ( rst ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0 <= 5'b00000;
    end
    else if ( run_wen & (~ return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse)
        ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0 <= MUX1HOT_v_5_3_2((out_u_rsci_q_d[15:11]),
          (z_out_58[15:11]), (in_u_rsci_q_d[15:11]), {return_add_generic_AC_RND_CONV_false_13_or_2_cse
          , or_1341_cse , stage_PE_1_tmp_re_d_or_3_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_0 <= 1'b0;
    end
    else if ( rst ) begin
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_0 <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_7_exp_and_ssc ) begin
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_0 <= MUX1HOT_s_1_11_2((drf_qr_lval_1_smx_lpi_3_dfm_mx0[10]),
          (drf_qr_lval_10_smx_lpi_3_dfm_mx2[10]), (drf_qr_lval_10_smx_lpi_3_dfm_mx3_10_1[9]),
          (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
          (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
          BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0, (return_extract_32_mux_cse[10]),
          (drf_qr_lval_10_smx_lpi_3_dfm_mx6[10]), (drf_qr_lval_10_smx_lpi_3_dfm_mx7_10_1[9]),
          (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
          (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
          {(fsm_output[5]) , (fsm_output[7]) , or_dcpl_208 , (fsm_output[13]) , return_add_generic_AC_RND_CONV_false_7_exp_and_6_nl
          , return_add_generic_AC_RND_CONV_false_7_exp_and_7_nl , (fsm_output[30])
          , (fsm_output[32]) , or_dcpl_235 , (fsm_output[37]) , (fsm_output[39])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_0 <= 4'b0000;
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1 <= 52'b0000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_0 <= 4'b0000;
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1 <= 52'b0000000000000000000000000000000000000000000000000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_12_res_mant_and_1_ssc ) begin
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_0 <= MUX_v_4_2_2((return_add_generic_AC_RND_CONV_false_12_res_mant_mux1h_1_itm[55:52]),
          (z_out_81[55:52]), or_dcpl_534);
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1 <= MUX1HOT_v_52_3_2(and_2619_nl,
          (return_add_generic_AC_RND_CONV_false_12_res_mant_mux1h_1_itm[51:0]), (z_out_81[51:0]),
          {or_1760_nl , or_1761_nl , or_dcpl_534});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0 <= 1'b0;
    end
    else if ( rst ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0 <= 1'b0;
    end
    else if ( and_3925_ssc & ((~ or_1866_ssc) | or_1864_ssc | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
        | return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse | (fsm_output[12])
        | return_extract_22_or_2_cse | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_32_cse
        | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse | (fsm_output[38])
        | return_add_generic_AC_RND_CONV_false_13_or_2_cse | BUTTERFLY_1_else_1_if_and_1_rgt
        | stage_PE_1_tmp_re_d_or_3_cse) ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0 <= MUX1HOT_s_1_11_2((out_u_rsci_q_d[10]),
          (z_out_58[10]), (stage_PE_1_tmp_re_d_sva[62]), (out_f_d_rsci_q_d[62]),
          return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_4_nl,
          (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
          (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
          drf_qr_lval_10_smx_lpi_3_dfm_rsp_0, (in_f_d_rsci_q_d[62]), (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
          (in_u_rsci_q_d[10]), {return_add_generic_AC_RND_CONV_false_13_or_2_cse
          , BUTTERFLY_1_else_1_if_and_1_rgt , BUTTERFLY_1_else_1_if_and_4_nl , BUTTERFLY_1_else_1_if_and_5_nl
          , BUTTERFLY_1_else_1_if_and_6_nl , BUTTERFLY_1_else_1_if_and_7_nl , BUTTERFLY_1_else_1_if_and_8_nl
          , BUTTERFLY_1_else_1_if_and_9_nl , BUTTERFLY_1_else_1_if_and_10_nl , BUTTERFLY_1_else_1_if_and_11_nl
          , stage_PE_1_tmp_re_d_or_3_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1 <= 10'b0000000000;
    end
    else if ( rst ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1 <= 10'b0000000000;
    end
    else if ( and_3925_ssc ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1 <= MUX1HOT_v_10_4_2((out_u_rsci_q_d[9:0]),
          ({BUTTERFLY_1_else_3_else_mux_2_nl , BUTTERFLY_1_else_3_else_mux_3_nl}),
          ({BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_1_9_1 , BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_1_0}),
          (in_u_rsci_q_d[9:0]), {return_add_generic_AC_RND_CONV_false_13_or_2_cse
          , or_1341_cse , or_1342_itm , stage_PE_1_tmp_re_d_or_3_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0 <= 9'b000000000;
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1 <= 1'b0;
    end
    else if ( rst ) begin
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0 <= 9'b000000000;
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1 <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_7_exp_and_2_ssc ) begin
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0 <= MUX1HOT_v_9_13_2((drf_qr_lval_1_smx_lpi_3_dfm_mx0[9:1]),
          (drf_qr_lval_10_smx_lpi_3_dfm_mx2[9:1]), (drf_qr_lval_10_smx_lpi_3_dfm_mx3_10_1[8:0]),
          (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_1[9:1]),
          (return_add_generic_AC_RND_CONV_false_7_exp_mux1h_4_itm_9_0[9:1]), (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1[9:1]),
          (stage_PE_1_tmp_re_d_sva[62:54]), (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[9:1]),
          (return_extract_32_mux_cse[9:1]), (drf_qr_lval_10_smx_lpi_3_dfm_mx6[9:1]),
          (drf_qr_lval_10_smx_lpi_3_dfm_mx7_10_1[8:0]), (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1[9:1]),
          (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[9:1]),
          {(fsm_output[5]) , (fsm_output[7]) , or_dcpl_208 , (fsm_output[13]) , (fsm_output[14])
          , or_tmp_946 , return_add_generic_AC_RND_CONV_false_18_exp_or_cse , or_1993_cse
          , (fsm_output[30]) , (fsm_output[32]) , or_dcpl_235 , (fsm_output[37])
          , (fsm_output[39])});
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1 <= MUX1HOT_s_1_13_2((drf_qr_lval_1_smx_lpi_3_dfm_mx0[0]),
          (drf_qr_lval_10_smx_lpi_3_dfm_mx2[0]), drf_qr_lval_10_smx_lpi_3_dfm_mx3_0,
          (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_1[0]),
          (return_add_generic_AC_RND_CONV_false_7_exp_mux1h_4_itm_9_0[0]), (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1[0]),
          (stage_PE_1_tmp_re_d_sva[53]), (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[0]),
          (return_extract_32_mux_cse[0]), (drf_qr_lval_10_smx_lpi_3_dfm_mx6[0]),
          drf_qr_lval_10_smx_lpi_3_dfm_mx7_0, (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1[0]),
          (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[0]),
          {(fsm_output[5]) , (fsm_output[7]) , or_dcpl_208 , (fsm_output[13]) , (fsm_output[14])
          , or_tmp_946 , return_add_generic_AC_RND_CONV_false_18_exp_or_cse , or_1993_cse
          , (fsm_output[30]) , (fsm_output[32]) , or_dcpl_235 , (fsm_output[37])
          , (fsm_output[39])});
    end
  end
  assign return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl = (~ return_mult_generic_AC_RND_CONV_false_6_e_incr_lpi_2_dfm_2)
      & return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_6_else_2_else_mux_nl = MUX_v_11_2_2((z_out_96[10:0]),
      return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3, return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl);
  assign return_mult_generic_AC_RND_CONV_false_6_else_2_else_return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl
      = MUX_v_11_2_2(11'b00000000000, return_mult_generic_AC_RND_CONV_false_6_else_2_else_mux_nl,
      return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_or_nl
      = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_6_else_2_else_return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_6_lor_lpi_2_dfm_1);
  assign BUTTERFLY_if_1_and_nl = (~ return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1)
      & out1_rsci_idat_63_0_mx0c1;
  assign BUTTERFLY_if_1_and_1_nl = return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1
      & out1_rsci_idat_63_0_mx0c1;
  assign return_mult_generic_AC_RND_CONV_false_6_oelse_3_not_1_nl = ~ return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1;
  assign return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_and_1_nl
      = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000, (z_out_88[50:0]),
      return_mult_generic_AC_RND_CONV_false_6_oelse_3_not_1_nl);
  assign return_add_generic_AC_RND_CONV_false_12_and_93_nl = (~ return_add_generic_AC_RND_CONV_false_16_do_sub_sva)
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_12_and_94_nl = return_add_generic_AC_RND_CONV_false_16_do_sub_sva
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_12_and_101_nl = (~ return_add_generic_AC_RND_CONV_false_16_do_sub_sva)
      & (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_12_and_102_nl = return_add_generic_AC_RND_CONV_false_16_do_sub_sva
      & (fsm_output[39]);
  assign t_in_mux_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_9, t_in_10_0_lpi_1_dfm_1_8,
      and_dcpl_160);
  assign t_in_mux_2_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_8, t_in_10_0_lpi_1_dfm_1_7,
      and_dcpl_160);
  assign t_in_mux_3_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_7, t_in_10_0_lpi_1_dfm_1_6,
      and_dcpl_160);
  assign t_in_mux_4_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_6, t_in_10_0_lpi_1_dfm_1_5,
      and_dcpl_160);
  assign t_in_mux_5_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_5, t_in_10_0_lpi_1_dfm_1_4,
      and_dcpl_160);
  assign t_in_mux_6_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_4, t_in_10_0_lpi_1_dfm_1_3,
      and_dcpl_160);
  assign t_in_mux_7_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_3, t_in_10_0_lpi_1_dfm_1_2,
      and_dcpl_160);
  assign t_in_mux_8_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_2, t_in_10_0_lpi_1_dfm_1_1,
      and_dcpl_160);
  assign t_in_mux_9_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_1, t_in_10_0_lpi_1_dfm_1_0,
      and_dcpl_160);
  assign need_ovf_1_need_ovf_1_and_nl = t_in_10_0_lpi_1_dfm_1_10 & and_dcpl_160;
  assign need_ovf_1_need_ovf_1_and_1_nl = m_in_0_lpi_1_dfm & and_dcpl_160;
  assign m_in_mux_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_13, m_in_15_1_lpi_1_dfm_1_14,
      and_dcpl_160);
  assign m_in_mux_14_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_12, m_in_15_1_lpi_1_dfm_1_13,
      and_dcpl_160);
  assign m_in_mux_13_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_11, m_in_15_1_lpi_1_dfm_1_12,
      and_dcpl_160);
  assign m_in_mux_12_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_10, m_in_15_1_lpi_1_dfm_1_11,
      and_dcpl_160);
  assign m_in_mux_11_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_9, m_in_15_1_lpi_1_dfm_1_10,
      and_dcpl_160);
  assign m_in_mux_10_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_8, m_in_15_1_lpi_1_dfm_1_9,
      and_dcpl_160);
  assign m_in_mux_9_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_7, m_in_15_1_lpi_1_dfm_1_8,
      and_dcpl_160);
  assign m_in_mux_8_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_6, m_in_15_1_lpi_1_dfm_1_7,
      and_dcpl_160);
  assign m_in_mux_7_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_5, m_in_15_1_lpi_1_dfm_1_6,
      and_dcpl_160);
  assign m_in_mux_6_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_4, m_in_15_1_lpi_1_dfm_1_5,
      and_dcpl_160);
  assign m_in_mux_5_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_3, m_in_15_1_lpi_1_dfm_1_4,
      and_dcpl_160);
  assign m_in_mux_4_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_2, m_in_15_1_lpi_1_dfm_1_3,
      and_dcpl_160);
  assign m_in_mux_3_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_1, m_in_15_1_lpi_1_dfm_1_2,
      and_dcpl_160);
  assign m_in_mux_2_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_0, m_in_15_1_lpi_1_dfm_1_1,
      and_dcpl_160);
  assign not_932_nl = ~ (fsm_output[1]);
  assign and_994_nl = stage_PE_1_and_1_tmp & (fsm_output[2]);
  assign and_996_nl = and_6_cse & (fsm_output[2]);
  assign stage_PE_qif_qelse_mux_nl = MUX_s_1_2_2(m_in_0_lpi_1_dfm, m_in_15_1_lpi_1_dfm_1_0,
      mode_lpi_1_dfm);
  assign stage_PE_qif_qelse_mux_1_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_13, m_in_15_1_lpi_1_dfm_1_14,
      mode_lpi_1_dfm);
  assign stage_PE_qif_qelse_mux_14_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_12, m_in_15_1_lpi_1_dfm_1_13,
      mode_lpi_1_dfm);
  assign stage_PE_qif_qelse_mux_13_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_11, m_in_15_1_lpi_1_dfm_1_12,
      mode_lpi_1_dfm);
  assign stage_PE_qif_qelse_mux_12_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_10, m_in_15_1_lpi_1_dfm_1_11,
      mode_lpi_1_dfm);
  assign stage_PE_qif_qelse_mux_11_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_9, m_in_15_1_lpi_1_dfm_1_10,
      mode_lpi_1_dfm);
  assign return_add_generic_AC_RND_CONV_false_3_return_add_generic_AC_RND_CONV_false_3_and_6_nl
      = MUX_v_10_2_2(10'b0000000000, (operator_33_true_32_acc_tmp[10:1]), return_add_generic_AC_RND_CONV_false_16_acc_3_itm_11_1);
  assign or_2741_nl = ((~ inverse_lpi_1_dfm_1) & or_dcpl_198 & nor_174_m1c) | (inverse_lpi_1_dfm_1
      & or_dcpl_198 & nor_174_m1c);
  assign and_2611_nl = (or_dcpl_224 | or_dcpl_476 | (fsm_output[22]) | (fsm_output[20])
      | or_dcpl_473 | or_dcpl_470 | (fsm_output[7]) | (fsm_output[54]) | (fsm_output[53])
      | (fsm_output[8]) | or_dcpl_466) & nor_174_m1c;
  assign or_2742_nl = ((~ (z_out_89[53])) & (fsm_output[9]) & nor_174_m1c) | ((~
      (z_out_89[53])) & (fsm_output[34]) & nor_174_m1c);
  assign BUTTERFLY_else_and_2_nl = (z_out_89[53]) & (fsm_output[9]) & nor_174_m1c;
  assign or_2744_nl = ((fsm_output[10]) & nor_174_m1c) | ((fsm_output[35]) & nor_174_m1c);
  assign and_2613_nl = and_1251_cse & nor_174_m1c;
  assign and_2614_nl = or_1302_cse & nor_174_m1c;
  assign BUTTERFLY_else_and_4_nl = (z_out_89[53]) & (fsm_output[34]) & nor_174_m1c;
  assign and_2616_nl = and_1057_cse & nor_174_m1c;
  assign and_2617_nl = (fsm_output[55]) & nor_174_m1c;
  assign mux1h_nl = MUX1HOT_v_10_12_2(z_out_66, return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0,
      (z_out_85[10:1]), (return_add_generic_AC_RND_CONV_false_2_exp_plus_1_12_1_lpi_3_dfm_1[9:0]),
      (return_add_generic_AC_RND_CONV_false_3_exp_plus_1_12_1_lpi_3_dfm_1[9:0]),
      return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1, (stage_PE_1_x_re_d_sva[62:53]),
      (return_add_generic_AC_RND_CONV_false_15_exp_plus_1_12_1_lpi_3_dfm_1[9:0]),
      return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1, (z_out_113[9:0]),
      return_add_generic_AC_RND_CONV_false_1_e_r_qelse_qr_10_1_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_3_return_add_generic_AC_RND_CONV_false_3_and_6_nl,
      {or_2741_nl , and_2611_nl , or_2742_nl , BUTTERFLY_else_and_2_nl , or_2744_nl
      , and_2613_nl , and_2614_nl , BUTTERFLY_else_and_4_nl , and_2616_nl , and_2617_nl
      , or_tmp , or_tmp_956});
  assign nand_153_nl = ~(BUTTERFLY_else_or_cse & nor_174_m1c);
  assign and_2618_nl = mux1h_nl & (signext_10_1(nand_153_nl)) & (signext_10_1(~ or_tmp_955));
  assign or_2026_nl = MUX_v_10_2_2(and_2618_nl, 10'b1111111111, or_tmp_954);
  assign and_1068_nl = and_dcpl_393 & (~((fsm_output[45]) | (fsm_output[26]))) &
      and_dcpl_323 & and_dcpl_389 & (~((fsm_output[49]) | (fsm_output[46]))) & (~((fsm_output[48])
      | (fsm_output[4]) | (fsm_output[29]))) & and_dcpl_382 & (~((fsm_output[14])
      | (fsm_output[39]))) & (~((fsm_output[13]) | (fsm_output[38]) | (fsm_output[15])))
      & (~((fsm_output[30]) | (fsm_output[36]))) & (~((fsm_output[40]) | (fsm_output[11])))
      & (~((fsm_output[5]) | (fsm_output[12]) | (fsm_output[37])));
  assign operator_33_true_12_or_1_nl = or_dcpl_493 | or_dcpl_485 | (fsm_output[19])
      | (fsm_output[21]) | (fsm_output[23]) | (fsm_output[25]) | (fsm_output[44])
      | (fsm_output[46]) | (fsm_output[48]) | (fsm_output[50]);
  assign BUTTERFLY_i_or_nl = or_dcpl_485 | BUTTERFLY_1_i_9_0_sva_mx0c3;
  assign return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_3_nl
      = BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx5 | return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp;
  assign return_extract_12_m_zero_return_extract_12_m_zero_nor_nl = ~(stage_PE_tmp_re_d_1_lpi_3_dfm_51_mx0
      | stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50 | (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx1[49:0]!=50'b00000000000000000000000000000000000000000000000000));
  assign return_extract_20_m_zero_return_extract_20_m_zero_nor_nl = ~(drf_qr_lval_15_smx_0_lpi_3_dfm_mx2
      | (return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_25_m_zero_return_extract_25_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_53_m_zero_return_extract_53_m_zero_nor_nl = ~(return_mult_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_mx1
      | (return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_59_m_zero_return_extract_59_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_21_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign operator_11_true_12_operator_11_true_12_and_nl = (drf_qr_lval_10_smx_lpi_3_dfm_mx3_10_1==10'b1111111111)
      & drf_qr_lval_10_smx_lpi_3_dfm_mx3_0;
  assign operator_11_true_52_operator_11_true_52_and_nl = (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1==11'b11111111111);
  assign operator_11_true_25_operator_11_true_25_and_nl = (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1;
  assign operator_11_true_44_operator_11_true_44_and_nl = (drf_qr_lval_10_smx_lpi_3_dfm_mx7_10_1==10'b1111111111)
      & drf_qr_lval_10_smx_lpi_3_dfm_mx7_0;
  assign operator_11_true_57_operator_11_true_57_and_nl = (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_25_r_nan_and_nl = operator_11_true_return_22_sva
      & operator_11_true_return_26_sva & return_add_generic_AC_RND_CONV_false_12_do_sub_sva;
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_or_6_nl = (fsm_output[4])
      | return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse;
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_and_2_nl = (~ and_517_tmp)
      & (fsm_output[6]);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_and_3_nl = and_517_tmp &
      (fsm_output[6]);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_or_8_nl = (fsm_output[29])
      | return_add_generic_AC_RND_CONV_false_13_op2_mu_or_5_cse;
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_and_4_nl = (~ return_extract_33_or_1_tmp)
      & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_and_5_nl = return_extract_33_or_1_tmp
      & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_or_3_nl = and_dcpl_448 |
      (~ inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_or_4_nl = (~ inverse_lpi_1_dfm_1)
      | (z_out_69[11]) | return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_and_1_cse;
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_nor_1_nl = ~((return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_or_1_tmp
      & (~ inverse_lpi_1_dfm_1)) | return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx8c1
      | return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx8c2);
  assign reg_return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_rgt_nl
      = MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_13_op2_mu_or_3_nl, (~
      inverse_lpi_1_dfm_1), return_add_generic_AC_RND_CONV_false_13_op2_mu_or_4_nl,
      and_dcpl_452, return_add_generic_AC_RND_CONV_false_13_op2_mu_nor_1_nl, {(fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[30]) , (fsm_output[32])});
  assign return_add_generic_AC_RND_CONV_false_18_exp_and_1_nl = (~ and_dcpl_460)
      & return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse;
  assign return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_2_nl
      = BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx2 | return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_21_nl = (~ return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp)
      & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_22_nl = return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp
      & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_16_nl = ((~ and_dcpl_467)
      & (fsm_output[14])) | ((~ and_dcpl_469) & (fsm_output[39]));
  assign return_add_generic_AC_RND_CONV_false_11_or_nl = ((~ return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1)
      & return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse) | ((~ return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1)
      & return_add_generic_AC_RND_CONV_false_11_or_5_cse);
  assign return_add_generic_AC_RND_CONV_false_11_or_6_nl = (return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1
      & return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse) | return_add_generic_AC_RND_CONV_false_11_and_9_itm;
  assign return_add_generic_AC_RND_CONV_false_11_or_7_nl = ((~ return_add_generic_AC_RND_CONV_false_16_do_sub_sva)
      & return_add_generic_AC_RND_CONV_false_10_ls_or_2_cse) | ((~ return_add_generic_AC_RND_CONV_false_11_do_sub_sva)
      & return_add_generic_AC_RND_CONV_false_11_or_4_cse);
  assign return_add_generic_AC_RND_CONV_false_11_or_8_nl = (return_add_generic_AC_RND_CONV_false_16_do_sub_sva
      & return_add_generic_AC_RND_CONV_false_10_ls_or_2_cse) | (return_add_generic_AC_RND_CONV_false_11_do_sub_sva
      & return_add_generic_AC_RND_CONV_false_11_or_4_cse);
  assign return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_3_nl
      = drf_qr_lval_15_smx_0_lpi_3_dfm_mx2 | return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp;
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_or_nl = or_dcpl_485 |
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx0c8;
  assign return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_and_2_nl
      = MUX_v_11_2_2(11'b00000000000, z_out_112, return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1);
  assign return_add_generic_AC_RND_CONV_false_4_if_2_return_add_generic_AC_RND_CONV_false_4_if_2_nor_1_nl
      = ~(inverse_lpi_1_dfm_1 | (~ (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[63])));
  assign or_756_nl = (fsm_output[12:11]!=2'b00);
  assign or_1538_nl = (fsm_output[37:36]!=2'b00);
  assign return_add_generic_AC_RND_CONV_false_5_if_2_return_add_generic_AC_RND_CONV_false_5_if_2_and_2_nl
      = inverse_lpi_1_dfm_1 & (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[63]);
  assign return_add_generic_AC_RND_CONV_false_9_do_sub_return_add_generic_AC_RND_CONV_false_9_do_sub_xor_nl
      = (stage_PE_1_x_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1;
  assign return_add_generic_AC_RND_CONV_false_23_do_sub_return_add_generic_AC_RND_CONV_false_23_do_sub_xor_nl
      = (stage_PE_1_tmp_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_17_mux_6_itm_mx4;
  assign return_add_generic_AC_RND_CONV_false_3_if_2_return_add_generic_AC_RND_CONV_false_3_if_2_nor_1_nl
      = ~((out_f_d_rsci_q_d[63]) | (~ (stage_PE_1_tmp_re_d_sva[63])));
  assign return_add_generic_AC_RND_CONV_false_15_if_2_return_add_generic_AC_RND_CONV_false_15_if_2_nor_1_nl
      = ~((stage_PE_1_tmp_re_d_sva[63]) | (~ (in_f_d_rsci_q_d[63])));
  assign return_add_generic_AC_RND_CONV_false_12_or_46_nl = return_add_generic_AC_RND_CONV_false_12_and_115_cse
      | return_add_generic_AC_RND_CONV_false_12_and_117_cse;
  assign return_add_generic_AC_RND_CONV_false_17_do_sub_return_add_generic_AC_RND_CONV_false_17_do_sub_return_add_generic_AC_RND_CONV_false_17_do_sub_xnor_nl
      = ~((BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[63]) ^ inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_10_do_sub_return_add_generic_AC_RND_CONV_false_10_do_sub_xor_nl
      = (stage_PE_1_tmp_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_17_mux_6_itm_mx2;
  assign return_add_generic_AC_RND_CONV_false_22_do_sub_return_add_generic_AC_RND_CONV_false_22_do_sub_xor_nl
      = (stage_PE_1_x_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2;
  assign return_add_generic_AC_RND_CONV_false_18_do_sub_return_add_generic_AC_RND_CONV_false_18_do_sub_xor_nl
      = (BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out[63]) ^ inverse_lpi_1_dfm_1;
  assign return_mult_generic_AC_RND_CONV_false_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0
      | (operator_11_true_15_operator_11_true_15_and_tmp & (~ return_extract_47_m_zero_return_extract_47_m_zero_nor_tmp))
      | (return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0 & return_mult_generic_AC_RND_CONV_false_op2_zero_sva_1)
      | (return_mult_generic_AC_RND_CONV_false_1_op1_zero_sva_1 & return_mult_generic_AC_RND_CONV_false_op2_inf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_1_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0
      | (operator_11_true_17_operator_11_true_17_and_tmp & (~ return_extract_49_m_zero_return_extract_49_m_zero_nor_tmp))
      | (return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0 & return_mult_generic_AC_RND_CONV_false_1_op2_zero_sva_1)
      | (return_mult_generic_AC_RND_CONV_false_1_op1_zero_sva_1 & return_mult_generic_AC_RND_CONV_false_1_op2_inf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_2_r_nan_or_nl = (operator_11_true_19_operator_11_true_19_and_tmp
      & (~ return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp)) | (return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1
      & return_mult_generic_AC_RND_CONV_false_2_op2_inf_sva_1);
  assign return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_xnor_nl
      = ~((stage_PE_1_x_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1);
  assign return_add_generic_AC_RND_CONV_false_11_r_nan_and_nl = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      & operator_11_true_return_26_sva & return_add_generic_AC_RND_CONV_false_11_do_sub_sva;
  assign return_mult_generic_AC_RND_CONV_false_3_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1
      | (operator_11_true_47_operator_11_true_47_and_tmp & (~ return_extract_47_m_zero_return_extract_47_m_zero_nor_tmp))
      | (return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1 & return_mult_generic_AC_RND_CONV_false_3_op2_zero_sva_1)
      | (return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0 & return_mult_generic_AC_RND_CONV_false_3_op2_inf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_4_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1
      | (operator_11_true_49_operator_11_true_49_and_tmp & (~ return_extract_49_m_zero_return_extract_49_m_zero_nor_tmp))
      | (return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1 & return_mult_generic_AC_RND_CONV_false_4_op2_zero_sva_1)
      | (return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0 & return_mult_generic_AC_RND_CONV_false_4_op2_inf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_5_r_nan_or_nl = (operator_11_true_51_operator_11_true_51_and_tmp
      & (~ return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp)) | (return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1
      & return_mult_generic_AC_RND_CONV_false_5_op2_inf_sva_1);
  assign return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_xnor_nl
      = ~((stage_PE_1_x_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2);
  assign return_add_generic_AC_RND_CONV_false_24_r_nan_and_nl = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva & return_add_generic_AC_RND_CONV_false_11_do_sub_sva;
  assign return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_xnor_nl
      = ~((stage_PE_1_tmp_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_17_mux_6_itm_mx2);
  assign return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_xnor_nl
      = ~((stage_PE_1_tmp_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_17_mux_6_itm_mx4);
  assign return_add_generic_AC_RND_CONV_false_8_do_sub_return_add_generic_AC_RND_CONV_false_8_do_sub_xor_nl
      = stage_d_mul_return_d_1_63_sva_1 ^ stage_d_mul_return_d_2_63_sva_1;
  assign return_add_generic_AC_RND_CONV_false_21_do_sub_return_add_generic_AC_RND_CONV_false_21_do_sub_xor_nl
      = stage_d_mul_return_d_4_63_sva_2 ^ stage_d_mul_return_d_5_63_sva_1;
  assign return_add_generic_AC_RND_CONV_false_10_r_zero_or_1_nl = or_dcpl_553 | return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse
      | (fsm_output[11]) | (fsm_output[14]) | (fsm_output[39]) | return_add_generic_AC_RND_CONV_false_10_r_zero_or_3_cse;
  assign return_extract_50_and_nl = return_add_generic_AC_RND_CONV_false_17_return_add_generic_AC_RND_CONV_false_17_if_1_return_add_generic_AC_RND_CONV_false_17_op2_normal_return_extract_41_nor_tmp
      & (r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out[51:0]==52'b0000000000000000000000000000000000000000000000000000);
  assign return_mult_generic_AC_RND_CONV_false_2_zero_m_return_mult_generic_AC_RND_CONV_false_2_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_2_r_zero_return_mult_generic_AC_RND_CONV_false_2_r_zero_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 | return_extract_19_and_cse);
  assign return_mult_generic_AC_RND_CONV_false_5_zero_m_return_mult_generic_AC_RND_CONV_false_5_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_5_r_zero_return_mult_generic_AC_RND_CONV_false_5_r_zero_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 | return_extract_51_and_cse);
  assign operator_11_true_53_operator_11_true_53_and_nl = (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1==11'b11111111111);
  assign operator_11_true_27_operator_11_true_27_and_nl = (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1;
  assign operator_11_true_59_operator_11_true_59_and_nl = (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1;
  assign return_extract_24_exception_or_1_nl = return_add_generic_AC_RND_CONV_false_12_and_115_cse
      | return_add_generic_AC_RND_CONV_false_12_and_117_cse | return_add_generic_AC_RND_CONV_false_12_and_111_cse;
  assign return_extract_21_m_zero_return_extract_21_m_zero_nor_nl = ~(return_mult_generic_AC_RND_CONV_false_2_m_r_51_lpi_3_dfm_mx1
      | (return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_27_m_zero_return_extract_27_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_8_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_44_m_zero_return_extract_44_m_zero_nor_nl = ~(stage_PE_1_tmp_im_d_1_lpi_3_dfm_51_mx1
      | stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50 | (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx2[49:0]!=50'b00000000000000000000000000000000000000000000000000));
  assign return_extract_52_m_zero_return_extract_52_m_zero_nor_nl = ~(BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx5
      | (return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_57_m_zero_return_extract_57_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign operator_6_false_17_and_2_nl = (~ return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1)
      & operator_6_false_17_or_cse;
  assign operator_6_false_17_or_9_nl = (return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1
      & operator_6_false_17_or_cse) | or_dcpl_534;
  assign return_add_generic_AC_RND_CONV_false_10_ls_or_6_nl = or_dcpl_553 | return_add_generic_AC_RND_CONV_false_10_ls_or_2_cse
      | return_add_generic_AC_RND_CONV_false_10_r_zero_or_3_cse;
  assign operator_32_false_1_or_1_nl = ((~ mode_lpi_1_dfm) & (fsm_output[6])) | (fsm_output[31]);
  assign operator_32_false_1_operator_32_false_1_nor_nl = ~(operator_6_false_7_or_rgt
      | (~((mode_lpi_1_dfm & (fsm_output[6])) | or_dcpl_645 | or_dcpl_208 | (fsm_output[8]))));
  assign return_add_generic_AC_RND_CONV_false_14_or_5_nl = (fsm_output[9]) | (fsm_output[10])
      | (fsm_output[34]) | (fsm_output[35]);
  assign return_add_generic_AC_RND_CONV_false_14_mux1h_11_nl = MUX1HOT_v_51_5_2(return_add_generic_AC_RND_CONV_false_14_return_add_generic_AC_RND_CONV_false_14_and_6_itm_mx1w0,
      (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1[50:0]),
      (return_add_generic_AC_RND_CONV_false_2_res_rounded_lpi_3_dfm_51_0_1[50:0]),
      return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1, return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1,
      {return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse , BUTTERFLY_else_or_cse
      , return_add_generic_AC_RND_CONV_false_14_or_5_nl , (fsm_output[12]) , (fsm_output[38])});
  assign nor_245_nl = ~(((return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva |
      return_add_generic_AC_RND_CONV_false_14_exception_sva_1) & (fsm_output[31]))
      | ((return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva | return_add_generic_AC_RND_CONV_false_16_exception_sva_1)
      & (fsm_output[35])) | ((return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva
      | return_add_generic_AC_RND_CONV_false_2_exception_sva_1) & (fsm_output[9]))
      | ((return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva | return_add_generic_AC_RND_CONV_false_1_exception_sva_1)
      & (fsm_output[6])) | ((return_add_generic_AC_RND_CONV_false_3_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_16_r_zero_1_sva) & (fsm_output[10]))
      | ((return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva | return_add_generic_AC_RND_CONV_false_15_exception_sva_1)
      & (fsm_output[34])));
  assign return_extract_22_or_nl = and_2393_rgt | and_2407_rgt;
  assign return_extract_22_or_1_nl = and_2395_rgt | and_2409_rgt;
  assign and_1245_nl = or_658_cse & return_add_generic_AC_RND_CONV_false_18_exp_or_1_cse;
  assign return_add_generic_AC_RND_CONV_false_1_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_mx1w0
      | return_add_generic_AC_RND_CONV_false_7_op2_nan_sva_mx2w0 | (return_add_generic_AC_RND_CONV_false_op2_inf_sva_mx1w0
      & return_add_generic_AC_RND_CONV_false_7_op2_inf_sva_mx2w0 & return_add_generic_AC_RND_CONV_false_12_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_2_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_unequal_tmp | (return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      & operator_11_true_return_26_sva & return_add_generic_AC_RND_CONV_false_12_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_3_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | (operator_11_true_return_22_sva
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva & return_add_generic_AC_RND_CONV_false_16_do_sub_sva);
  assign return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_or_nl
      = ((z_out_104[105]) & (~ (z_out_107[52]))) | ((z_out_104[104]) & (~ (z_out_107[51])))
      | ((z_out_104[103]) & (~ (z_out_107[50]))) | ((z_out_104[102]) & (~ (z_out_107[49])))
      | ((z_out_104[101]) & (~ (z_out_107[48]))) | ((z_out_104[100]) & (~ (z_out_107[47])))
      | ((z_out_104[99]) & (~ (z_out_107[46]))) | ((z_out_104[98]) & (~ (z_out_107[45])))
      | ((z_out_104[97]) & (~ (z_out_107[44]))) | ((z_out_104[96]) & (~ (z_out_107[43])))
      | ((z_out_104[95]) & (~ (z_out_107[42]))) | ((z_out_104[94]) & (~ (z_out_107[41])))
      | ((z_out_104[93]) & (~ (z_out_107[40]))) | ((z_out_104[92]) & (~ (z_out_107[39])))
      | ((z_out_104[91]) & (~ (z_out_107[38]))) | ((z_out_104[90]) & (~ (z_out_107[37])))
      | ((z_out_104[89]) & (~ (z_out_107[36]))) | ((z_out_104[88]) & (~ (z_out_107[35])))
      | ((z_out_104[87]) & (~ (z_out_107[34]))) | ((z_out_104[86]) & (~ (z_out_107[33])))
      | ((z_out_104[85]) & (~ (z_out_107[32]))) | ((z_out_104[84]) & (~ (z_out_107[31])))
      | ((z_out_104[83]) & (~ (z_out_107[30]))) | ((z_out_104[82]) & (~ (z_out_107[29])))
      | ((z_out_104[81]) & (~ (z_out_107[28]))) | ((z_out_104[80]) & (~ (z_out_107[27])))
      | ((z_out_104[79]) & (~ (z_out_107[26]))) | ((z_out_104[78]) & (~ (z_out_107[25])))
      | ((z_out_104[77]) & (~ (z_out_107[24]))) | ((z_out_104[76]) & (~ (z_out_107[23])))
      | ((z_out_104[75]) & (~ (z_out_107[22]))) | ((z_out_104[74]) & (~ (z_out_107[21])))
      | ((z_out_104[73]) & (~ (z_out_107[20]))) | ((z_out_104[72]) & (~ (z_out_107[19])))
      | ((z_out_104[71]) & (~ (z_out_107[18]))) | ((z_out_104[70]) & (~ (z_out_107[17])))
      | ((z_out_104[69]) & (~ (z_out_107[16]))) | ((z_out_104[68]) & (~ (z_out_107[15])))
      | ((z_out_104[67]) & (~ (z_out_107[14]))) | ((z_out_104[66]) & (~ (z_out_107[13])))
      | ((z_out_104[65]) & (~ (z_out_107[12]))) | ((z_out_104[64]) & (~ (z_out_107[11])))
      | ((z_out_104[63]) & (~ (z_out_107[10]))) | ((z_out_104[62]) & (~ (z_out_107[9])))
      | ((z_out_104[61]) & (~ (z_out_107[8]))) | ((z_out_104[60]) & (~ (z_out_107[7])))
      | ((z_out_104[59]) & (~ (z_out_107[6]))) | ((z_out_104[58]) & (~ (z_out_107[5])))
      | ((z_out_104[57]) & (~ (z_out_107[4]))) | ((z_out_104[56]) & (~ (z_out_107[3])))
      | ((z_out_104[55]) & (~ (z_out_107[2]))) | ((z_out_104[54]) & (~ (z_out_107[1])))
      | ((z_out_104[53]) & (~ (z_out_107[0]))) | (z_out_104[52:0]!=53'b00000000000000000000000000000000000000000000000000000);
  assign return_add_generic_AC_RND_CONV_false_16_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_unequal_tmp | (return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      & operator_11_true_return_26_sva & return_add_generic_AC_RND_CONV_false_16_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_11_exp_or_nl = ((~ and_572_tmp) & (fsm_output[6]))
      | ((~ and_584_tmp) & (fsm_output[31]));
  assign return_add_generic_AC_RND_CONV_false_11_exp_or_2_nl = (and_572_tmp & (fsm_output[6]))
      | (and_584_tmp & (fsm_output[31]));
  assign return_add_generic_AC_RND_CONV_false_11_exp_and_3_nl = (~ and_577_tmp) &
      (fsm_output[9]);
  assign return_add_generic_AC_RND_CONV_false_11_exp_or_3_nl = (and_577_tmp & (fsm_output[9]))
      | (and_588_tmp & (fsm_output[34]));
  assign return_add_generic_AC_RND_CONV_false_11_exp_and_5_nl = (~ and_582_tmp) &
      (fsm_output[10]);
  assign return_add_generic_AC_RND_CONV_false_11_exp_or_4_nl = (and_582_tmp & (fsm_output[10]))
      | (and_591_tmp & (fsm_output[35]));
  assign return_add_generic_AC_RND_CONV_false_11_exp_and_9_nl = (~ and_588_tmp) &
      (fsm_output[34]);
  assign return_add_generic_AC_RND_CONV_false_11_exp_and_11_nl = (~ and_591_tmp)
      & (fsm_output[35]);
  assign return_add_generic_AC_RND_CONV_false_12_exp_and_1_nl = (~ return_add_generic_AC_RND_CONV_false_11_do_sub_sva)
      & BUTTERFLY_else_or_cse;
  assign return_add_generic_AC_RND_CONV_false_12_exp_and_2_nl = return_add_generic_AC_RND_CONV_false_11_do_sub_sva
      & BUTTERFLY_else_or_cse;
  assign or_352_nl = and_276_cse | operator_11_true_return_1_sva | or_dcpl_285;
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs, or_352_nl);
  assign return_add_generic_AC_RND_CONV_false_1_e_r_return_add_generic_AC_RND_CONV_false_1_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_30 & (~ return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_nl))
      | return_add_generic_AC_RND_CONV_false_1_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_and_2_nl
      = (z_out_85[0]) & return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_2_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_and_2_nl,
      return_add_generic_AC_RND_CONV_false_2_exp_plus_1_0_lpi_3_dfm_1, z_out_89[53]);
  assign or_370_nl = or_dcpl_301 | and_dcpl_216 | return_add_generic_AC_RND_CONV_false_2_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva;
  assign return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs, or_370_nl);
  assign return_add_generic_AC_RND_CONV_false_2_e_r_return_add_generic_AC_RND_CONV_false_2_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_2_mux_13_nl & (~ return_add_generic_AC_RND_CONV_false_2_e_r_qelse_mux_1_nl))
      | return_add_generic_AC_RND_CONV_false_2_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_3_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_3_return_add_generic_AC_RND_CONV_false_3_and_9,
      return_add_generic_AC_RND_CONV_false_3_exp_plus_1_0_lpi_3_dfm_1, z_out_89[53]);
  assign or_382_nl = return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2 | or_dcpl_311
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_14_op1_nan_sva
      | and_dcpl_217;
  assign return_add_generic_AC_RND_CONV_false_16_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs, or_382_nl);
  assign return_add_generic_AC_RND_CONV_false_3_e_r_return_add_generic_AC_RND_CONV_false_3_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_3_mux_13_nl & (~ return_add_generic_AC_RND_CONV_false_16_e_r_qelse_mux_1_nl))
      | return_add_generic_AC_RND_CONV_false_3_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_6_if_5_return_add_generic_AC_RND_CONV_false_6_if_5_and_nl
      = (return_add_generic_AC_RND_CONV_false_6_exp_plus_1_12_1_lpi_3_dfm_1[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_6_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_6_exp_plus_1_12_1_lpi_3_dfm_1[11:10]==2'b00);
  assign or_409_nl = and_311_cse | operator_11_true_return_1_sva | or_dcpl_285;
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_4_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs_mx0w1,
      return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs, or_409_nl);
  assign return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_30 & (~ return_add_generic_AC_RND_CONV_false_e_r_qelse_mux_4_nl))
      | return_add_generic_AC_RND_CONV_false_14_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_15_return_add_generic_AC_RND_CONV_false_15_and_2_nl
      = (z_out_85[0]) & return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1;
  assign return_add_generic_AC_RND_CONV_false_15_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_15_return_add_generic_AC_RND_CONV_false_15_and_2_nl,
      return_add_generic_AC_RND_CONV_false_15_exp_plus_1_0_lpi_3_dfm_1, z_out_89[53]);
  assign or_426_nl = return_add_generic_AC_RND_CONV_false_15_r_inf_lpi_3_dfm_2 |
      or_dcpl_311 | and_dcpl_251 | or_dcpl_359;
  assign return_add_generic_AC_RND_CONV_false_15_e_r_qelse_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs, or_426_nl);
  assign return_add_generic_AC_RND_CONV_false_15_e_r_return_add_generic_AC_RND_CONV_false_15_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_15_mux_13_nl & (~ return_add_generic_AC_RND_CONV_false_15_e_r_qelse_mux_1_nl))
      | return_add_generic_AC_RND_CONV_false_15_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_16_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_3_return_add_generic_AC_RND_CONV_false_3_and_9,
      return_add_generic_AC_RND_CONV_false_16_exp_plus_1_0_lpi_3_dfm_1, z_out_89[53]);
  assign or_434_nl = return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2 | or_dcpl_93
      | or_dcpl_367 | and_dcpl_253;
  assign return_add_generic_AC_RND_CONV_false_16_e_r_qelse_mux_3_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs_mx0w0,
      return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs, or_434_nl);
  assign return_add_generic_AC_RND_CONV_false_16_e_r_return_add_generic_AC_RND_CONV_false_16_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_16_mux_13_nl & (~ return_add_generic_AC_RND_CONV_false_16_e_r_qelse_mux_3_nl))
      | return_add_generic_AC_RND_CONV_false_16_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_19_if_5_return_add_generic_AC_RND_CONV_false_19_if_5_and_nl
      = (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_2[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_19_exp_plus_1_0_lpi_3_dfm_1 & (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_2[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_5_return_add_generic_AC_RND_CONV_false_5_or_nl
      = (operator_6_false_11_acc_psp_1_sva_1[0]) | (~ return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1);
  assign return_add_generic_AC_RND_CONV_false_16_r_zero_or_nl = BUTTERFLY_else_or_cse
      | (fsm_output[16]) | (fsm_output[20]) | (fsm_output[44]);
  assign operator_11_true_54_operator_11_true_54_and_nl = (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_1==11'b11111111111);
  assign return_extract_58_and_1_nl = operator_11_true_return_26_sva & return_extract_26_m_zero_sva;
  assign or_1826_nl = or_dcpl_906 | (fsm_output[6]);
  assign return_add_generic_AC_RND_CONV_false_18_return_add_generic_AC_RND_CONV_false_18_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_11_do_sub_sva | return_add_generic_AC_RND_CONV_false_18_mux_1_itm_mx1c2);
  assign return_add_generic_AC_RND_CONV_false_18_and_9_nl = return_add_generic_AC_RND_CONV_false_11_do_sub_sva
      & (~ return_add_generic_AC_RND_CONV_false_18_mux_1_itm_mx1c2);
  assign return_add_generic_AC_RND_CONV_false_6_or_nl = return_add_generic_AC_RND_CONV_false_13_and_2_cse
      | return_add_generic_AC_RND_CONV_false_13_and_4_cse;
  assign return_add_generic_AC_RND_CONV_false_2_if_2_return_add_generic_AC_RND_CONV_false_2_if_2_nor_1_nl
      = ~((stage_PE_1_tmp_re_d_sva[63]) | (~ (out_f_d_rsci_q_d[63])));
  assign and_596_nl = inverse_lpi_1_dfm_1 & return_add_generic_AC_RND_CONV_false_e1_eq_e2_equal_tmp
      & return_add_generic_AC_RND_CONV_false_2_aif_equal_tmp & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_2_if_2_and_nl = (~ return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse)
      & and_597_m1c & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_2_if_2_and_1_nl = return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse
      & and_597_m1c & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_11_or_9_nl = return_add_generic_AC_RND_CONV_false_11_and_19_cse
      | return_add_generic_AC_RND_CONV_false_11_and_21_cse;
  assign return_add_generic_AC_RND_CONV_false_16_if_2_return_add_generic_AC_RND_CONV_false_16_if_2_nor_1_nl
      = ~((in_f_d_rsci_q_d[63]) | (~ (stage_PE_1_tmp_re_d_sva[63])));
  assign return_add_generic_AC_RND_CONV_false_16_and_1_nl = (~ or_dcpl_967) & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_16_and_9_nl = (~ return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse)
      & return_add_generic_AC_RND_CONV_false_16_and_2_m1c;
  assign return_add_generic_AC_RND_CONV_false_16_or_nl = (return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse
      & return_add_generic_AC_RND_CONV_false_16_and_2_m1c) | return_add_generic_AC_RND_CONV_false_11_and_19_cse
      | return_add_generic_AC_RND_CONV_false_11_and_21_cse;
  assign return_add_generic_AC_RND_CONV_false_7_do_sub_return_add_generic_AC_RND_CONV_false_7_do_sub_xor_nl
      = stage_d_mul_return_d_63_sva_1 ^ stage_d_mul_return_d_2_63_sva_1;
  assign return_add_generic_AC_RND_CONV_false_20_do_sub_return_add_generic_AC_RND_CONV_false_20_do_sub_xor_nl
      = stage_d_mul_return_d_63_sva_1 ^ stage_d_mul_return_d_5_63_sva_1;
  assign return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_or_1_nl
      = (operator_6_false_9_acc_psp_1_sva_1[0]) | (~ return_add_generic_AC_RND_CONV_false_17_acc_3_itm_10);
  assign return_extract_56_and_1_nl = operator_11_true_return_24_sva & return_add_generic_AC_RND_CONV_false_12_mux_itm;
  assign stage_PE_1_tmp_re_d_and_3_nl = (~ inverse_lpi_1_dfm_1) & (fsm_output[10]);
  assign stage_PE_1_tmp_re_d_and_4_nl = inverse_lpi_1_dfm_1 & (fsm_output[10]);
  assign stage_PE_1_tmp_re_d_and_5_nl = (~ inverse_lpi_1_dfm_1) & (fsm_output[35]);
  assign stage_PE_1_tmp_re_d_and_6_nl = inverse_lpi_1_dfm_1 & (fsm_output[35]);
  assign return_add_generic_AC_RND_CONV_false_7_exp_and_6_nl = (~ and_dcpl_469) &
      (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_7_exp_and_7_nl = and_dcpl_469 & (fsm_output[14]);
  assign nor_nl = ~(((z_out_88[53]) & (fsm_output[15])) | ((z_out_88[53]) & (fsm_output[5]))
      | ((z_out_88[53]) & (fsm_output[17])) | ((z_out_88[53]) & (fsm_output[30]))
      | ((z_out_88[53]) & (fsm_output[42])) | ((z_out_88[53]) & (fsm_output[40])));
  assign and_2619_nl = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (z_out_88[51:0]), nor_nl);
  assign or_1760_nl = or_dcpl_485 | (fsm_output[15]) | or_dcpl_528;
  assign or_1761_nl = or_dcpl_625 | or_dcpl_598 | or_dcpl_597;
  assign return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_4_nl
      = (z_out_112[10]) & return_add_generic_AC_RND_CONV_false_17_acc_3_itm_10;
  assign BUTTERFLY_1_else_1_if_and_4_nl = or_1864_ssc & BUTTERFLY_1_else_1_if_or_rgt;
  assign BUTTERFLY_1_else_1_if_and_5_nl = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
      & BUTTERFLY_1_else_1_if_or_rgt;
  assign BUTTERFLY_1_else_1_if_and_6_nl = return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse
      & BUTTERFLY_1_else_1_if_or_rgt;
  assign BUTTERFLY_1_else_1_if_and_7_nl = (fsm_output[12]) & BUTTERFLY_1_else_1_if_or_rgt;
  assign BUTTERFLY_1_else_1_if_and_8_nl = return_extract_22_or_2_cse & BUTTERFLY_1_else_1_if_or_rgt;
  assign BUTTERFLY_1_else_1_if_and_9_nl = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_32_cse
      & BUTTERFLY_1_else_1_if_or_rgt;
  assign BUTTERFLY_1_else_1_if_and_10_nl = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse
      & BUTTERFLY_1_else_1_if_or_rgt;
  assign BUTTERFLY_1_else_1_if_and_11_nl = (fsm_output[38]) & BUTTERFLY_1_else_1_if_or_rgt;
  assign BUTTERFLY_1_else_3_else_mux_2_nl = MUX_v_9_2_2((z_out_58[9:1]), BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_1_9_1,
      inverse_lpi_1_dfm_1);
  assign BUTTERFLY_1_else_3_else_mux_3_nl = MUX_s_1_2_2((z_out_58[0]), BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_1_0,
      inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_22_ma1_lt_ma2_mux_4_nl = MUX_s_1_2_2((~
      return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0), (~ return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0),
      fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_22_ma1_lt_ma2_mux_5_nl = MUX_v_51_2_2((~
      return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1), (~ return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1),
      fsm_output[16]);
  assign nl_acc_nl = ({1'b1 , (stage_PE_1_x_re_d_sva[51:0]) , 1'b1}) + conv_u2u_53_54({return_add_generic_AC_RND_CONV_false_22_ma1_lt_ma2_mux_4_nl
      , return_add_generic_AC_RND_CONV_false_22_ma1_lt_ma2_mux_5_nl , 1'b1});
  assign acc_nl = nl_acc_nl[53:0];
  assign z_out_53_52 = readslicef_54_1_53(acc_nl);
  assign return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_mux1h_4_nl = MUX1HOT_s_1_4_2((~
      return_add_generic_AC_RND_CONV_false_21_m_r_51_lpi_3_dfm_mx0), (~ (out_f_d_rsci_q_d[51])),
      (~ return_add_generic_AC_RND_CONV_false_8_m_r_51_lpi_3_dfm_mx0), (~ (in_f_d_rsci_q_d[51])),
      {(fsm_output[43]) , (fsm_output[5]) , (fsm_output[18]) , (fsm_output[30])});
  assign return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_mux1h_5_nl = MUX1HOT_v_51_4_2((~
      return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1), (~ (out_f_d_rsci_q_d[50:0])),
      (~ return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1), (~ (in_f_d_rsci_q_d[50:0])),
      {(fsm_output[43]) , (fsm_output[5]) , (fsm_output[18]) , (fsm_output[30])});
  assign nl_acc_1_nl = ({1'b1 , (stage_PE_1_tmp_re_d_sva[51:0]) , 1'b1}) + conv_u2u_53_54({return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_mux1h_4_nl
      , return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_mux1h_5_nl , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[53:0];
  assign z_out_54_52 = readslicef_54_1_53(acc_1_nl);
  assign return_add_generic_AC_RND_CONV_false_6_ma1_lt_ma2_mux_5_nl = MUX_s_1_2_2((~
      stage_PE_tmp_re_d_1_lpi_3_dfm_51_mx0), (~ stage_PE_1_tmp_im_d_1_lpi_3_dfm_51_mx1),
      fsm_output[36]);
  assign return_add_generic_AC_RND_CONV_false_6_ma1_lt_ma2_mux_6_nl = MUX_v_51_2_2((~
      return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx1),
      (~ return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm_mx2),
      fsm_output[36]);
  assign nl_acc_4_nl = ({1'b1 , stage_PE_1_tmp_im_d_1_lpi_3_dfm_51 , return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm
      , 1'b1}) + conv_u2u_53_54({return_add_generic_AC_RND_CONV_false_6_ma1_lt_ma2_mux_5_nl
      , return_add_generic_AC_RND_CONV_false_6_ma1_lt_ma2_mux_6_nl , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[53:0];
  assign z_out_57_52 = readslicef_54_1_53(acc_4_nl);
  assign BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_9_nl = MUX_v_16_2_2((signext_16_14(z_out_98[15:2])),
      z_out_60, BUTTERFLY_else_or_cse);
  assign BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_10_nl = MUX_v_2_2_2((z_out_98[1:0]),
      2'b01, BUTTERFLY_else_or_cse);
  assign BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_or_1_nl = (~ or_1341_cse)
      | (fsm_output[6]) | (fsm_output[31]);
  assign BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_and_2_nl
      = MUX_v_2_2_2(2'b00, (z_out_61_15_0[15:14]), BUTTERFLY_else_or_cse);
  assign BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_11_nl = MUX_v_2_2_2((signext_2_1(z_out_98[17])),
      (z_out_61_15_0[13:12]), BUTTERFLY_else_or_cse);
  assign BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_and_3_nl
      = MUX_v_11_2_2(11'b00000000000, (z_out_61_15_0[11:1]), BUTTERFLY_else_or_cse);
  assign BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_12_nl = MUX_s_1_2_2((z_out_98[17]),
      (z_out_61_15_0[0]), BUTTERFLY_else_or_cse);
  assign nl_z_out_58 = ({BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_9_nl
      , BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_10_nl}) + conv_s2u_17_18({BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_or_1_nl
      , BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_and_2_nl
      , BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_11_nl , BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_and_3_nl
      , BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_12_nl});
  assign z_out_58 = nl_z_out_58[17:0];
  assign BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_13_nl = MUX_v_16_2_2((operator_32_false_3_acc_psp_sva_1[15:0]),
      (z_out_98[15:0]), BUTTERFLY_else_or_cse);
  assign nl_z_out_59 = BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_13_nl
      + conv_u2u_14_16(signext_14_13({BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_4_cse
      , 11'b00000000000 , BUTTERFLY_1_else_3_else_BUTTERFLY_1_else_3_else_mux_4_cse}));
  assign z_out_59 = nl_z_out_59[15:0];
  assign nl_z_out_60 = (~ (z_out_105[15:0])) + ({(~ (z_out_105[3:0])) , 12'b000000000001})
      + ({(z_out_105[1:0]) , 14'b01000000000000});
  assign z_out_60 = nl_z_out_60[15:0];
  assign nl_z_out_61_15_0 = conv_u2u_4_16(z_out_60[15:12]) + (~ z_out_60);
  assign z_out_61_15_0 = nl_z_out_61_15_0[15:0];
  assign BUTTERFLY_else_1_if_mux_6_nl = MUX_v_16_2_2(out_u_rsci_q_d, in_u_rsci_q_d,
      fsm_output[31]);
  assign nl_acc_9_nl = ({1'b1 , BUTTERFLY_else_1_if_mux_6_nl , 1'b1}) + conv_u2u_17_18({(~
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0) , (~ BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0)
      , (~ BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1) , 1'b1});
  assign acc_9_nl = nl_acc_9_nl[17:0];
  assign z_out_62 = readslicef_18_17_1(acc_9_nl);
  assign nl_operator_32_false_acc_7_nl = z_out_105 + conv_u2u_30_32({z_out_58 , (z_out_60[11:0])});
  assign operator_32_false_acc_7_nl = nl_operator_32_false_acc_7_nl[31:0];
  assign nl_z_out_64 = conv_u2u_16_17(readslicef_32_16_16(operator_32_false_acc_7_nl))
      + 17'b11100111111111111;
  assign z_out_64 = nl_z_out_64[16:0];
  assign stage_PE_stage_PE_stage_PE_mux_3_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_10,
      t_in_10_0_lpi_1_dfm_1_9, return_extract_26_m_zero_sva);
  assign BUTTERFLY_else_mux_10_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_8,
      stage_PE_stage_PE_stage_PE_mux_3_nl, and_3379_cse);
  assign BUTTERFLY_else_mux_11_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_7,
      stage_PE_1_qr_1_10_1_lpi_2_dfm_8, and_3379_cse);
  assign BUTTERFLY_else_mux_12_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_6,
      stage_PE_1_qr_1_10_1_lpi_2_dfm_7, and_3379_cse);
  assign BUTTERFLY_else_mux_13_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_5,
      stage_PE_1_qr_1_10_1_lpi_2_dfm_6, and_3379_cse);
  assign BUTTERFLY_else_mux_14_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_4,
      stage_PE_1_qr_1_10_1_lpi_2_dfm_5, and_3379_cse);
  assign BUTTERFLY_else_mux_15_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_3,
      stage_PE_1_qr_1_10_1_lpi_2_dfm_4, and_3379_cse);
  assign BUTTERFLY_else_mux_16_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_2,
      stage_PE_1_qr_1_10_1_lpi_2_dfm_3, and_3379_cse);
  assign BUTTERFLY_else_mux_17_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_1,
      stage_PE_1_qr_1_10_1_lpi_2_dfm_2, and_3379_cse);
  assign BUTTERFLY_else_mux_18_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_0,
      stage_PE_1_qr_1_10_1_lpi_2_dfm_1, and_3379_cse);
  assign BUTTERFLY_else_mux_19_nl = MUX_s_1_2_2(stage_PE_1_qr_1_0_lpi_2_dfm, stage_PE_1_qr_1_10_1_lpi_2_dfm_0,
      and_3379_cse);
  assign nl_z_out_66 = ({BUTTERFLY_else_mux_10_nl , BUTTERFLY_else_mux_11_nl , BUTTERFLY_else_mux_12_nl
      , BUTTERFLY_else_mux_13_nl , BUTTERFLY_else_mux_14_nl , BUTTERFLY_else_mux_15_nl
      , BUTTERFLY_else_mux_16_nl , BUTTERFLY_else_mux_17_nl , BUTTERFLY_else_mux_18_nl
      , BUTTERFLY_else_mux_19_nl}) + conv_u2u_9_10(BUTTERFLY_i_div_psp_sva_1);
  assign z_out_66 = nl_z_out_66[9:0];
  assign BUTTERFLY_fry_mux_10_nl = MUX_s_1_2_2(stage_PE_1_qr_0_lpi_2_dfm, stage_PE_1_qr_10_1_lpi_2_dfm_8,
      and_3379_cse);
  assign BUTTERFLY_fry_mux_11_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_8, stage_PE_1_qr_10_1_lpi_2_dfm_7,
      and_3379_cse);
  assign BUTTERFLY_fry_mux_12_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_7, stage_PE_1_qr_10_1_lpi_2_dfm_6,
      and_3379_cse);
  assign BUTTERFLY_fry_mux_13_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_6, stage_PE_1_qr_10_1_lpi_2_dfm_5,
      and_3379_cse);
  assign BUTTERFLY_fry_mux_14_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_5, stage_PE_1_qr_10_1_lpi_2_dfm_4,
      and_3379_cse);
  assign BUTTERFLY_fry_mux_15_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_4, stage_PE_1_qr_10_1_lpi_2_dfm_3,
      and_3379_cse);
  assign BUTTERFLY_fry_mux_16_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_3, stage_PE_1_qr_10_1_lpi_2_dfm_2,
      and_3379_cse);
  assign BUTTERFLY_fry_mux_17_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_2, stage_PE_1_qr_10_1_lpi_2_dfm_1,
      and_3379_cse);
  assign BUTTERFLY_fry_mux_18_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_1, stage_PE_1_qr_10_1_lpi_2_dfm_0,
      and_3379_cse);
  assign BUTTERFLY_fry_mux_19_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_0, stage_PE_1_qr_0_lpi_2_dfm,
      and_3379_cse);
  assign nl_z_out_67 = BUTTERFLY_i_9_0_sva_1 + ({BUTTERFLY_fry_mux_10_nl , BUTTERFLY_fry_mux_11_nl
      , BUTTERFLY_fry_mux_12_nl , BUTTERFLY_fry_mux_13_nl , BUTTERFLY_fry_mux_14_nl
      , BUTTERFLY_fry_mux_15_nl , BUTTERFLY_fry_mux_16_nl , BUTTERFLY_fry_mux_17_nl
      , BUTTERFLY_fry_mux_18_nl , BUTTERFLY_fry_mux_19_nl});
  assign z_out_67 = nl_z_out_67[9:0];
  assign return_mult_generic_AC_RND_CONV_false_2_exp_mux_7_nl = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1, fsm_output[38]);
  assign return_mult_generic_AC_RND_CONV_false_2_exp_mux_8_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1, fsm_output[38]);
  assign nl_acc_10_nl = conv_u2u_12_13({return_mult_generic_AC_RND_CONV_false_2_exp_mux_7_nl
      , return_mult_generic_AC_RND_CONV_false_2_exp_mux_8_nl , 1'b1}) + conv_u2u_2_13({(~
      return_extract_41_return_extract_41_or_1_cse_sva) , 1'b1});
  assign acc_10_nl = nl_acc_10_nl[12:0];
  assign return_mult_generic_AC_RND_CONV_false_2_exp_mux_9_nl = MUX_s_1_2_2(return_extract_19_return_extract_19_nor_tmp,
      return_extract_51_return_extract_51_nor_tmp, fsm_output[38]);
  assign nl_acc_14_nl = conv_u2u_13_14({(readslicef_13_12_1(acc_10_nl)) , return_mult_generic_AC_RND_CONV_false_2_exp_mux_9_nl})
      + conv_s2u_12_14({1'b1 , (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[61:52]) , 1'b1});
  assign acc_14_nl = nl_acc_14_nl[13:0];
  assign z_out_68 = readslicef_14_13_1(acc_14_nl);
  assign return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_6_nl = MUX1HOT_s_1_5_2((out_f_d_rsci_q_d[62]),
      (stage_PE_1_x_re_d_sva[62]), (in_f_d_rsci_q_d[62]), drf_qr_lval_10_smx_lpi_3_dfm_rsp_0,
      (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[9]), {return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse
      , (fsm_output[16]) , (fsm_output[32]) , (fsm_output[36]) , (fsm_output[43])});
  assign return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_7_nl = MUX1HOT_v_9_5_2((out_f_d_rsci_q_d[61:53]),
      (stage_PE_1_x_re_d_sva[61:53]), (in_f_d_rsci_q_d[61:53]), drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0,
      (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[8:0]), {return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse
      , (fsm_output[16]) , (fsm_output[32]) , (fsm_output[36]) , (fsm_output[43])});
  assign return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_8_nl = MUX1HOT_s_1_5_2((out_f_d_rsci_q_d[52]),
      (stage_PE_1_x_re_d_sva[52]), (in_f_d_rsci_q_d[52]), drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1,
      return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1, {return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse
      , (fsm_output[16]) , (fsm_output[32]) , (fsm_output[36]) , (fsm_output[43])});
  assign return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_9_nl = MUX1HOT_v_10_3_2((~
      (stage_PE_1_tmp_re_d_sva[62:53])), (~ return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1),
      (~ drf_qr_lval_10_smx_lpi_3_dfm_mx7_10_1), {return_add_generic_AC_RND_CONV_false_e_dif1_or_1_cse
      , (fsm_output[16]) , (fsm_output[36])});
  assign return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_10_nl = MUX1HOT_s_1_3_2((~
      (stage_PE_1_tmp_re_d_sva[52])), (~ return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1),
      (~ drf_qr_lval_10_smx_lpi_3_dfm_mx7_0), {return_add_generic_AC_RND_CONV_false_e_dif1_or_1_cse
      , (fsm_output[16]) , (fsm_output[36])});
  assign nl_acc_15_nl = ({1'b1 , return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_6_nl
      , return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_7_nl , return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_8_nl
      , 1'b1}) + conv_u2u_12_13({return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_9_nl
      , return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_10_nl , 1'b1});
  assign acc_15_nl = nl_acc_15_nl[12:0];
  assign z_out_69 = readslicef_13_12_1(acc_15_nl);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_and_4_nl = (~ inverse_lpi_1_dfm_1)
      & (fsm_output[11]);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_or_5_nl = (inverse_lpi_1_dfm_1
      & (fsm_output[11])) | (inverse_lpi_1_dfm_1 & (fsm_output[36]));
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_or_6_nl = return_add_generic_AC_RND_CONV_false_11_or_5_cse
      | ((~ inverse_lpi_1_dfm_1) & (fsm_output[36]));
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_6_nl = MUX1HOT_v_10_5_2((stage_PE_1_tmp_re_d_sva[62:53]),
      (out_f_d_rsci_q_d[62:53]), return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0,
      return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1, (in_f_d_rsci_q_d[62:53]),
      {return_add_generic_AC_RND_CONV_false_1_e_dif1_or_cse , return_add_generic_AC_RND_CONV_false_1_e_dif1_and_4_nl
      , return_add_generic_AC_RND_CONV_false_1_e_dif1_or_5_nl , (fsm_output[16])
      , return_add_generic_AC_RND_CONV_false_1_e_dif1_or_6_nl});
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_7_nl = MUX1HOT_s_1_5_2((stage_PE_1_tmp_re_d_sva[52]),
      drf_qr_lval_10_smx_lpi_3_dfm_mx3_0, return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1,
      (in_f_d_rsci_q_d[52]), drf_qr_lval_10_smx_lpi_3_dfm_mx7_0, {return_add_generic_AC_RND_CONV_false_1_e_dif1_or_cse
      , (fsm_output[11]) , (fsm_output[16]) , return_add_generic_AC_RND_CONV_false_11_or_5_cse
      , (fsm_output[36])});
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_8_nl = MUX1HOT_s_1_5_2((~
      (out_f_d_rsci_q_d[62])), (~ drf_qr_lval_10_smx_lpi_3_dfm_rsp_0), (~ (stage_PE_1_x_re_d_sva[62])),
      (~ (stage_PE_1_tmp_re_d_sva[62])), (~ (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[9])),
      {return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse , or_dcpl_680 , (fsm_output[16])
      , return_add_generic_AC_RND_CONV_false_11_or_5_cse , (fsm_output[43])});
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_9_nl = MUX1HOT_v_9_5_2((~
      (out_f_d_rsci_q_d[61:53])), (~ drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0), (~
      (stage_PE_1_x_re_d_sva[61:53])), (~ (stage_PE_1_tmp_re_d_sva[61:53])), (~ (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[8:0])),
      {return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse , or_dcpl_680 , (fsm_output[16])
      , return_add_generic_AC_RND_CONV_false_11_or_5_cse , (fsm_output[43])});
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_10_nl = MUX1HOT_s_1_5_2((~
      (out_f_d_rsci_q_d[52])), (~ drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1), (~ (stage_PE_1_x_re_d_sva[52])),
      (~ (stage_PE_1_tmp_re_d_sva[52])), (~ return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1),
      {return_add_generic_AC_RND_CONV_false_13_op2_mu_or_cse , or_dcpl_680 , (fsm_output[16])
      , return_add_generic_AC_RND_CONV_false_11_or_5_cse , (fsm_output[43])});
  assign nl_acc_16_nl = ({1'b1 , return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_6_nl
      , return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_7_nl , 1'b1}) + conv_u2u_12_13({return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_8_nl
      , return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_9_nl , return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_10_nl
      , 1'b1});
  assign acc_16_nl = nl_acc_16_nl[12:0];
  assign z_out_70 = readslicef_13_12_1(acc_16_nl);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif_mux_3_nl = MUX_v_11_2_2((~
      (out_f_d_rsci_q_d[62:52])), (~ (in_f_d_rsci_q_d[62:52])), fsm_output[30]);
  assign nl_acc_17_nl = ({1'b1 , (stage_PE_1_tmp_re_d_sva[62:52]) , 1'b1}) + conv_u2u_12_13({return_add_generic_AC_RND_CONV_false_1_e_dif_mux_3_nl
      , 1'b1});
  assign acc_17_nl = nl_acc_17_nl[12:0];
  assign z_out_71_11 = readslicef_13_1_12(acc_17_nl);
  assign nl_acc_18_cse_6_1 = ({1'b1 , (~ (rtn_out_2[5:1]))}) + 6'b000001;
  assign acc_18_cse_6_1 = nl_acc_18_cse_6_1[5:0];
  assign return_add_generic_AC_RND_CONV_false_1_or_17_nl = (return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1
      & (~ return_add_generic_AC_RND_CONV_false_11_or_5_cse)) | return_add_generic_AC_RND_CONV_false_11_and_9_itm;
  assign return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_mux_1_nl
      = MUX_v_56_2_2((z_out_73[56:1]), (~ (z_out_73[56:1])), return_add_generic_AC_RND_CONV_false_1_or_17_nl);
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_15_nl = MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_1_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_1_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_14_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_14_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_13_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_13_res_mant_3_0_sva_1), {return_add_generic_AC_RND_CONV_false_12_and_89_cse
      , return_add_generic_AC_RND_CONV_false_12_and_90_cse , return_add_generic_AC_RND_CONV_false_12_and_91_cse
      , return_add_generic_AC_RND_CONV_false_12_and_92_cse , return_add_generic_AC_RND_CONV_false_12_and_97_cse
      , return_add_generic_AC_RND_CONV_false_12_and_98_cse , return_add_generic_AC_RND_CONV_false_12_and_99_cse
      , return_add_generic_AC_RND_CONV_false_12_and_100_cse});
  assign return_add_generic_AC_RND_CONV_false_1_mux_35_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_do_sub_sva_1,
      return_add_generic_AC_RND_CONV_false_14_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_11_or_5_cse);
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_16_nl = MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_1_op1_mu_52_lpi_3_dfm_1, drf_qr_lval_13_smx_0_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_52_lpi_3_dfm_1, {return_add_generic_AC_RND_CONV_false_1_or_6_cse
      , return_add_generic_AC_RND_CONV_false_1_or_7_cse , or_1864_ssc , return_add_generic_AC_RND_CONV_false_1_or_9_cse});
  assign return_add_generic_AC_RND_CONV_false_1_or_18_nl = return_add_generic_AC_RND_CONV_false_1_and_16_cse
      | and_2172_cse | return_add_generic_AC_RND_CONV_false_1_and_20_cse | and_2173_cse;
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_17_nl = MUX1HOT_v_51_3_2(return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm,
      return_extract_2_mux_4_cse, return_extract_33_mux_3_cse, {return_add_generic_AC_RND_CONV_false_1_or_18_nl
      , return_add_generic_AC_RND_CONV_false_1_or_7_cse , return_add_generic_AC_RND_CONV_false_1_or_9_cse});
  assign return_add_generic_AC_RND_CONV_false_1_mux1h_18_nl = MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_13_op2_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1, {return_add_generic_AC_RND_CONV_false_1_or_6_cse
      , return_add_generic_AC_RND_CONV_false_1_or_7_cse , or_1864_ssc , return_add_generic_AC_RND_CONV_false_1_or_9_cse});
  assign nl_acc_19_nl = ({return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_mux_1_nl
      , return_add_generic_AC_RND_CONV_false_1_mux1h_15_nl , return_add_generic_AC_RND_CONV_false_1_mux_35_nl})
      + conv_u2u_57_58({return_add_generic_AC_RND_CONV_false_1_mux1h_16_nl , return_add_generic_AC_RND_CONV_false_1_mux1h_17_nl
      , return_add_generic_AC_RND_CONV_false_1_mux1h_18_nl , 4'b0001});
  assign acc_19_nl = nl_acc_19_nl[57:0];
  assign z_out_80 = readslicef_58_57_1(acc_19_nl);
  assign return_add_generic_AC_RND_CONV_false_12_mux1h_26_nl = MUX1HOT_v_4_8_2(return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_0,
      (return_add_generic_AC_RND_CONV_false_11_mux_1_itm[55:52]), (return_add_generic_AC_RND_CONV_false_18_mux_1_itm_55_50[5:2]),
      (return_add_generic_AC_RND_CONV_false_9_mux_28_cse[55:52]), (return_add_generic_AC_RND_CONV_false_6_res_mant_conc_2_itm_56_1[55:52]),
      (return_add_generic_AC_RND_CONV_false_7_mux_31_cse[55:52]), (return_add_generic_AC_RND_CONV_false_10_mux_28_cse[55:52]),
      (return_add_generic_AC_RND_CONV_false_19_res_mant_conc_2_itm_56_1[55:52]),
      {return_add_generic_AC_RND_CONV_false_12_or_41_cse , return_add_generic_AC_RND_CONV_false_12_or_9_cse
      , operator_6_false_17_or_cse , return_add_generic_AC_RND_CONV_false_12_or_11_cse_1
      , (fsm_output[11]) , return_add_generic_AC_RND_CONV_false_10_ls_or_2_cse ,
      return_add_generic_AC_RND_CONV_false_10_r_zero_or_2_cse , (fsm_output[36])});
  assign return_add_generic_AC_RND_CONV_false_12_mux1h_27_nl = MUX1HOT_v_2_8_2((return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1[51:50]),
      (return_add_generic_AC_RND_CONV_false_11_mux_1_itm[51:50]), (return_add_generic_AC_RND_CONV_false_18_mux_1_itm_55_50[1:0]),
      (return_add_generic_AC_RND_CONV_false_9_mux_28_cse[51:50]), (return_add_generic_AC_RND_CONV_false_6_res_mant_conc_2_itm_56_1[51:50]),
      (return_add_generic_AC_RND_CONV_false_7_mux_31_cse[51:50]), (return_add_generic_AC_RND_CONV_false_10_mux_28_cse[51:50]),
      (return_add_generic_AC_RND_CONV_false_19_res_mant_conc_2_itm_56_1[51:50]),
      {return_add_generic_AC_RND_CONV_false_12_or_41_cse , return_add_generic_AC_RND_CONV_false_12_or_9_cse
      , operator_6_false_17_or_cse , return_add_generic_AC_RND_CONV_false_12_or_11_cse_1
      , (fsm_output[11]) , return_add_generic_AC_RND_CONV_false_10_ls_or_2_cse ,
      return_add_generic_AC_RND_CONV_false_10_r_zero_or_2_cse , (fsm_output[36])});
  assign return_add_generic_AC_RND_CONV_false_12_mux1h_28_nl = MUX1HOT_v_50_8_2((return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_55_0_rsp_1[49:0]),
      (return_add_generic_AC_RND_CONV_false_11_mux_1_itm[49:0]), return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0,
      (return_add_generic_AC_RND_CONV_false_9_mux_28_cse[49:0]), (return_add_generic_AC_RND_CONV_false_6_res_mant_conc_2_itm_56_1[49:0]),
      (return_add_generic_AC_RND_CONV_false_7_mux_31_cse[49:0]), (return_add_generic_AC_RND_CONV_false_10_mux_28_cse[49:0]),
      (return_add_generic_AC_RND_CONV_false_19_res_mant_conc_2_itm_56_1[49:0]), {return_add_generic_AC_RND_CONV_false_12_or_41_cse
      , return_add_generic_AC_RND_CONV_false_12_or_9_cse , operator_6_false_17_or_cse
      , return_add_generic_AC_RND_CONV_false_12_or_11_cse_1 , (fsm_output[11]) ,
      return_add_generic_AC_RND_CONV_false_10_ls_or_2_cse , return_add_generic_AC_RND_CONV_false_10_r_zero_or_2_cse
      , (fsm_output[36])});
  assign return_add_generic_AC_RND_CONV_false_12_or_47_nl = or_dcpl_534 | BUTTERFLY_else_or_cse
      | or_dcpl_553 | or_dcpl_493;
  assign return_add_generic_AC_RND_CONV_false_12_and_121_nl = (~ return_add_generic_AC_RND_CONV_false_18_mux_itm)
      & (fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_12_and_122_nl = return_add_generic_AC_RND_CONV_false_18_mux_itm
      & (fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_12_and_123_nl = (~ return_add_generic_AC_RND_CONV_false_11_do_sub_sva)
      & or_tmp_1400;
  assign return_add_generic_AC_RND_CONV_false_12_and_124_nl = return_add_generic_AC_RND_CONV_false_11_do_sub_sva
      & or_tmp_1400;
  assign return_add_generic_AC_RND_CONV_false_12_and_125_nl = (~ return_add_generic_AC_RND_CONV_false_18_mux_itm)
      & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_12_and_126_nl = return_add_generic_AC_RND_CONV_false_18_mux_itm
      & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_12_and_127_nl = (~ not_tmp_376) & (fsm_output[11]);
  assign return_add_generic_AC_RND_CONV_false_12_and_128_nl = not_tmp_376 & (fsm_output[11]);
  assign return_add_generic_AC_RND_CONV_false_12_and_129_nl = (~ return_add_generic_AC_RND_CONV_false_20_do_sub_sva)
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_12_and_130_nl = return_add_generic_AC_RND_CONV_false_20_do_sub_sva
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_12_and_131_nl = (~ return_add_generic_AC_RND_CONV_false_10_do_sub_sva)
      & (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_12_and_132_nl = return_add_generic_AC_RND_CONV_false_10_do_sub_sva
      & (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_12_and_133_nl = (~ not_tmp_395) & (fsm_output[36]);
  assign return_add_generic_AC_RND_CONV_false_12_and_134_nl = not_tmp_395 & (fsm_output[36]);
  assign return_add_generic_AC_RND_CONV_false_12_and_135_nl = (~ return_add_generic_AC_RND_CONV_false_20_do_sub_sva)
      & (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_12_and_136_nl = return_add_generic_AC_RND_CONV_false_20_do_sub_sva
      & (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_12_and_137_nl = (~ return_add_generic_AC_RND_CONV_false_10_do_sub_sva)
      & (fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_12_and_138_nl = return_add_generic_AC_RND_CONV_false_10_do_sub_sva
      & (fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_12_mux1h_29_nl = MUX1HOT_s_1_21_2(return_add_generic_AC_RND_CONV_false_12_mux_2_itm,
      drf_qr_lval_15_smx_0_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_9_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_9_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_11_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_11_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_23_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_23_res_mant_3_0_sva_1), BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm,
      (~ return_add_generic_AC_RND_CONV_false_6_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_6_res_mant_3_0_sva_1,
      return_add_generic_AC_RND_CONV_false_7_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_7_res_mant_3_0_sva_1),
      return_add_generic_AC_RND_CONV_false_10_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_10_res_mant_3_0_sva_1),
      (~ return_add_generic_AC_RND_CONV_false_19_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_19_res_mant_3_0_sva_1,
      return_add_generic_AC_RND_CONV_false_20_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_20_res_mant_3_0_sva_1),
      return_add_generic_AC_RND_CONV_false_22_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_22_res_mant_3_0_sva_1),
      {return_add_generic_AC_RND_CONV_false_12_or_47_nl , operator_6_false_17_or_cse
      , return_add_generic_AC_RND_CONV_false_12_and_121_nl , return_add_generic_AC_RND_CONV_false_12_and_122_nl
      , return_add_generic_AC_RND_CONV_false_12_and_123_nl , return_add_generic_AC_RND_CONV_false_12_and_124_nl
      , return_add_generic_AC_RND_CONV_false_12_and_125_nl , return_add_generic_AC_RND_CONV_false_12_and_126_nl
      , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse , return_add_generic_AC_RND_CONV_false_12_and_127_nl
      , return_add_generic_AC_RND_CONV_false_12_and_128_nl , return_add_generic_AC_RND_CONV_false_12_and_129_nl
      , return_add_generic_AC_RND_CONV_false_12_and_130_nl , return_add_generic_AC_RND_CONV_false_12_and_131_nl
      , return_add_generic_AC_RND_CONV_false_12_and_132_nl , return_add_generic_AC_RND_CONV_false_12_and_133_nl
      , return_add_generic_AC_RND_CONV_false_12_and_134_nl , return_add_generic_AC_RND_CONV_false_12_and_135_nl
      , return_add_generic_AC_RND_CONV_false_12_and_136_nl , return_add_generic_AC_RND_CONV_false_12_and_137_nl
      , return_add_generic_AC_RND_CONV_false_12_and_138_nl});
  assign return_add_generic_AC_RND_CONV_false_12_or_48_nl = or_dcpl_534 | or_dcpl_553;
  assign return_add_generic_AC_RND_CONV_false_12_or_49_nl = BUTTERFLY_else_or_cse
      | or_dcpl_493;
  assign return_add_generic_AC_RND_CONV_false_12_or_50_nl = operator_6_false_17_or_cse
      | or_tmp_1400;
  assign return_add_generic_AC_RND_CONV_false_12_or_51_nl = return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse
      | (fsm_output[18]) | (fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_12_mux1h_30_nl = MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_12_do_sub_sva,
      return_add_generic_AC_RND_CONV_false_16_do_sub_sva, return_add_generic_AC_RND_CONV_false_11_do_sub_sva,
      return_add_generic_AC_RND_CONV_false_18_mux_itm, return_add_generic_AC_RND_CONV_false_10_do_sub_sva,
      return_add_generic_AC_RND_CONV_false_6_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_20_do_sub_sva,
      return_add_generic_AC_RND_CONV_false_19_do_sub_sva_1, {return_add_generic_AC_RND_CONV_false_12_or_48_nl
      , return_add_generic_AC_RND_CONV_false_12_or_49_nl , return_add_generic_AC_RND_CONV_false_12_or_50_nl
      , return_add_generic_AC_RND_CONV_false_12_or_11_cse_1 , return_add_generic_AC_RND_CONV_false_12_or_51_nl
      , (fsm_output[11]) , return_add_generic_AC_RND_CONV_false_10_ls_or_2_cse ,
      (fsm_output[36])});
  assign return_add_generic_AC_RND_CONV_false_12_or_52_nl = BUTTERFLY_else_or_cse
      | or_dcpl_553 | or_dcpl_493;
  assign return_add_generic_AC_RND_CONV_false_12_or_53_nl = return_add_generic_AC_RND_CONV_false_12_and_29_cse
      | return_add_generic_AC_RND_CONV_false_12_and_31_cse | return_add_generic_AC_RND_CONV_false_12_and_39_cse;
  assign return_add_generic_AC_RND_CONV_false_12_or_54_nl = return_add_generic_AC_RND_CONV_false_12_and_33_cse
      | return_add_generic_AC_RND_CONV_false_12_and_35_cse | return_add_generic_AC_RND_CONV_false_12_and_37_cse;
  assign return_add_generic_AC_RND_CONV_false_12_mux1h_31_nl = MUX1HOT_s_1_15_2(return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_itm,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm, return_add_generic_AC_RND_CONV_false_23_op1_mu_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm,
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm_mx1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1, drf_qr_lval_13_smx_0_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx0, drf_qr_lval_13_smx_0_lpi_3_dfm_mx3,
      return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0,
      {return_add_generic_AC_RND_CONV_false_12_or_22_cse , return_add_generic_AC_RND_CONV_false_12_or_52_nl
      , return_add_generic_AC_RND_CONV_false_12_or_24_cse , and_1251_cse , or_tmp_1400
      , or_1993_cse , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse ,
      return_add_generic_AC_RND_CONV_false_12_or_53_nl , return_add_generic_AC_RND_CONV_false_12_and_30_cse
      , return_add_generic_AC_RND_CONV_false_12_and_32_cse , return_add_generic_AC_RND_CONV_false_12_or_54_nl
      , or_tmp_946 , return_add_generic_AC_RND_CONV_false_12_and_36_cse , return_add_generic_AC_RND_CONV_false_12_and_38_cse
      , and_1057_cse});
  assign return_add_generic_AC_RND_CONV_false_12_mux1h_32_nl = MUX1HOT_s_1_16_2(return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm,
      (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[50]), return_add_generic_AC_RND_CONV_false_18_op_bigger_mux_1_itm_50,
      (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[50]), return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm, return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_50, return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm_mx1,
      return_add_generic_AC_RND_CONV_false_7_mux_27_cse, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm,
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm_mx3,
      return_add_generic_AC_RND_CONV_false_20_mux_27_cse, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0,
      {or_dcpl_534 , return_add_generic_AC_RND_CONV_false_12_or_27_cse , operator_6_false_17_or_cse
      , return_add_generic_AC_RND_CONV_false_12_or_24_cse , and_1251_cse , or_tmp_1400
      , or_1993_cse , return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse ,
      return_add_generic_AC_RND_CONV_false_12_or_29_cse , return_add_generic_AC_RND_CONV_false_12_and_30_cse
      , return_add_generic_AC_RND_CONV_false_12_and_32_cse , or_dcpl_493 , or_tmp_946
      , return_add_generic_AC_RND_CONV_false_12_and_36_cse , return_add_generic_AC_RND_CONV_false_12_and_38_cse
      , and_1057_cse});
  assign return_add_generic_AC_RND_CONV_false_12_or_55_nl = or_tmp_1400 | return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse
      | or_dcpl_493;
  assign return_add_generic_AC_RND_CONV_false_12_mux1h_33_nl = MUX1HOT_v_50_12_2(return_add_generic_AC_RND_CONV_false_18_op_bigger_mux_1_itm_49_0,
      (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49:0]), (return_add_generic_AC_RND_CONV_false_23_op1_mu_51_1_lpi_3_dfm[49:0]),
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_1_itm_49_0,
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_18_mux_1_itm_49_0,
      return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_49_0_mx0, return_extract_21_mux_cse,
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0_mx0,
      return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0, {return_add_generic_AC_RND_CONV_false_12_or_22_cse
      , return_add_generic_AC_RND_CONV_false_12_or_27_cse , return_add_generic_AC_RND_CONV_false_12_or_24_cse
      , and_1251_cse , return_add_generic_AC_RND_CONV_false_12_or_55_nl , or_1993_cse
      , return_add_generic_AC_RND_CONV_false_12_or_29_cse , return_add_generic_AC_RND_CONV_false_12_and_30_cse
      , return_add_generic_AC_RND_CONV_false_12_or_44_cse , or_tmp_946 , return_add_generic_AC_RND_CONV_false_12_and_36_cse
      , and_1057_cse});
  assign return_add_generic_AC_RND_CONV_false_12_or_56_nl = BUTTERFLY_else_or_cse
      | or_tmp_1400 | or_dcpl_553;
  assign return_add_generic_AC_RND_CONV_false_12_or_57_nl = return_add_generic_AC_RND_CONV_false_12_and_25_cse
      | return_add_generic_AC_RND_CONV_false_12_and_39_cse;
  assign return_add_generic_AC_RND_CONV_false_12_or_58_nl = return_add_generic_AC_RND_CONV_false_12_and_27_cse
      | return_add_generic_AC_RND_CONV_false_12_and_33_cse;
  assign return_add_generic_AC_RND_CONV_false_12_or_59_nl = return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse
      | or_dcpl_493;
  assign return_add_generic_AC_RND_CONV_false_12_or_60_nl = return_add_generic_AC_RND_CONV_false_12_and_29_cse
      | return_add_generic_AC_RND_CONV_false_12_and_35_cse;
  assign return_add_generic_AC_RND_CONV_false_12_mux1h_34_nl = MUX1HOT_s_1_15_2(return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm, return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm,
      return_add_generic_AC_RND_CONV_false_6_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_19_op2_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1,
      {return_add_generic_AC_RND_CONV_false_12_or_22_cse , return_add_generic_AC_RND_CONV_false_12_or_56_nl
      , return_add_generic_AC_RND_CONV_false_12_or_57_nl , and_1251_cse , return_add_generic_AC_RND_CONV_false_12_or_58_nl
      , or_1993_cse , return_add_generic_AC_RND_CONV_false_12_or_59_nl , return_add_generic_AC_RND_CONV_false_12_or_60_nl
      , return_add_generic_AC_RND_CONV_false_12_and_30_cse , return_add_generic_AC_RND_CONV_false_12_and_31_cse
      , return_add_generic_AC_RND_CONV_false_12_or_44_cse , or_tmp_946 , return_add_generic_AC_RND_CONV_false_12_and_36_cse
      , return_add_generic_AC_RND_CONV_false_12_and_37_cse , and_1057_cse});
  assign nl_acc_20_nl = ({return_add_generic_AC_RND_CONV_false_12_mux1h_26_nl , return_add_generic_AC_RND_CONV_false_12_mux1h_27_nl
      , return_add_generic_AC_RND_CONV_false_12_mux1h_28_nl , return_add_generic_AC_RND_CONV_false_12_mux1h_29_nl
      , return_add_generic_AC_RND_CONV_false_12_mux1h_30_nl}) + conv_u2u_57_58({return_add_generic_AC_RND_CONV_false_12_mux1h_31_nl
      , return_add_generic_AC_RND_CONV_false_12_mux1h_32_nl , return_add_generic_AC_RND_CONV_false_12_mux1h_33_nl
      , return_add_generic_AC_RND_CONV_false_12_mux1h_34_nl , 4'b0001});
  assign acc_20_nl = nl_acc_20_nl[57:0];
  assign z_out_81 = readslicef_58_57_1(acc_20_nl);
  assign nl_z_out_82 = conv_s2u_17_18(z_out_62) + conv_u2u_14_18(signext_14_13({(z_out_62[16])
      , 11'b00000000000 , (z_out_62[16])}));
  assign z_out_82 = nl_z_out_82[17:0];
  assign operator_6_false_2_mux1h_3_nl = MUX1HOT_v_11_4_2(drf_qr_lval_1_smx_lpi_3_dfm_mx0,
      drf_qr_lval_10_smx_lpi_3_dfm_mx2, return_extract_32_mux_cse, drf_qr_lval_10_smx_lpi_3_dfm_mx6,
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[30]) , (fsm_output[32])});
  assign nl_operator_6_false_2_acc_1_nl = ({1'b1 , (~ (rtn_out_1[5:1]))}) + 6'b000001;
  assign operator_6_false_2_acc_1_nl = nl_operator_6_false_2_acc_1_nl[5:0];
  assign nl_operator_6_false_acc_1_nl = ({1'b1 , (~ (rtn_out_1[5:1]))}) + 6'b000001;
  assign operator_6_false_acc_1_nl = nl_operator_6_false_acc_1_nl[5:0];
  assign nl_operator_6_false_31_acc_1_nl = ({1'b1 , (~ (rtn_out_1[5:1]))}) + 6'b000001;
  assign operator_6_false_31_acc_1_nl = nl_operator_6_false_31_acc_1_nl[5:0];
  assign nl_operator_6_false_29_acc_1_nl = ({1'b1 , (~ (rtn_out_1[5:1]))}) + 6'b000001;
  assign operator_6_false_29_acc_1_nl = nl_operator_6_false_29_acc_1_nl[5:0];
  assign operator_6_false_2_mux1h_4_nl = MUX1HOT_v_6_4_2(operator_6_false_2_acc_1_nl,
      operator_6_false_acc_1_nl, operator_6_false_31_acc_1_nl, operator_6_false_29_acc_1_nl,
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[30]) , (fsm_output[32])});
  assign nl_z_out_84 = conv_u2u_11_13(operator_6_false_2_mux1h_3_nl) + conv_s2u_7_13({operator_6_false_2_mux1h_4_nl
      , (~ (rtn_out_1[0]))});
  assign z_out_84 = nl_z_out_84[12:0];
  assign operator_6_false_33_mux1h_6_nl = MUX1HOT_s_1_6_2(drf_qr_lval_10_smx_lpi_3_dfm_rsp_0,
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0, (operator_14_false_1_acc_psp_sva_9_0[9]),
      (drf_qr_lval_21_smx_9_0_lpi_3_dfm[9]), (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[9]),
      (drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0[8]), {or_tmp_1439 , or_tmp_1440 ,
      operator_6_false_33_or_5_cse , operator_6_false_33_or_7_cse , operator_6_false_33_or_1_cse
      , operator_6_false_33_or_3_cse});
  assign operator_6_false_33_mux1h_7_nl = MUX1HOT_v_8_6_2((drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0[8:1]),
      (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1[9:2]), (operator_14_false_1_acc_psp_sva_9_0[8:1]),
      (drf_qr_lval_21_smx_9_0_lpi_3_dfm[8:1]), (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[8:1]),
      (drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0[7:0]), {or_tmp_1439 , or_tmp_1440
      , operator_6_false_33_or_5_cse , operator_6_false_33_or_7_cse , operator_6_false_33_or_1_cse
      , operator_6_false_33_or_3_cse});
  assign operator_6_false_33_mux1h_8_nl = MUX1HOT_s_1_6_2((drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0[0]),
      (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1[1]), (operator_14_false_1_acc_psp_sva_9_0[0]),
      (drf_qr_lval_21_smx_9_0_lpi_3_dfm[0]), (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[0]),
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1, {or_tmp_1439 , or_tmp_1440 , operator_6_false_33_or_5_cse
      , operator_6_false_33_or_7_cse , operator_6_false_33_or_1_cse , operator_6_false_33_or_3_cse});
  assign operator_6_false_33_or_22_nl = (fsm_output[23]) | (fsm_output[48]);
  assign operator_6_false_33_mux1h_9_nl = MUX1HOT_s_1_6_2(drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1,
      (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1[0]), BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm,
      drf_qr_lval_13_smx_0_lpi_3_dfm, drf_qr_lval_14_smx_0_lpi_3_dfm, drf_qr_lval_15_smx_0_lpi_3_dfm,
      {or_tmp_1439 , or_tmp_1440 , or_dcpl_534 , or_tmp_450 , operator_6_false_33_or_22_nl
      , BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx0c8});
  assign nl_operator_6_false_23_acc_3_nl = ({1'b1 , (~ (return_add_generic_AC_RND_CONV_false_10_ls_sva[5:1]))})
      + 6'b000001;
  assign operator_6_false_23_acc_3_nl = nl_operator_6_false_23_acc_3_nl[5:0];
  assign nl_operator_6_false_27_acc_3_nl = ({1'b1 , (~ (operator_6_false_17_acc_itm_6_1[5:1]))})
      + 6'b000001;
  assign operator_6_false_27_acc_3_nl = nl_operator_6_false_27_acc_3_nl[5:0];
  assign operator_6_false_33_mux1h_10_nl = MUX1HOT_v_6_5_2(operator_6_false_17_acc_itm_6_1,
      operator_6_false_21_acc_itm_6_1, operator_6_false_23_acc_3_nl, (z_out_101[5:0]),
      operator_6_false_27_acc_3_nl, {operator_6_false_33_or_12_cse , or_dcpl_534
      , operator_6_false_33_or_14_cse , operator_6_false_33_or_15_cse , BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx0c8});
  assign operator_6_false_33_mux1h_11_nl = MUX1HOT_s_1_5_2(operator_6_false_17_acc_itm_0,
      operator_6_false_21_acc_itm_0, (~ (return_add_generic_AC_RND_CONV_false_10_ls_sva[0])),
      (~ (return_add_generic_AC_RND_CONV_false_11_ls_sva[0])), (~ (operator_6_false_17_acc_itm_6_1[0])),
      {operator_6_false_33_or_12_cse , or_dcpl_534 , operator_6_false_33_or_14_cse
      , operator_6_false_33_or_15_cse , BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx0c8});
  assign nl_z_out_85 = conv_u2u_11_13({operator_6_false_33_mux1h_6_nl , operator_6_false_33_mux1h_7_nl
      , operator_6_false_33_mux1h_8_nl , operator_6_false_33_mux1h_9_nl}) + conv_s2u_7_13({operator_6_false_33_mux1h_10_nl
      , operator_6_false_33_mux1h_11_nl});
  assign z_out_85 = nl_z_out_85[12:0];
  assign return_mult_generic_AC_RND_CONV_false_exp_mux1h_6_nl = MUX1HOT_v_10_4_2(return_add_generic_AC_RND_CONV_false_4_e_r_qr_10_1_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_5_e_r_qr_10_1_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_17_e_r_qr_10_1_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_18_e_r_qr_10_1_lpi_3_dfm_1, {(fsm_output[11])
      , (fsm_output[12]) , (fsm_output[36]) , (fsm_output[37])});
  assign return_mult_generic_AC_RND_CONV_false_exp_mux1h_7_nl = MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_18_e_r_qr_0_lpi_3_dfm_1, {(fsm_output[11])
      , (fsm_output[12]) , (fsm_output[36]) , (fsm_output[37])});
  assign nl_acc_22_nl = conv_u2u_12_13({return_mult_generic_AC_RND_CONV_false_exp_mux1h_6_nl
      , return_mult_generic_AC_RND_CONV_false_exp_mux1h_7_nl , 1'b1}) + conv_s2u_12_13({10'b1000000000
      , (~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm) , 1'b1});
  assign acc_22_nl = nl_acc_22_nl[12:0];
  assign return_mult_generic_AC_RND_CONV_false_exp_mux1h_8_nl = MUX1HOT_s_1_4_2(return_extract_15_return_extract_15_nor_tmp,
      return_extract_17_return_extract_17_nor_tmp, return_extract_47_return_extract_47_nor_tmp,
      return_extract_49_return_extract_49_nor_tmp, {(fsm_output[11]) , (fsm_output[12])
      , (fsm_output[36]) , (fsm_output[37])});
  assign nl_acc_25_nl = conv_s2u_13_14({(readslicef_13_12_1(acc_22_nl)) , return_mult_generic_AC_RND_CONV_false_exp_mux1h_8_nl})
      + conv_u2u_12_14({drf_qr_lval_10_smx_lpi_3_dfm_rsp_0 , drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0
      , drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1 , 1'b1});
  assign acc_25_nl = nl_acc_25_nl[13:0];
  assign z_out_86 = readslicef_14_13_1(acc_25_nl);
  assign mux1h_29_nl = MUX1HOT_s_1_3_2((z_out_106[104]), (z_out_106[103]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_1,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_23_nl = MUX1HOT_s_1_3_2((z_out_106[103]), (z_out_106[102]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_2,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_34_nl = MUX1HOT_s_1_3_2((z_out_106[102]), (z_out_106[101]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_3,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_27_nl = MUX1HOT_s_1_3_2((z_out_106[101]), (z_out_106[100]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_4,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_31_nl = MUX1HOT_s_1_3_2((z_out_106[100]), (z_out_106[99]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_5,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_24_nl = MUX1HOT_s_1_3_2((z_out_106[99]), (z_out_106[98]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_6,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_22_nl = MUX1HOT_s_1_3_2((z_out_106[98]), (z_out_106[97]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_7,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_33_nl = MUX1HOT_s_1_3_2((z_out_106[97]), (z_out_106[96]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_8,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_26_nl = MUX1HOT_s_1_3_2((z_out_106[96]), (z_out_106[95]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_9,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_36_nl = MUX1HOT_s_1_3_2((z_out_106[95]), (z_out_106[94]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_10,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_35_nl = MUX1HOT_s_1_3_2((z_out_106[94]), (z_out_106[93]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_11,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_56_nl = MUX1HOT_s_1_3_2((z_out_106[93]), (z_out_106[92]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_12,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_57_nl = MUX1HOT_s_1_3_2((z_out_106[92]), (z_out_106[91]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_13,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_38_nl = MUX1HOT_s_1_3_2((z_out_106[91]), (z_out_106[90]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_14,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_58_nl = MUX1HOT_s_1_3_2((z_out_106[90]), (z_out_106[89]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_15,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_55_nl = MUX1HOT_s_1_3_2((z_out_106[89]), (z_out_106[88]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_16,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_45_nl = MUX1HOT_s_1_3_2((z_out_106[88]), (z_out_106[87]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_17,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_54_nl = MUX1HOT_s_1_3_2((z_out_106[87]), (z_out_106[86]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_18,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_60_nl = MUX1HOT_s_1_3_2((z_out_106[86]), (z_out_106[85]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_19,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_59_nl = MUX1HOT_s_1_3_2((z_out_106[85]), (z_out_106[84]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_20,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_32_nl = MUX1HOT_s_1_3_2((z_out_106[84]), (z_out_106[83]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_21,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_28_nl = MUX1HOT_s_1_3_2((z_out_106[83]), (z_out_106[82]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_22,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_51_nl = MUX1HOT_s_1_3_2((z_out_106[82]), (z_out_106[81]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_23,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_46_nl = MUX1HOT_s_1_3_2((z_out_106[81]), (z_out_106[80]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_24,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_8_nl = MUX1HOT_s_1_3_2((z_out_106[80]), (z_out_106[79]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_25,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_9_nl = MUX1HOT_s_1_3_2((z_out_106[79]), (z_out_106[78]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_26,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_10_nl = MUX1HOT_s_1_3_2((z_out_106[78]), (z_out_106[77]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_27,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_11_nl = MUX1HOT_s_1_3_2((z_out_106[77]), (z_out_106[76]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_28,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_30_nl = MUX1HOT_s_1_3_2((z_out_106[76]), (z_out_106[75]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_29,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_20_nl = MUX1HOT_s_1_3_2((z_out_106[75]), (z_out_106[74]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_30,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_19_nl = MUX1HOT_s_1_3_2((z_out_106[74]), (z_out_106[73]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_31,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_18_nl = MUX1HOT_s_1_3_2((z_out_106[73]), (z_out_106[72]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_32,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_17_nl = MUX1HOT_s_1_3_2((z_out_106[72]), (z_out_106[71]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_33,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_16_nl = MUX1HOT_s_1_3_2((z_out_106[71]), (z_out_106[70]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_34,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_15_nl = MUX1HOT_s_1_3_2((z_out_106[70]), (z_out_106[69]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_35,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_14_nl = MUX1HOT_s_1_3_2((z_out_106[69]), (z_out_106[68]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_36,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_13_nl = MUX1HOT_s_1_3_2((z_out_106[68]), (z_out_106[67]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_37,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_12_nl = MUX1HOT_s_1_3_2((z_out_106[67]), (z_out_106[66]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_38,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_49_nl = MUX1HOT_s_1_3_2((z_out_106[66]), (z_out_106[65]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_39,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_44_nl = MUX1HOT_s_1_3_2((z_out_106[65]), (z_out_106[64]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_40,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_41_nl = MUX1HOT_s_1_3_2((z_out_106[64]), (z_out_106[63]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_41,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_52_nl = MUX1HOT_s_1_3_2((z_out_106[63]), (z_out_106[62]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_42,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_53_nl = MUX1HOT_s_1_3_2((z_out_106[62]), (z_out_106[61]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_43,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_47_nl = MUX1HOT_s_1_3_2((z_out_106[61]), (z_out_106[60]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_44,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_42_nl = MUX1HOT_s_1_3_2((z_out_106[60]), (z_out_106[59]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_45,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_39_nl = MUX1HOT_s_1_3_2((z_out_106[59]), (z_out_106[58]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_46,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_43_nl = MUX1HOT_s_1_3_2((z_out_106[58]), (z_out_106[57]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_47,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_50_nl = MUX1HOT_s_1_3_2((z_out_106[57]), (z_out_106[56]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_48,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_48_nl = MUX1HOT_s_1_3_2((z_out_106[56]), (z_out_106[55]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_49,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_40_nl = MUX1HOT_s_1_3_2((z_out_106[55]), (z_out_106[54]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_50,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_37_nl = MUX1HOT_s_1_3_2((z_out_106[54]), (z_out_106[53]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_51,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign mux1h_25_nl = MUX1HOT_s_1_3_2((z_out_106[52]), (z_out_106[51]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_53,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign return_mult_generic_AC_RND_CONV_false_if_1_or_3_nl = (z_out_106[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_if_1_aelse_return_mult_generic_AC_RND_CONV_false_if_1_aelse_or_2
      & (z_out_106[51]));
  assign return_mult_generic_AC_RND_CONV_false_mux_16_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_if_1_or_3_nl,
      drf_qr_lval_14_smx_0_lpi_3_dfm, operator_14_false_1_acc_psp_sva_12_10[2]);
  assign return_mult_generic_AC_RND_CONV_false_and_3_nl = mux1h_25_nl & (return_mult_generic_AC_RND_CONV_false_mux_16_nl
      | z_out_13);
  assign nl_z_out_87 = ({mux1h_29_nl , mux1h_23_nl , mux1h_34_nl , mux1h_27_nl ,
      mux1h_31_nl , mux1h_24_nl , mux1h_22_nl , mux1h_33_nl , mux1h_26_nl , mux1h_36_nl
      , mux1h_35_nl , mux1h_56_nl , mux1h_57_nl , mux1h_38_nl , mux1h_58_nl , mux1h_55_nl
      , mux1h_45_nl , mux1h_54_nl , mux1h_60_nl , mux1h_59_nl , mux1h_32_nl , mux1h_28_nl
      , mux1h_51_nl , mux1h_46_nl , mux1h_8_nl , mux1h_9_nl , mux1h_10_nl , mux1h_11_nl
      , mux1h_30_nl , mux1h_20_nl , mux1h_19_nl , mux1h_18_nl , mux1h_17_nl , mux1h_16_nl
      , mux1h_15_nl , mux1h_14_nl , mux1h_13_nl , mux1h_12_nl , mux1h_49_nl , mux1h_44_nl
      , mux1h_41_nl , mux1h_52_nl , mux1h_53_nl , mux1h_47_nl , mux1h_42_nl , mux1h_39_nl
      , mux1h_43_nl , mux1h_50_nl , mux1h_48_nl , mux1h_40_nl , mux1h_37_nl , z_out_13})
      + conv_u2u_1_52(return_mult_generic_AC_RND_CONV_false_and_3_nl);
  assign z_out_87 = nl_z_out_87[51:0];
  assign return_add_generic_AC_RND_CONV_false_1_res_rounded_mux_1_nl = MUX_s_1_2_2((z_out_77[56]),
      (z_out_79[56]), return_add_generic_AC_RND_CONV_false_1_res_rounded_or_2_cse);
  assign return_add_generic_AC_RND_CONV_false_1_res_rounded_return_add_generic_AC_RND_CONV_false_1_res_rounded_and_1_nl
      = return_add_generic_AC_RND_CONV_false_1_res_rounded_mux_1_nl & (~ (fsm_output[54]));
  assign return_add_generic_AC_RND_CONV_false_1_res_rounded_mux1h_3_nl = MUX1HOT_v_52_3_2((z_out_77[55:4]),
      (z_out_79[55:4]), (return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1[52:1]),
      {return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse , return_add_generic_AC_RND_CONV_false_1_res_rounded_or_2_cse
      , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_1_res_rounded_and_1_nl = (z_out_77[3])
      & ((z_out_77[0]) | (z_out_77[1]) | (z_out_77[2]) | (z_out_77[4]));
  assign return_mult_generic_AC_RND_CONV_false_6_if_1_or_1_nl = (z_out_106[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_or_2
      & (z_out_106[51]));
  assign return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_or_1_tmp
      & (~ (z_out_107[51]))) | ((out_f_d_rsci_q_d[51]) & (~ (z_out_107[50]))) | ((out_f_d_rsci_q_d[50])
      & (~ (z_out_107[49]))) | ((out_f_d_rsci_q_d[49]) & (~ (z_out_107[48]))) | ((out_f_d_rsci_q_d[48])
      & (~ (z_out_107[47]))) | ((out_f_d_rsci_q_d[47]) & (~ (z_out_107[46]))) | ((out_f_d_rsci_q_d[46])
      & (~ (z_out_107[45]))) | ((out_f_d_rsci_q_d[45]) & (~ (z_out_107[44]))) | ((out_f_d_rsci_q_d[44])
      & (~ (z_out_107[43]))) | ((out_f_d_rsci_q_d[43]) & (~ (z_out_107[42]))) | ((out_f_d_rsci_q_d[42])
      & (~ (z_out_107[41]))) | ((out_f_d_rsci_q_d[41]) & (~ (z_out_107[40]))) | ((out_f_d_rsci_q_d[40])
      & (~ (z_out_107[39]))) | ((out_f_d_rsci_q_d[39]) & (~ (z_out_107[38]))) | ((out_f_d_rsci_q_d[38])
      & (~ (z_out_107[37]))) | ((out_f_d_rsci_q_d[37]) & (~ (z_out_107[36]))) | ((out_f_d_rsci_q_d[36])
      & (~ (z_out_107[35]))) | ((out_f_d_rsci_q_d[35]) & (~ (z_out_107[34]))) | ((out_f_d_rsci_q_d[34])
      & (~ (z_out_107[33]))) | ((out_f_d_rsci_q_d[33]) & (~ (z_out_107[32]))) | ((out_f_d_rsci_q_d[32])
      & (~ (z_out_107[31]))) | ((out_f_d_rsci_q_d[31]) & (~ (z_out_107[30]))) | ((out_f_d_rsci_q_d[30])
      & (~ (z_out_107[29]))) | ((out_f_d_rsci_q_d[29]) & (~ (z_out_107[28]))) | ((out_f_d_rsci_q_d[28])
      & (~ (z_out_107[27]))) | ((out_f_d_rsci_q_d[27]) & (~ (z_out_107[26]))) | ((out_f_d_rsci_q_d[26])
      & (~ (z_out_107[25]))) | ((out_f_d_rsci_q_d[25]) & (~ (z_out_107[24]))) | ((out_f_d_rsci_q_d[24])
      & (~ (z_out_107[23]))) | ((out_f_d_rsci_q_d[23]) & (~ (z_out_107[22]))) | ((out_f_d_rsci_q_d[22])
      & (~ (z_out_107[21]))) | ((out_f_d_rsci_q_d[21]) & (~ (z_out_107[20]))) | ((out_f_d_rsci_q_d[20])
      & (~ (z_out_107[19]))) | ((out_f_d_rsci_q_d[19]) & (~ (z_out_107[18]))) | ((out_f_d_rsci_q_d[18])
      & (~ (z_out_107[17]))) | ((out_f_d_rsci_q_d[17]) & (~ (z_out_107[16]))) | ((out_f_d_rsci_q_d[16])
      & (~ (z_out_107[15]))) | ((out_f_d_rsci_q_d[15]) & (~ (z_out_107[14]))) | ((out_f_d_rsci_q_d[14])
      & (~ (z_out_107[13]))) | ((out_f_d_rsci_q_d[13]) & (~ (z_out_107[12]))) | ((out_f_d_rsci_q_d[12])
      & (~ (z_out_107[11]))) | ((out_f_d_rsci_q_d[11]) & (~ (z_out_107[10]))) | ((out_f_d_rsci_q_d[10])
      & (~ (z_out_107[9]))) | ((out_f_d_rsci_q_d[9]) & (~ (z_out_107[8]))) | ((out_f_d_rsci_q_d[8])
      & (~ (z_out_107[7]))) | ((out_f_d_rsci_q_d[7]) & (~ (z_out_107[6]))) | ((out_f_d_rsci_q_d[6])
      & (~ (z_out_107[5]))) | ((out_f_d_rsci_q_d[5]) & (~ (z_out_107[4]))) | ((out_f_d_rsci_q_d[4])
      & (~ (z_out_107[3]))) | ((out_f_d_rsci_q_d[3]) & (~ (z_out_107[2]))) | ((out_f_d_rsci_q_d[2])
      & (~ (z_out_107[1]))) | ((out_f_d_rsci_q_d[1]) & (~ (z_out_107[0]))) | (out_f_d_rsci_q_d[0]);
  assign return_mult_generic_AC_RND_CONV_false_6_mux_12_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_6_if_1_or_1_nl,
      return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_or_1_nl,
      return_mult_generic_AC_RND_CONV_false_6_exp_acc_tmp[11]);
  assign return_mult_generic_AC_RND_CONV_false_6_and_3_nl = (return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1[0])
      & (return_mult_generic_AC_RND_CONV_false_6_mux_12_nl | (return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1[1]));
  assign return_add_generic_AC_RND_CONV_false_1_res_rounded_mux1h_4_nl = MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_1_res_rounded_and_1_nl,
      return_add_generic_AC_RND_CONV_false_7_res_rounded_and_cse, return_mult_generic_AC_RND_CONV_false_6_and_3_nl,
      {return_add_generic_AC_RND_CONV_false_10_r_zero_or_cse , return_add_generic_AC_RND_CONV_false_1_res_rounded_or_2_cse
      , (fsm_output[54])});
  assign nl_z_out_88 = conv_u2u_53_54({return_add_generic_AC_RND_CONV_false_1_res_rounded_return_add_generic_AC_RND_CONV_false_1_res_rounded_and_1_nl
      , return_add_generic_AC_RND_CONV_false_1_res_rounded_mux1h_3_nl}) + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_1_res_rounded_mux1h_4_nl);
  assign z_out_88 = nl_z_out_88[53:0];
  assign return_add_generic_AC_RND_CONV_false_10_res_rounded_return_add_generic_AC_RND_CONV_false_10_res_rounded_mux_3_nl
      = MUX_v_53_2_2((z_out_79[56:4]), (z_out_78[56:4]), BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx0c8);
  assign return_add_generic_AC_RND_CONV_false_12_res_rounded_and_1_nl = (z_out_78[3])
      & ((z_out_78[0]) | (z_out_78[1]) | (z_out_78[2]) | (z_out_78[4]));
  assign return_add_generic_AC_RND_CONV_false_10_res_rounded_return_add_generic_AC_RND_CONV_false_10_res_rounded_mux_4_nl
      = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_res_rounded_and_cse, return_add_generic_AC_RND_CONV_false_12_res_rounded_and_1_nl,
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm_mx0c8);
  assign nl_z_out_89 = conv_u2u_53_54(return_add_generic_AC_RND_CONV_false_10_res_rounded_return_add_generic_AC_RND_CONV_false_10_res_rounded_mux_3_nl)
      + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_10_res_rounded_return_add_generic_AC_RND_CONV_false_10_res_rounded_mux_4_nl);
  assign z_out_89 = nl_z_out_89[53:0];
  assign operator_6_false_3_mux1h_6_nl = MUX1HOT_s_1_6_2(drf_qr_lval_10_smx_lpi_3_dfm_rsp_0,
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0, (operator_14_false_1_acc_psp_sva_9_0[9]),
      (drf_qr_lval_21_smx_9_0_lpi_3_dfm[9]), (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[9]),
      (drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0[8]), {or_tmp_1491 , operator_6_false_3_or_1_ssc
      , operator_6_false_3_or_6_cse , operator_6_false_3_or_8_cse , operator_6_false_3_or_2_cse
      , operator_6_false_3_or_4_cse});
  assign operator_6_false_3_mux1h_7_nl = MUX1HOT_v_8_6_2((drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0[8:1]),
      (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1[9:2]), (operator_14_false_1_acc_psp_sva_9_0[8:1]),
      (drf_qr_lval_21_smx_9_0_lpi_3_dfm[8:1]), (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[8:1]),
      (drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0[7:0]), {or_tmp_1491 , operator_6_false_3_or_1_ssc
      , operator_6_false_3_or_6_cse , operator_6_false_3_or_8_cse , operator_6_false_3_or_2_cse
      , operator_6_false_3_or_4_cse});
  assign operator_6_false_3_mux1h_8_nl = MUX1HOT_s_1_6_2((drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0[0]),
      (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1[1]), (operator_14_false_1_acc_psp_sva_9_0[0]),
      (drf_qr_lval_21_smx_9_0_lpi_3_dfm[0]), (return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0[0]),
      drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1, {or_tmp_1491 , operator_6_false_3_or_1_ssc
      , operator_6_false_3_or_6_cse , operator_6_false_3_or_8_cse , operator_6_false_3_or_2_cse
      , operator_6_false_3_or_4_cse});
  assign operator_6_false_3_or_16_nl = (fsm_output[22]) | (fsm_output[47]);
  assign operator_6_false_3_or_17_nl = (fsm_output[24]) | (fsm_output[49]);
  assign operator_6_false_3_mux1h_9_nl = MUX1HOT_s_1_6_2(drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1,
      (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1[0]), BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm,
      drf_qr_lval_13_smx_0_lpi_3_dfm, drf_qr_lval_14_smx_0_lpi_3_dfm, drf_qr_lval_15_smx_0_lpi_3_dfm,
      {or_tmp_1491 , operator_6_false_3_or_1_ssc , or_tmp_1400 , operator_6_false_3_or_16_nl
      , operator_6_false_3_or_17_nl , operator_6_false_3_or_12_cse});
  assign operator_6_false_3_or_18_nl = or_tmp_1491 | or_tmp_1492 | (fsm_output[22])
      | (fsm_output[45]) | (fsm_output[49]);
  assign operator_6_false_3_or_19_nl = or_dcpl_625 | (fsm_output[24]) | (fsm_output[47]);
  assign operator_6_false_3_mux1h_10_nl = MUX1HOT_v_6_4_2((~ return_add_generic_AC_RND_CONV_false_10_ls_sva),
      (~ return_add_generic_AC_RND_CONV_false_11_ls_sva), (~ return_add_generic_AC_RND_CONV_false_9_ls_sva),
      (~ operator_6_false_17_acc_itm_6_1), {operator_6_false_3_or_18_nl , operator_6_false_3_or_19_nl
      , (fsm_output[20]) , operator_6_false_3_or_12_cse});
  assign nl_acc_29_nl = conv_u2u_12_13({operator_6_false_3_mux1h_6_nl , operator_6_false_3_mux1h_7_nl
      , operator_6_false_3_mux1h_8_nl , operator_6_false_3_mux1h_9_nl , 1'b1}) +
      conv_s2u_8_13({1'b1 , operator_6_false_3_mux1h_10_nl , 1'b1});
  assign acc_29_nl = nl_acc_29_nl[12:0];
  assign z_out_94 = readslicef_13_12_1(acc_29_nl);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif1_return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_3_nl
      = MUX_s_1_2_2(drf_qr_lval_10_smx_lpi_3_dfm_rsp_0, (stage_PE_1_tmp_re_d_sva[62]),
      return_add_generic_AC_RND_CONV_false_6_e_dif1_or_1_cse);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif1_return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_4_nl
      = MUX_v_9_2_2(drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_0, (stage_PE_1_tmp_re_d_sva[61:53]),
      return_add_generic_AC_RND_CONV_false_6_e_dif1_or_1_cse);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif1_return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_5_nl
      = MUX_s_1_2_2(drf_qr_lval_10_smx_lpi_3_dfm_rsp_1_rsp_1, (stage_PE_1_tmp_re_d_sva[52]),
      return_add_generic_AC_RND_CONV_false_6_e_dif1_or_1_cse);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif1_mux1h_5_nl = MUX1HOT_v_10_3_2((~
      drf_qr_lval_10_smx_lpi_3_dfm_mx3_10_1), (~ return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1),
      (~ (in_f_d_rsci_q_d[62:53])), {(fsm_output[11]) , (fsm_output[18]) , return_add_generic_AC_RND_CONV_false_11_or_5_cse});
  assign return_add_generic_AC_RND_CONV_false_6_e_dif1_mux1h_6_nl = MUX1HOT_s_1_3_2((~
      drf_qr_lval_10_smx_lpi_3_dfm_mx3_0), (~ return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1),
      (~ (in_f_d_rsci_q_d[52])), {(fsm_output[11]) , (fsm_output[18]) , return_add_generic_AC_RND_CONV_false_11_or_5_cse});
  assign nl_acc_30_nl = ({1'b1 , return_add_generic_AC_RND_CONV_false_6_e_dif1_return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_3_nl
      , return_add_generic_AC_RND_CONV_false_6_e_dif1_return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_4_nl
      , return_add_generic_AC_RND_CONV_false_6_e_dif1_return_add_generic_AC_RND_CONV_false_6_e_dif1_mux_5_nl
      , 1'b1}) + conv_u2u_12_13({return_add_generic_AC_RND_CONV_false_6_e_dif1_mux1h_5_nl
      , return_add_generic_AC_RND_CONV_false_6_e_dif1_mux1h_6_nl , 1'b1});
  assign acc_30_nl = nl_acc_30_nl[12:0];
  assign z_out_95 = readslicef_13_12_1(acc_30_nl);
  assign return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_or_2_nl
      = (return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3[10]) | (fsm_output[18])
      | (fsm_output[41]);
  assign return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_mux1h_5_nl = MUX1HOT_v_10_3_2((return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3[10:1]),
      return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1, (stage_PE_1_x_re_d_sva[62:53]),
      {(fsm_output[54]) , (fsm_output[18]) , (fsm_output[41])});
  assign return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_mux1h_6_nl = MUX1HOT_s_1_3_2((return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3[0]),
      return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1, (stage_PE_1_x_re_d_sva[52]),
      {(fsm_output[54]) , (fsm_output[18]) , (fsm_output[41])});
  assign return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_or_1_nl = (~ (fsm_output[54]))
      | (fsm_output[18]) | (fsm_output[41]);
  assign return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_mux_2_nl = MUX_v_10_2_2((stage_PE_1_tmp_re_d_sva[62:53]),
      return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1, fsm_output[41]);
  assign return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_nor_1_nl
      = ~(MUX_v_10_2_2(return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_mux_2_nl,
      10'b1111111111, (fsm_output[54])));
  assign return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_mux_3_nl = MUX_s_1_2_2((~
      (stage_PE_1_tmp_re_d_sva[52])), (~ return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1),
      fsm_output[41]);
  assign return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_or_3_nl
      = return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_mux_3_nl | (fsm_output[54]);
  assign nl_acc_31_nl = ({return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_or_2_nl
      , return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_mux1h_5_nl , return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_mux1h_6_nl
      , return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_or_1_nl}) + conv_u2u_12_13({return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_nor_1_nl
      , return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_or_3_nl
      , 1'b1});
  assign acc_31_nl = nl_acc_31_nl[12:0];
  assign z_out_96 = readslicef_13_12_1(acc_31_nl);
  assign stage_u_add_stage_u_add_mux_2_nl = MUX_v_5_2_2(operator_32_false_1_acc_psp_sva_16_12,
      (~ (z_out_111[16:12])), or_1341_cse);
  assign stage_u_add_or_6_nl = MUX_v_5_2_2(stage_u_add_stage_u_add_mux_2_nl, 5'b11111,
      (fsm_output[41]));
  assign stage_u_add_stage_u_add_mux_3_nl = MUX_s_1_2_2((operator_32_false_1_acc_psp_sva_11_0[11]),
      (~ (z_out_111[11])), or_1341_cse);
  assign stage_u_add_or_7_nl = stage_u_add_stage_u_add_mux_3_nl | (fsm_output[41]);
  assign stage_u_add_mux1h_7_nl = MUX1HOT_v_10_3_2((operator_32_false_1_acc_psp_sva_11_0[10:1]),
      (~ (z_out_111[10:1])), return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1,
      {BUTTERFLY_else_or_cse , or_1341_cse , (fsm_output[41])});
  assign stage_u_add_mux1h_8_nl = MUX1HOT_s_1_3_2((operator_32_false_1_acc_psp_sva_11_0[0]),
      (~ (z_out_111[0])), return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1,
      {BUTTERFLY_else_or_cse , or_1341_cse , (fsm_output[41])});
  assign stage_u_add_or_8_nl = (~((fsm_output[6]) | (fsm_output[31]))) | or_1341_cse
      | (fsm_output[41]);
  assign stage_u_add_mux1h_9_nl = MUX1HOT_v_5_3_2((out_u_rsci_q_d[15:11]), (in_u_rsci_q_d[15:11]),
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0, {(fsm_output[6]) , (fsm_output[31])
      , or_1341_cse});
  assign not_1086_nl = ~ (fsm_output[41]);
  assign stage_u_add_and_1_nl = MUX_v_5_2_2(5'b00000, stage_u_add_mux1h_9_nl, not_1086_nl);
  assign stage_u_add_mux1h_10_nl = MUX1HOT_s_1_4_2((out_u_rsci_q_d[10]), (in_u_rsci_q_d[10]),
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0, (~ (stage_PE_1_x_re_d_sva[62])),
      {(fsm_output[6]) , (fsm_output[31]) , or_1341_cse , (fsm_output[41])});
  assign stage_u_add_mux1h_11_nl = MUX1HOT_v_10_4_2((out_u_rsci_q_d[9:0]), (in_u_rsci_q_d[9:0]),
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1, (~ (stage_PE_1_x_re_d_sva[61:52])),
      {(fsm_output[6]) , (fsm_output[31]) , or_1341_cse , (fsm_output[41])});
  assign nl_acc_33_nl = conv_s2u_18_19({stage_u_add_or_6_nl , stage_u_add_or_7_nl
      , stage_u_add_mux1h_7_nl , stage_u_add_mux1h_8_nl , stage_u_add_or_8_nl}) +
      conv_u2u_17_19({stage_u_add_and_1_nl , stage_u_add_mux1h_10_nl , stage_u_add_mux1h_11_nl
      , 1'b1});
  assign acc_33_nl = nl_acc_33_nl[18:0];
  assign z_out_98 = readslicef_19_18_1(acc_33_nl);
  assign BUTTERFLY_BUTTERFLY_or_2_nl = (~((in_u_rsci_q_d[9]) | t_in_or_3_cse)) |
      operator_6_false_33_or_15_cse;
  assign BUTTERFLY_mux_1546_nl = MUX_v_4_2_2((BUTTERFLY_1_n_9_0_sva_8_0[8:5]), (~
      (in_u_rsci_q_d[8:5])), fsm_output[54]);
  assign BUTTERFLY_BUTTERFLY_or_3_nl = MUX_v_4_2_2(BUTTERFLY_mux_1546_nl, 4'b1111,
      operator_6_false_33_or_15_cse);
  assign BUTTERFLY_mux1h_3_nl = MUX1HOT_v_5_3_2((BUTTERFLY_1_n_9_0_sva_8_0[4:0]),
      (~ (in_u_rsci_q_d[4:0])), (~ (return_add_generic_AC_RND_CONV_false_11_ls_sva[5:1])),
      {t_in_or_3_cse , (fsm_output[54]) , operator_6_false_33_or_15_cse});
  assign nl_z_out_101 = ({BUTTERFLY_BUTTERFLY_or_2_nl , BUTTERFLY_BUTTERFLY_or_3_nl
      , BUTTERFLY_mux1h_3_nl}) + 10'b0000000001;
  assign z_out_101 = nl_z_out_101[9:0];
  assign operator_6_false_10_mux_3_nl = MUX_v_10_2_2(drf_qr_lval_21_smx_9_0_lpi_3_dfm,
      operator_14_false_1_acc_psp_sva_9_0, return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse);
  assign nl_z_out_102 = conv_u2u_10_12(operator_6_false_10_mux_3_nl) + conv_s2u_7_12({acc_18_cse_6_1
      , (~ (rtn_out_2[0]))});
  assign z_out_102 = nl_z_out_102[11:0];
  assign operator_33_true_7_or_1_nl = (fsm_output[20]) | (fsm_output[22]) | (fsm_output[24])
      | (fsm_output[26]) | (fsm_output[45]) | (fsm_output[47]) | (fsm_output[49])
      | (fsm_output[51]) | (fsm_output[33]) | (fsm_output[9]);
  assign operator_33_true_7_mux1h_1_nl = MUX1HOT_v_11_3_2((operator_32_false_1_acc_psp_sva_11_0[11:1]),
      (z_out_94[11:1]), (operator_33_true_36_acc_psp_1_sva[11:1]), {(fsm_output[10])
      , operator_33_true_7_or_1_nl , (fsm_output[35])});
  assign nl_z_out_103 = conv_s2u_11_12(operator_33_true_7_mux1h_1_nl) + 12'b000000000001;
  assign z_out_103 = nl_z_out_103[11:0];
  assign BUTTERFLY_i_BUTTERFLY_i_mux_3_nl = MUX_s_1_2_2(BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm,
      return_extract_41_return_extract_41_or_1_cse_sva, return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse);
  assign BUTTERFLY_i_and_5_nl = BUTTERFLY_i_BUTTERFLY_i_mux_3_nl & (~ or_dcpl_198);
  assign BUTTERFLY_i_BUTTERFLY_i_mux_4_nl = MUX_s_1_2_2(stage_PE_1_tmp_im_d_1_lpi_3_dfm_51,
      (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[51]), return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse);
  assign BUTTERFLY_i_and_6_nl = BUTTERFLY_i_BUTTERFLY_i_mux_4_nl & (~ or_dcpl_198);
  assign BUTTERFLY_i_mux_1_nl = MUX_v_42_2_2((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[50:9]),
      (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[50:9]), return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse);
  assign not_1089_nl = ~ or_dcpl_198;
  assign BUTTERFLY_i_BUTTERFLY_i_and_1_nl = MUX_v_42_2_2(42'b000000000000000000000000000000000000000000,
      BUTTERFLY_i_mux_1_nl, not_1089_nl);
  assign BUTTERFLY_i_mux1h_17_nl = MUX1HOT_v_9_3_2(BUTTERFLY_i_div_psp_sva_1, (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[8:0]),
      (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[8:0]), {or_dcpl_198 , operator_14_false_1_or_cse
      , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse});
  assign BUTTERFLY_i_mux1h_18_nl = MUX1HOT_s_1_6_2(return_extract_15_return_extract_15_or_sva_1,
      return_extract_17_return_extract_17_or_sva_1, return_extract_19_return_extract_19_or_sva_1,
      return_extract_47_return_extract_47_or_sva_1, return_extract_49_return_extract_49_or_sva_1,
      return_extract_51_return_extract_51_or_sva_1, {(fsm_output[11]) , (fsm_output[12])
      , (fsm_output[13]) , (fsm_output[36]) , (fsm_output[37]) , (fsm_output[38])});
  assign BUTTERFLY_i_and_7_nl = BUTTERFLY_i_mux1h_18_nl & (~ or_dcpl_198);
  assign BUTTERFLY_i_mux1h_19_nl = MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_4_m_r_51_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0, {or_dcpl_680
      , or_dcpl_484 , (fsm_output[13]) , (fsm_output[38])});
  assign BUTTERFLY_i_and_8_nl = BUTTERFLY_i_mux1h_19_nl & (~ or_dcpl_198);
  assign BUTTERFLY_i_mux1h_20_nl = MUX1HOT_v_41_4_2((return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[50:10]),
      (return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[50:10]), (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[50:10]),
      (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[50:10]), {or_dcpl_680
      , or_dcpl_484 , (fsm_output[13]) , (fsm_output[38])});
  assign not_1092_nl = ~ or_dcpl_198;
  assign BUTTERFLY_i_and_9_nl = MUX_v_41_2_2(41'b00000000000000000000000000000000000000000,
      BUTTERFLY_i_mux1h_20_nl, not_1092_nl);
  assign BUTTERFLY_i_mux1h_21_nl = MUX1HOT_s_1_5_2(stage_PE_1_index_const_9_1_lpi_2_dfm_8,
      (return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[9]), (return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[9]),
      (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[9]), (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[9]),
      {or_dcpl_198 , or_dcpl_680 , or_dcpl_484 , (fsm_output[13]) , (fsm_output[38])});
  assign BUTTERFLY_i_mux1h_22_nl = MUX1HOT_s_1_5_2(stage_PE_1_index_const_9_1_lpi_2_dfm_7,
      (return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[8]), (return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[8]),
      (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[8]), (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[8]),
      {or_dcpl_198 , or_dcpl_680 , or_dcpl_484 , (fsm_output[13]) , (fsm_output[38])});
  assign BUTTERFLY_i_mux1h_23_nl = MUX1HOT_s_1_5_2(stage_PE_1_index_const_9_1_lpi_2_dfm_6,
      (return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[7]), (return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[7]),
      (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[7]), (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[7]),
      {or_dcpl_198 , or_dcpl_680 , or_dcpl_484 , (fsm_output[13]) , (fsm_output[38])});
  assign BUTTERFLY_i_mux1h_24_nl = MUX1HOT_s_1_5_2(stage_PE_1_index_const_9_1_lpi_2_dfm_5,
      (return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[6]), (return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[6]),
      (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[6]), (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[6]),
      {or_dcpl_198 , or_dcpl_680 , or_dcpl_484 , (fsm_output[13]) , (fsm_output[38])});
  assign BUTTERFLY_i_mux1h_25_nl = MUX1HOT_s_1_5_2(stage_PE_1_index_const_9_1_lpi_2_dfm_4,
      (return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[5]), (return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[5]),
      (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[5]), (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[5]),
      {or_dcpl_198 , or_dcpl_680 , or_dcpl_484 , (fsm_output[13]) , (fsm_output[38])});
  assign BUTTERFLY_i_mux1h_26_nl = MUX1HOT_s_1_5_2(stage_PE_1_index_const_9_1_lpi_2_dfm_3,
      (return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[4]), (return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[4]),
      (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[4]), (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[4]),
      {or_dcpl_198 , or_dcpl_680 , or_dcpl_484 , (fsm_output[13]) , (fsm_output[38])});
  assign BUTTERFLY_i_mux1h_27_nl = MUX1HOT_s_1_5_2(stage_PE_1_index_const_9_1_lpi_2_dfm_2,
      (return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[3]), (return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[3]),
      (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[3]), (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[3]),
      {or_dcpl_198 , or_dcpl_680 , or_dcpl_484 , (fsm_output[13]) , (fsm_output[38])});
  assign BUTTERFLY_i_mux1h_28_nl = MUX1HOT_s_1_5_2(stage_PE_1_index_const_9_1_lpi_2_dfm_1,
      (return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[2]), (return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[2]),
      (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[2]), (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[2]),
      {or_dcpl_198 , or_dcpl_680 , or_dcpl_484 , (fsm_output[13]) , (fsm_output[38])});
  assign BUTTERFLY_i_mux1h_29_nl = MUX1HOT_s_1_5_2(stage_PE_1_index_const_9_1_lpi_2_dfm_0,
      (return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[1]), (return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[1]),
      (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[1]), (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[1]),
      {or_dcpl_198 , or_dcpl_680 , or_dcpl_484 , (fsm_output[13]) , (fsm_output[38])});
  assign BUTTERFLY_i_mux1h_30_nl = MUX1HOT_s_1_5_2(stage_PE_1_index_const_0_lpi_2_dfm,
      (return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[0]), (return_add_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[0]),
      (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[0]), (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[0]),
      {or_dcpl_198 , or_dcpl_680 , or_dcpl_484 , (fsm_output[13]) , (fsm_output[38])});
  assign z_out_104 = ({BUTTERFLY_i_and_5_nl , BUTTERFLY_i_and_6_nl , BUTTERFLY_i_BUTTERFLY_i_and_1_nl
      , BUTTERFLY_i_mux1h_17_nl}) * ({BUTTERFLY_i_and_7_nl , BUTTERFLY_i_and_8_nl
      , BUTTERFLY_i_and_9_nl , BUTTERFLY_i_mux1h_21_nl , BUTTERFLY_i_mux1h_22_nl
      , BUTTERFLY_i_mux1h_23_nl , BUTTERFLY_i_mux1h_24_nl , BUTTERFLY_i_mux1h_25_nl
      , BUTTERFLY_i_mux1h_26_nl , BUTTERFLY_i_mux1h_27_nl , BUTTERFLY_i_mux1h_28_nl
      , BUTTERFLY_i_mux1h_29_nl , BUTTERFLY_i_mux1h_30_nl});
  assign BUTTERFLY_else_2_mux_4_nl = MUX_v_14_4_2(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out,
      BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out, BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out,
      BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out, {(fsm_output[31]) ,
      inverse_lpi_1_dfm_1});
  assign BUTTERFLY_else_1_BUTTERFLY_else_1_and_1_nl = MUX_v_2_2_2(2'b00, (z_out_82[17:16]),
      inverse_lpi_1_dfm_1);
  assign BUTTERFLY_else_1_mux_9_nl = MUX_v_5_2_2(BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0,
      (z_out_82[15:11]), inverse_lpi_1_dfm_1);
  assign BUTTERFLY_else_1_mux_10_nl = MUX_s_1_2_2(BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_0,
      (z_out_82[10]), inverse_lpi_1_dfm_1);
  assign BUTTERFLY_else_1_mux_11_nl = MUX_v_10_2_2(BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1,
      (z_out_82[9:0]), inverse_lpi_1_dfm_1);
  assign nl_z_out_105 = $signed(conv_u2s_14_15(BUTTERFLY_else_2_mux_4_nl)) * $signed(({BUTTERFLY_else_1_BUTTERFLY_else_1_and_1_nl
      , BUTTERFLY_else_1_mux_9_nl , BUTTERFLY_else_1_mux_10_nl , BUTTERFLY_else_1_mux_11_nl}));
  assign z_out_105 = nl_z_out_105[31:0];
  assign not_1093_nl = ~ or_1341_cse;
  assign operator_6_false_15_operator_6_false_15_or_2_nl = MUX_v_5_2_2(operator_32_false_1_acc_psp_sva_16_12,
      5'b11111, not_1093_nl);
  assign not_1094_nl = ~ or_1341_cse;
  assign operator_6_false_15_operator_6_false_15_or_3_nl = MUX_v_6_2_2((operator_32_false_1_acc_psp_sva_11_0[11:6]),
      6'b111111, not_1094_nl);
  assign operator_6_false_15_mux_4_nl = MUX_v_6_2_2((~ return_add_generic_AC_RND_CONV_false_10_ls_sva),
      (operator_32_false_1_acc_psp_sva_11_0[5:0]), or_1341_cse);
  assign operator_6_false_15_or_1_nl = (~ or_1341_cse) | (fsm_output[37]) | (fsm_output[38])
      | (fsm_output[39]) | (fsm_output[14]) | (fsm_output[13]) | (fsm_output[12]);
  assign operator_6_false_15_mux_5_nl = MUX_s_1_2_2((operator_14_false_1_acc_psp_sva_12_10[2]),
      (operator_32_false_1_acc_psp_sva_16_12[4]), or_1341_cse);
  assign not_1096_nl = ~ or_1341_cse;
  assign operator_6_false_15_operator_6_false_15_and_2_nl = MUX_v_2_2_2(2'b00, (operator_14_false_1_acc_psp_sva_12_10[1:0]),
      not_1096_nl);
  assign not_1097_nl = ~ or_1341_cse;
  assign operator_6_false_15_operator_6_false_15_and_3_nl = MUX_v_9_2_2(9'b000000000,
      (operator_14_false_1_acc_psp_sva_9_0[9:1]), not_1097_nl);
  assign operator_6_false_15_mux_6_nl = MUX_s_1_2_2((operator_14_false_1_acc_psp_sva_9_0[0]),
      (operator_32_false_1_acc_psp_sva_16_12[4]), or_1341_cse);
  assign nl_acc_39_nl = ({operator_6_false_15_operator_6_false_15_or_2_nl , operator_6_false_15_operator_6_false_15_or_3_nl
      , operator_6_false_15_mux_4_nl , operator_6_false_15_or_1_nl}) + conv_u2u_15_18(signext_15_14({operator_6_false_15_mux_5_nl
      , operator_6_false_15_operator_6_false_15_and_2_nl , operator_6_false_15_operator_6_false_15_and_3_nl
      , operator_6_false_15_mux_6_nl , 1'b1}));
  assign acc_39_nl = nl_acc_39_nl[17:0];
  assign z_out_111 = readslicef_18_17_1(acc_39_nl);
  assign operator_33_true_11_mux_1_nl = MUX_v_10_2_2((operator_6_false_11_acc_psp_1_sva_1[10:1]),
      (operator_6_false_9_acc_psp_1_sva_1[10:1]), return_add_generic_AC_RND_CONV_false_17_e_dif_sat_or_cse);
  assign nl_z_out_112 = conv_s2u_10_11(operator_33_true_11_mux_1_nl) + 11'b00000000001;
  assign z_out_112 = nl_z_out_112[10:0];
  assign operator_32_false_2_operator_32_false_2_and_1_nl = (operator_32_false_2_acc_5_itm[10])
      & (~ (fsm_output[55]));
  assign operator_32_false_2_mux_3_nl = MUX_v_10_2_2((operator_32_false_2_acc_5_itm[9:0]),
      return_add_generic_AC_RND_CONV_false_19_exp_plus_1_12_1_lpi_3_dfm_9_0, fsm_output[55]);
  assign nl_z_out_113 = ({operator_32_false_2_operator_32_false_2_and_1_nl , operator_32_false_2_mux_3_nl})
      + ({(~ (fsm_output[55])) , 10'b0000000001});
  assign z_out_113 = nl_z_out_113[10:0];
  assign nl_z_out_114 = conv_s2u_11_12(z_out_94[11:1]) + 12'b000000000001;
  assign z_out_114 = nl_z_out_114[11:0];
  assign z_out_13 = MUX1HOT_s_1_3_2((z_out_106[53]), (z_out_106[52]), reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd_52,
      {return_mult_generic_AC_RND_CONV_false_mux1h_cse , return_mult_generic_AC_RND_CONV_false_mux1h_1_cse
      , (operator_14_false_1_acc_psp_sva_12_10[2])});
  assign z_out_90 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_11,
      (return_add_generic_AC_RND_CONV_false_1_return_add_generic_AC_RND_CONV_false_1_and_5_cse[9:0]),
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_4_or_8_tmp = (fsm_output[12]) | (fsm_output[36]);
  assign return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_4_or_8_tmp | (z_out_89[53]));
  assign return_add_generic_AC_RND_CONV_false_4_and_1_nl = return_add_generic_AC_RND_CONV_false_4_or_8_tmp
      & (~ (z_out_89[53]));
  assign return_add_generic_AC_RND_CONV_false_4_and_2_nl = (~ or_dcpl_484) & (z_out_89[53]);
  assign return_add_generic_AC_RND_CONV_false_4_and_3_nl = or_dcpl_484 & (z_out_89[53]);
  assign z_out_91 = MUX1HOT_v_10_4_2((operator_33_true_36_acc_psp_1_sva[10:1]), (operator_32_false_1_acc_psp_sva_11_0[10:1]),
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1_rsp_1, (drf_qr_lval_19_smx_lpi_3_dfm[9:0]),
      {return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_nor_nl
      , return_add_generic_AC_RND_CONV_false_4_and_1_nl , return_add_generic_AC_RND_CONV_false_4_and_2_nl
      , return_add_generic_AC_RND_CONV_false_4_and_3_nl});
  function automatic [8:0] div_9_u9_u16;
    input [8:0] l;
    input [15:0] r;
    reg [8:0] rdiv;
    reg [16:0] diff;
    reg [17:0] diff_tmp;
    reg [24:0] lbuf;
    integer i;
  begin
    lbuf = 25'b0;
    lbuf[8:0] = l;
    for(i=8; i>=0; i=i-1)
    begin
      diff_tmp = (lbuf[24:8] - {1'b0,r});
      diff = diff_tmp[16:0];
      rdiv[i] = ~diff[16];
      if(diff[16] == 0)
        lbuf[24:8] = diff;
      lbuf[24:1] = lbuf[23:0];
    end
    div_9_u9_u16 = rdiv;
  end
  endfunction
  function automatic MUX1HOT_s_1_10_2;
    input input_9;
    input input_8;
    input input_7;
    input input_6;
    input input_5;
    input input_4;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [9:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    MUX1HOT_s_1_10_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_11_2;
    input input_10;
    input input_9;
    input input_8;
    input input_7;
    input input_6;
    input input_5;
    input input_4;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [10:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    MUX1HOT_s_1_11_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_12_2;
    input input_11;
    input input_10;
    input input_9;
    input input_8;
    input input_7;
    input input_6;
    input input_5;
    input input_4;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [11:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    MUX1HOT_s_1_12_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_13_2;
    input input_12;
    input input_11;
    input input_10;
    input input_9;
    input input_8;
    input input_7;
    input input_6;
    input input_5;
    input input_4;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [12:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    MUX1HOT_s_1_13_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_14_2;
    input input_13;
    input input_12;
    input input_11;
    input input_10;
    input input_9;
    input input_8;
    input input_7;
    input input_6;
    input input_5;
    input input_4;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [13:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    MUX1HOT_s_1_14_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_15_2;
    input input_14;
    input input_13;
    input input_12;
    input input_11;
    input input_10;
    input input_9;
    input input_8;
    input input_7;
    input input_6;
    input input_5;
    input input_4;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [14:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    MUX1HOT_s_1_15_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_16_2;
    input input_15;
    input input_14;
    input input_13;
    input input_12;
    input input_11;
    input input_10;
    input input_9;
    input input_8;
    input input_7;
    input input_6;
    input input_5;
    input input_4;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [15:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    MUX1HOT_s_1_16_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_20_2;
    input input_19;
    input input_18;
    input input_17;
    input input_16;
    input input_15;
    input input_14;
    input input_13;
    input input_12;
    input input_11;
    input input_10;
    input input_9;
    input input_8;
    input input_7;
    input input_6;
    input input_5;
    input input_4;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [19:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    result = result | (input_18 & sel[18]);
    result = result | (input_19 & sel[19]);
    MUX1HOT_s_1_20_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_21_2;
    input input_20;
    input input_19;
    input input_18;
    input input_17;
    input input_16;
    input input_15;
    input input_14;
    input input_13;
    input input_12;
    input input_11;
    input input_10;
    input input_9;
    input input_8;
    input input_7;
    input input_6;
    input input_5;
    input input_4;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [20:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    result = result | (input_18 & sel[18]);
    result = result | (input_19 & sel[19]);
    result = result | (input_20 & sel[20]);
    MUX1HOT_s_1_21_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_3_2;
    input input_2;
    input input_1;
    input input_0;
    input [2:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_4_2;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [3:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_5_2;
    input input_4;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [4:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_6_2;
    input input_5;
    input input_4;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [5:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_7_2;
    input input_6;
    input input_5;
    input input_4;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [6:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_8_2;
    input input_7;
    input input_6;
    input input_5;
    input input_4;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [7:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    MUX1HOT_s_1_8_2 = result;
  end
  endfunction
  function automatic MUX1HOT_s_1_9_2;
    input input_8;
    input input_7;
    input input_6;
    input input_5;
    input input_4;
    input input_3;
    input input_2;
    input input_1;
    input input_0;
    input [8:0] sel;
    reg result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    MUX1HOT_s_1_9_2 = result;
  end
  endfunction
  function automatic [9:0] MUX1HOT_v_10_12_2;
    input [9:0] input_11;
    input [9:0] input_10;
    input [9:0] input_9;
    input [9:0] input_8;
    input [9:0] input_7;
    input [9:0] input_6;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [11:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    result = result | (input_3 & {10{sel[3]}});
    result = result | (input_4 & {10{sel[4]}});
    result = result | (input_5 & {10{sel[5]}});
    result = result | (input_6 & {10{sel[6]}});
    result = result | (input_7 & {10{sel[7]}});
    result = result | (input_8 & {10{sel[8]}});
    result = result | (input_9 & {10{sel[9]}});
    result = result | (input_10 & {10{sel[10]}});
    result = result | (input_11 & {10{sel[11]}});
    MUX1HOT_v_10_12_2 = result;
  end
  endfunction
  function automatic [9:0] MUX1HOT_v_10_3_2;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [2:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    MUX1HOT_v_10_3_2 = result;
  end
  endfunction
  function automatic [9:0] MUX1HOT_v_10_4_2;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [3:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    result = result | (input_3 & {10{sel[3]}});
    MUX1HOT_v_10_4_2 = result;
  end
  endfunction
  function automatic [9:0] MUX1HOT_v_10_5_2;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [4:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    result = result | (input_3 & {10{sel[3]}});
    result = result | (input_4 & {10{sel[4]}});
    MUX1HOT_v_10_5_2 = result;
  end
  endfunction
  function automatic [9:0] MUX1HOT_v_10_6_2;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [5:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    result = result | (input_3 & {10{sel[3]}});
    result = result | (input_4 & {10{sel[4]}});
    result = result | (input_5 & {10{sel[5]}});
    MUX1HOT_v_10_6_2 = result;
  end
  endfunction
  function automatic [9:0] MUX1HOT_v_10_7_2;
    input [9:0] input_6;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [6:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    result = result | (input_3 & {10{sel[3]}});
    result = result | (input_4 & {10{sel[4]}});
    result = result | (input_5 & {10{sel[5]}});
    result = result | (input_6 & {10{sel[6]}});
    MUX1HOT_v_10_7_2 = result;
  end
  endfunction
  function automatic [10:0] MUX1HOT_v_11_3_2;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [2:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    MUX1HOT_v_11_3_2 = result;
  end
  endfunction
  function automatic [10:0] MUX1HOT_v_11_4_2;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [3:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    result = result | (input_3 & {11{sel[3]}});
    MUX1HOT_v_11_4_2 = result;
  end
  endfunction
  function automatic [11:0] MUX1HOT_v_12_4_2;
    input [11:0] input_3;
    input [11:0] input_2;
    input [11:0] input_1;
    input [11:0] input_0;
    input [3:0] sel;
    reg [11:0] result;
  begin
    result = input_0 & {12{sel[0]}};
    result = result | (input_1 & {12{sel[1]}});
    result = result | (input_2 & {12{sel[2]}});
    result = result | (input_3 & {12{sel[3]}});
    MUX1HOT_v_12_4_2 = result;
  end
  endfunction
  function automatic [12:0] MUX1HOT_v_13_4_2;
    input [12:0] input_3;
    input [12:0] input_2;
    input [12:0] input_1;
    input [12:0] input_0;
    input [3:0] sel;
    reg [12:0] result;
  begin
    result = input_0 & {13{sel[0]}};
    result = result | (input_1 & {13{sel[1]}});
    result = result | (input_2 & {13{sel[2]}});
    result = result | (input_3 & {13{sel[3]}});
    MUX1HOT_v_13_4_2 = result;
  end
  endfunction
  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction
  function automatic [15:0] MUX1HOT_v_16_4_2;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [3:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    MUX1HOT_v_16_4_2 = result;
  end
  endfunction
  function automatic [1:0] MUX1HOT_v_2_8_2;
    input [1:0] input_7;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [7:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    result = result | (input_7 & {2{sel[7]}});
    MUX1HOT_v_2_8_2 = result;
  end
  endfunction
  function automatic [2:0] MUX1HOT_v_3_11_2;
    input [2:0] input_10;
    input [2:0] input_9;
    input [2:0] input_8;
    input [2:0] input_7;
    input [2:0] input_6;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [10:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    result = result | (input_5 & {3{sel[5]}});
    result = result | (input_6 & {3{sel[6]}});
    result = result | (input_7 & {3{sel[7]}});
    result = result | (input_8 & {3{sel[8]}});
    result = result | (input_9 & {3{sel[9]}});
    result = result | (input_10 & {3{sel[10]}});
    MUX1HOT_v_3_11_2 = result;
  end
  endfunction
  function automatic [40:0] MUX1HOT_v_41_4_2;
    input [40:0] input_3;
    input [40:0] input_2;
    input [40:0] input_1;
    input [40:0] input_0;
    input [3:0] sel;
    reg [40:0] result;
  begin
    result = input_0 & {41{sel[0]}};
    result = result | (input_1 & {41{sel[1]}});
    result = result | (input_2 & {41{sel[2]}});
    result = result | (input_3 & {41{sel[3]}});
    MUX1HOT_v_41_4_2 = result;
  end
  endfunction
  function automatic [3:0] MUX1HOT_v_4_14_2;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [13:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    MUX1HOT_v_4_14_2 = result;
  end
  endfunction
  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction
  function automatic [3:0] MUX1HOT_v_4_8_2;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [7:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    MUX1HOT_v_4_8_2 = result;
  end
  endfunction
  function automatic [49:0] MUX1HOT_v_50_10_2;
    input [49:0] input_9;
    input [49:0] input_8;
    input [49:0] input_7;
    input [49:0] input_6;
    input [49:0] input_5;
    input [49:0] input_4;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [9:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    result = result | (input_3 & {50{sel[3]}});
    result = result | (input_4 & {50{sel[4]}});
    result = result | (input_5 & {50{sel[5]}});
    result = result | (input_6 & {50{sel[6]}});
    result = result | (input_7 & {50{sel[7]}});
    result = result | (input_8 & {50{sel[8]}});
    result = result | (input_9 & {50{sel[9]}});
    MUX1HOT_v_50_10_2 = result;
  end
  endfunction
  function automatic [49:0] MUX1HOT_v_50_12_2;
    input [49:0] input_11;
    input [49:0] input_10;
    input [49:0] input_9;
    input [49:0] input_8;
    input [49:0] input_7;
    input [49:0] input_6;
    input [49:0] input_5;
    input [49:0] input_4;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [11:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    result = result | (input_3 & {50{sel[3]}});
    result = result | (input_4 & {50{sel[4]}});
    result = result | (input_5 & {50{sel[5]}});
    result = result | (input_6 & {50{sel[6]}});
    result = result | (input_7 & {50{sel[7]}});
    result = result | (input_8 & {50{sel[8]}});
    result = result | (input_9 & {50{sel[9]}});
    result = result | (input_10 & {50{sel[10]}});
    result = result | (input_11 & {50{sel[11]}});
    MUX1HOT_v_50_12_2 = result;
  end
  endfunction
  function automatic [49:0] MUX1HOT_v_50_5_2;
    input [49:0] input_4;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [4:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    result = result | (input_3 & {50{sel[3]}});
    result = result | (input_4 & {50{sel[4]}});
    MUX1HOT_v_50_5_2 = result;
  end
  endfunction
  function automatic [49:0] MUX1HOT_v_50_7_2;
    input [49:0] input_6;
    input [49:0] input_5;
    input [49:0] input_4;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [6:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    result = result | (input_3 & {50{sel[3]}});
    result = result | (input_4 & {50{sel[4]}});
    result = result | (input_5 & {50{sel[5]}});
    result = result | (input_6 & {50{sel[6]}});
    MUX1HOT_v_50_7_2 = result;
  end
  endfunction
  function automatic [49:0] MUX1HOT_v_50_8_2;
    input [49:0] input_7;
    input [49:0] input_6;
    input [49:0] input_5;
    input [49:0] input_4;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [7:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    result = result | (input_3 & {50{sel[3]}});
    result = result | (input_4 & {50{sel[4]}});
    result = result | (input_5 & {50{sel[5]}});
    result = result | (input_6 & {50{sel[6]}});
    result = result | (input_7 & {50{sel[7]}});
    MUX1HOT_v_50_8_2 = result;
  end
  endfunction
  function automatic [50:0] MUX1HOT_v_51_3_2;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [2:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | (input_1 & {51{sel[1]}});
    result = result | (input_2 & {51{sel[2]}});
    MUX1HOT_v_51_3_2 = result;
  end
  endfunction
  function automatic [50:0] MUX1HOT_v_51_4_2;
    input [50:0] input_3;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [3:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | (input_1 & {51{sel[1]}});
    result = result | (input_2 & {51{sel[2]}});
    result = result | (input_3 & {51{sel[3]}});
    MUX1HOT_v_51_4_2 = result;
  end
  endfunction
  function automatic [50:0] MUX1HOT_v_51_5_2;
    input [50:0] input_4;
    input [50:0] input_3;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [4:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | (input_1 & {51{sel[1]}});
    result = result | (input_2 & {51{sel[2]}});
    result = result | (input_3 & {51{sel[3]}});
    result = result | (input_4 & {51{sel[4]}});
    MUX1HOT_v_51_5_2 = result;
  end
  endfunction
  function automatic [50:0] MUX1HOT_v_51_6_2;
    input [50:0] input_5;
    input [50:0] input_4;
    input [50:0] input_3;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [5:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | (input_1 & {51{sel[1]}});
    result = result | (input_2 & {51{sel[2]}});
    result = result | (input_3 & {51{sel[3]}});
    result = result | (input_4 & {51{sel[4]}});
    result = result | (input_5 & {51{sel[5]}});
    MUX1HOT_v_51_6_2 = result;
  end
  endfunction
  function automatic [50:0] MUX1HOT_v_51_7_2;
    input [50:0] input_6;
    input [50:0] input_5;
    input [50:0] input_4;
    input [50:0] input_3;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [6:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | (input_1 & {51{sel[1]}});
    result = result | (input_2 & {51{sel[2]}});
    result = result | (input_3 & {51{sel[3]}});
    result = result | (input_4 & {51{sel[4]}});
    result = result | (input_5 & {51{sel[5]}});
    result = result | (input_6 & {51{sel[6]}});
    MUX1HOT_v_51_7_2 = result;
  end
  endfunction
  function automatic [51:0] MUX1HOT_v_52_3_2;
    input [51:0] input_2;
    input [51:0] input_1;
    input [51:0] input_0;
    input [2:0] sel;
    reg [51:0] result;
  begin
    result = input_0 & {52{sel[0]}};
    result = result | (input_1 & {52{sel[1]}});
    result = result | (input_2 & {52{sel[2]}});
    MUX1HOT_v_52_3_2 = result;
  end
  endfunction
  function automatic [52:0] MUX1HOT_v_53_3_2;
    input [52:0] input_2;
    input [52:0] input_1;
    input [52:0] input_0;
    input [2:0] sel;
    reg [52:0] result;
  begin
    result = input_0 & {53{sel[0]}};
    result = result | (input_1 & {53{sel[1]}});
    result = result | (input_2 & {53{sel[2]}});
    MUX1HOT_v_53_3_2 = result;
  end
  endfunction
  function automatic [55:0] MUX1HOT_v_56_3_2;
    input [55:0] input_2;
    input [55:0] input_1;
    input [55:0] input_0;
    input [2:0] sel;
    reg [55:0] result;
  begin
    result = input_0 & {56{sel[0]}};
    result = result | (input_1 & {56{sel[1]}});
    result = result | (input_2 & {56{sel[2]}});
    MUX1HOT_v_56_3_2 = result;
  end
  endfunction
  function automatic [55:0] MUX1HOT_v_56_4_2;
    input [55:0] input_3;
    input [55:0] input_2;
    input [55:0] input_1;
    input [55:0] input_0;
    input [3:0] sel;
    reg [55:0] result;
  begin
    result = input_0 & {56{sel[0]}};
    result = result | (input_1 & {56{sel[1]}});
    result = result | (input_2 & {56{sel[2]}});
    result = result | (input_3 & {56{sel[3]}});
    MUX1HOT_v_56_4_2 = result;
  end
  endfunction
  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction
  function automatic [4:0] MUX1HOT_v_5_7_2;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [6:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    MUX1HOT_v_5_7_2 = result;
  end
  endfunction
  function automatic [4:0] MUX1HOT_v_5_8_2;
    input [4:0] input_7;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [7:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    result = result | (input_7 & {5{sel[7]}});
    MUX1HOT_v_5_8_2 = result;
  end
  endfunction
  function automatic [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction
  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction
  function automatic [5:0] MUX1HOT_v_6_5_2;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [4:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    MUX1HOT_v_6_5_2 = result;
  end
  endfunction
  function automatic [5:0] MUX1HOT_v_6_9_2;
    input [5:0] input_8;
    input [5:0] input_7;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [8:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    result = result | (input_6 & {6{sel[6]}});
    result = result | (input_7 & {6{sel[7]}});
    result = result | (input_8 & {6{sel[8]}});
    MUX1HOT_v_6_9_2 = result;
  end
  endfunction
  function automatic [7:0] MUX1HOT_v_8_6_2;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [5:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    MUX1HOT_v_8_6_2 = result;
  end
  endfunction
  function automatic [8:0] MUX1HOT_v_9_13_2;
    input [8:0] input_12;
    input [8:0] input_11;
    input [8:0] input_10;
    input [8:0] input_9;
    input [8:0] input_8;
    input [8:0] input_7;
    input [8:0] input_6;
    input [8:0] input_5;
    input [8:0] input_4;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [12:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | (input_1 & {9{sel[1]}});
    result = result | (input_2 & {9{sel[2]}});
    result = result | (input_3 & {9{sel[3]}});
    result = result | (input_4 & {9{sel[4]}});
    result = result | (input_5 & {9{sel[5]}});
    result = result | (input_6 & {9{sel[6]}});
    result = result | (input_7 & {9{sel[7]}});
    result = result | (input_8 & {9{sel[8]}});
    result = result | (input_9 & {9{sel[9]}});
    result = result | (input_10 & {9{sel[10]}});
    result = result | (input_11 & {9{sel[11]}});
    result = result | (input_12 & {9{sel[12]}});
    MUX1HOT_v_9_13_2 = result;
  end
  endfunction
  function automatic [8:0] MUX1HOT_v_9_3_2;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [2:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | (input_1 & {9{sel[1]}});
    result = result | (input_2 & {9{sel[2]}});
    MUX1HOT_v_9_3_2 = result;
  end
  endfunction
  function automatic [8:0] MUX1HOT_v_9_4_2;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [3:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | (input_1 & {9{sel[1]}});
    result = result | (input_2 & {9{sel[2]}});
    result = result | (input_3 & {9{sel[3]}});
    MUX1HOT_v_9_4_2 = result;
  end
  endfunction
  function automatic [8:0] MUX1HOT_v_9_5_2;
    input [8:0] input_4;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [4:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | (input_1 & {9{sel[1]}});
    result = result | (input_2 & {9{sel[2]}});
    result = result | (input_3 & {9{sel[3]}});
    result = result | (input_4 & {9{sel[4]}});
    MUX1HOT_v_9_5_2 = result;
  end
  endfunction
  function automatic [8:0] MUX1HOT_v_9_9_2;
    input [8:0] input_8;
    input [8:0] input_7;
    input [8:0] input_6;
    input [8:0] input_5;
    input [8:0] input_4;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [8:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | (input_1 & {9{sel[1]}});
    result = result | (input_2 & {9{sel[2]}});
    result = result | (input_3 & {9{sel[3]}});
    result = result | (input_4 & {9{sel[4]}});
    result = result | (input_5 & {9{sel[5]}});
    result = result | (input_6 & {9{sel[6]}});
    result = result | (input_7 & {9{sel[7]}});
    result = result | (input_8 & {9{sel[8]}});
    MUX1HOT_v_9_9_2 = result;
  end
  endfunction
  function automatic MUX_s_1_2_2;
    input input_0;
    input input_1;
    input sel;
    reg result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction
  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction
  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction
  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction
  function automatic [13:0] MUX_v_14_4_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [13:0] input_2;
    input [13:0] input_3;
    input [1:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_14_4_2 = result;
  end
  endfunction
  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction
  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction
  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction
  function automatic [40:0] MUX_v_41_2_2;
    input [40:0] input_0;
    input [40:0] input_1;
    input sel;
    reg [40:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_41_2_2 = result;
  end
  endfunction
  function automatic [41:0] MUX_v_42_2_2;
    input [41:0] input_0;
    input [41:0] input_1;
    input sel;
    reg [41:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_42_2_2 = result;
  end
  endfunction
  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction
  function automatic [49:0] MUX_v_50_2_2;
    input [49:0] input_0;
    input [49:0] input_1;
    input sel;
    reg [49:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_50_2_2 = result;
  end
  endfunction
  function automatic [50:0] MUX_v_51_2_2;
    input [50:0] input_0;
    input [50:0] input_1;
    input sel;
    reg [50:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_51_2_2 = result;
  end
  endfunction
  function automatic [51:0] MUX_v_52_2_2;
    input [51:0] input_0;
    input [51:0] input_1;
    input sel;
    reg [51:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_52_2_2 = result;
  end
  endfunction
  function automatic [52:0] MUX_v_53_2_2;
    input [52:0] input_0;
    input [52:0] input_1;
    input sel;
    reg [52:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_53_2_2 = result;
  end
  endfunction
  function automatic [55:0] MUX_v_56_2_2;
    input [55:0] input_0;
    input [55:0] input_1;
    input sel;
    reg [55:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_56_2_2 = result;
  end
  endfunction
  function automatic [56:0] MUX_v_57_2_2;
    input [56:0] input_0;
    input [56:0] input_1;
    input sel;
    reg [56:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_57_2_2 = result;
  end
  endfunction
  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction
  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction
  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction
  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction
  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction
  function automatic [0:0] readslicef_12_1_11;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_12_1_11 = tmp[0:0];
  end
  endfunction
  function automatic [11:0] readslicef_13_12_1;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_13_12_1 = tmp[11:0];
  end
  endfunction
  function automatic [0:0] readslicef_13_1_12;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 12;
    readslicef_13_1_12 = tmp[0:0];
  end
  endfunction
  function automatic [12:0] readslicef_14_13_1;
    input [13:0] vector;
    reg [13:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_14_13_1 = tmp[12:0];
  end
  endfunction
  function automatic [16:0] readslicef_18_17_1;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_18_17_1 = tmp[16:0];
  end
  endfunction
  function automatic [17:0] readslicef_19_18_1;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_19_18_1 = tmp[17:0];
  end
  endfunction
  function automatic [13:0] readslicef_24_14_10;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_24_14_10 = tmp[13:0];
  end
  endfunction
  function automatic [15:0] readslicef_32_16_16;
    input [31:0] vector;
    reg [31:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_32_16_16 = tmp[15:0];
  end
  endfunction
  function automatic [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction
  function automatic [0:0] readslicef_53_1_52;
    input [52:0] vector;
    reg [52:0] tmp;
  begin
    tmp = vector >> 52;
    readslicef_53_1_52 = tmp[0:0];
  end
  endfunction
  function automatic [0:0] readslicef_54_1_53;
    input [53:0] vector;
    reg [53:0] tmp;
  begin
    tmp = vector >> 53;
    readslicef_54_1_53 = tmp[0:0];
  end
  endfunction
  function automatic [56:0] readslicef_58_57_1;
    input [57:0] vector;
    reg [57:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_58_57_1 = tmp[56:0];
  end
  endfunction
  function automatic [9:0] signext_10_1;
    input vector;
  begin
    signext_10_1= {{9{vector}}, vector};
  end
  endfunction
  function automatic [13:0] signext_14_13;
    input [12:0] vector;
  begin
    signext_14_13= {{1{vector[12]}}, vector};
  end
  endfunction
  function automatic [14:0] signext_15_14;
    input [13:0] vector;
  begin
    signext_15_14= {{1{vector[13]}}, vector};
  end
  endfunction
  function automatic [15:0] signext_16_14;
    input [13:0] vector;
  begin
    signext_16_14= {{2{vector[13]}}, vector};
  end
  endfunction
  function automatic [1:0] signext_2_1;
    input vector;
  begin
    signext_2_1= {{1{vector}}, vector};
  end
  endfunction
  function automatic [54:0] signext_55_54;
    input [53:0] vector;
  begin
    signext_55_54= {{1{vector[53]}}, vector};
  end
  endfunction
  function automatic [11:0] conv_s2s_5_12 ;
    input [4:0] vector ;
  begin
    conv_s2s_5_12 = {{7{vector[4]}}, vector};
  end
  endfunction
  function automatic [10:0] conv_s2s_7_11 ;
    input [6:0] vector ;
  begin
    conv_s2s_7_11 = {{4{vector[6]}}, vector};
  end
  endfunction
  function automatic [11:0] conv_s2s_7_12 ;
    input [6:0] vector ;
  begin
    conv_s2s_7_12 = {{5{vector[6]}}, vector};
  end
  endfunction
  function automatic [12:0] conv_s2s_7_13 ;
    input [6:0] vector ;
  begin
    conv_s2s_7_13 = {{6{vector[6]}}, vector};
  end
  endfunction
  function automatic [11:0] conv_s2s_11_12 ;
    input [10:0] vector ;
  begin
    conv_s2s_11_12 = {vector[10], vector};
  end
  endfunction
  function automatic [17:0] conv_s2s_17_18 ;
    input [16:0] vector ;
  begin
    conv_s2s_17_18 = {vector[16], vector};
  end
  endfunction
  function automatic [11:0] conv_s2u_7_12 ;
    input [6:0] vector ;
  begin
    conv_s2u_7_12 = {{5{vector[6]}}, vector};
  end
  endfunction
  function automatic [12:0] conv_s2u_7_13 ;
    input [6:0] vector ;
  begin
    conv_s2u_7_13 = {{6{vector[6]}}, vector};
  end
  endfunction
  function automatic [12:0] conv_s2u_8_13 ;
    input [7:0] vector ;
  begin
    conv_s2u_8_13 = {{5{vector[7]}}, vector};
  end
  endfunction
  function automatic [10:0] conv_s2u_10_11 ;
    input [9:0] vector ;
  begin
    conv_s2u_10_11 = {vector[9], vector};
  end
  endfunction
  function automatic [11:0] conv_s2u_11_12 ;
    input [10:0] vector ;
  begin
    conv_s2u_11_12 = {vector[10], vector};
  end
  endfunction
  function automatic [12:0] conv_s2u_12_13 ;
    input [11:0] vector ;
  begin
    conv_s2u_12_13 = {vector[11], vector};
  end
  endfunction
  function automatic [13:0] conv_s2u_12_14 ;
    input [11:0] vector ;
  begin
    conv_s2u_12_14 = {{2{vector[11]}}, vector};
  end
  endfunction
  function automatic [13:0] conv_s2u_13_14 ;
    input [12:0] vector ;
  begin
    conv_s2u_13_14 = {vector[12], vector};
  end
  endfunction
  function automatic [17:0] conv_s2u_17_18 ;
    input [16:0] vector ;
  begin
    conv_s2u_17_18 = {vector[16], vector};
  end
  endfunction
  function automatic [18:0] conv_s2u_18_19 ;
    input [17:0] vector ;
  begin
    conv_s2u_18_19 = {vector[17], vector};
  end
  endfunction
  function automatic [23:0] conv_s2u_23_24 ;
    input [22:0] vector ;
  begin
    conv_s2u_23_24 = {vector[22], vector};
  end
  endfunction
  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0] vector ;
  begin
    conv_u2s_3_4 = {1'b0, vector};
  end
  endfunction
  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0] vector ;
  begin
    conv_u2s_10_11 = {1'b0, vector};
  end
  endfunction
  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0] vector ;
  begin
    conv_u2s_11_12 = {1'b0, vector};
  end
  endfunction
  function automatic [12:0] conv_u2s_11_13 ;
    input [10:0] vector ;
  begin
    conv_u2s_11_13 = {{2{1'b0}}, vector};
  end
  endfunction
  function automatic [14:0] conv_u2s_14_15 ;
    input [13:0] vector ;
  begin
    conv_u2s_14_15 = {1'b0, vector};
  end
  endfunction
  function automatic [16:0] conv_u2s_16_17 ;
    input [15:0] vector ;
  begin
    conv_u2s_16_17 = {1'b0, vector};
  end
  endfunction
  function automatic [51:0] conv_u2u_1_52 ;
    input [0:0] vector ;
  begin
    conv_u2u_1_52 = {{51{1'b0}}, vector};
  end
  endfunction
  function automatic [53:0] conv_u2u_1_54 ;
    input [0:0] vector ;
  begin
    conv_u2u_1_54 = {{53{1'b0}}, vector};
  end
  endfunction
  function automatic [12:0] conv_u2u_2_13 ;
    input [1:0] vector ;
  begin
    conv_u2u_2_13 = {{11{1'b0}}, vector};
  end
  endfunction
  function automatic [10:0] conv_u2u_4_11 ;
    input [3:0] vector ;
  begin
    conv_u2u_4_11 = {{7{1'b0}}, vector};
  end
  endfunction
  function automatic [15:0] conv_u2u_4_16 ;
    input [3:0] vector ;
  begin
    conv_u2u_4_16 = {{12{1'b0}}, vector};
  end
  endfunction
  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0] vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction
  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0] vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction
  function automatic [11:0] conv_u2u_10_12 ;
    input [9:0] vector ;
  begin
    conv_u2u_10_12 = {{2{1'b0}}, vector};
  end
  endfunction
  function automatic [11:0] conv_u2u_11_12 ;
    input [10:0] vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction
  function automatic [12:0] conv_u2u_11_13 ;
    input [10:0] vector ;
  begin
    conv_u2u_11_13 = {{2{1'b0}}, vector};
  end
  endfunction
  function automatic [12:0] conv_u2u_12_13 ;
    input [11:0] vector ;
  begin
    conv_u2u_12_13 = {1'b0, vector};
  end
  endfunction
  function automatic [13:0] conv_u2u_12_14 ;
    input [11:0] vector ;
  begin
    conv_u2u_12_14 = {{2{1'b0}}, vector};
  end
  endfunction
  function automatic [13:0] conv_u2u_13_14 ;
    input [12:0] vector ;
  begin
    conv_u2u_13_14 = {1'b0, vector};
  end
  endfunction
  function automatic [15:0] conv_u2u_14_16 ;
    input [13:0] vector ;
  begin
    conv_u2u_14_16 = {{2{1'b0}}, vector};
  end
  endfunction
  function automatic [17:0] conv_u2u_14_18 ;
    input [13:0] vector ;
  begin
    conv_u2u_14_18 = {{4{1'b0}}, vector};
  end
  endfunction
  function automatic [17:0] conv_u2u_15_18 ;
    input [14:0] vector ;
  begin
    conv_u2u_15_18 = {{3{1'b0}}, vector};
  end
  endfunction
  function automatic [16:0] conv_u2u_16_17 ;
    input [15:0] vector ;
  begin
    conv_u2u_16_17 = {1'b0, vector};
  end
  endfunction
  function automatic [17:0] conv_u2u_17_18 ;
    input [16:0] vector ;
  begin
    conv_u2u_17_18 = {1'b0, vector};
  end
  endfunction
  function automatic [18:0] conv_u2u_17_19 ;
    input [16:0] vector ;
  begin
    conv_u2u_17_19 = {{2{1'b0}}, vector};
  end
  endfunction
  function automatic [31:0] conv_u2u_30_32 ;
    input [29:0] vector ;
  begin
    conv_u2u_30_32 = {{2{1'b0}}, vector};
  end
  endfunction
  function automatic [52:0] conv_u2u_52_53 ;
    input [51:0] vector ;
  begin
    conv_u2u_52_53 = {1'b0, vector};
  end
  endfunction
  function automatic [53:0] conv_u2u_53_54 ;
    input [52:0] vector ;
  begin
    conv_u2u_53_54 = {1'b0, vector};
  end
  endfunction
  function automatic [57:0] conv_u2u_57_58 ;
    input [56:0] vector ;
  begin
    conv_u2u_57_58 = {1'b0, vector};
  end
  endfunction
endmodule
module stage_struct (
  clk, rst, arst_n, ap_start_rsc_dat, ap_start_rsc_vld, ap_start_rsc_rdy, ap_done_rsc_dat,
      ap_done_rsc_vld, ap_done_rsc_rdy, mode1_rsc_dat, mode1_triosy_lz, in_f_d_rsc_adr,
      in_f_d_rsc_d, in_f_d_rsc_we, in_f_d_rsc_q, in_f_d_rsc_en, in_f_d_triosy_lz,
      in_u_rsc_adr, in_u_rsc_d, in_u_rsc_we, in_u_rsc_q, in_u_rsc_en, in_u_triosy_lz,
      out_f_d_rsc_adr, out_f_d_rsc_d, out_f_d_rsc_we, out_f_d_rsc_q, out_f_d_rsc_en,
      out_f_d_triosy_lz, out_u_rsc_adr, out_u_rsc_d, out_u_rsc_we, out_u_rsc_q, out_u_rsc_en,
      out_u_triosy_lz, out1_rsc_dat_u, out1_rsc_dat_d, out1_rsc_vld, out1_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input [15:0] mode1_rsc_dat;
  output mode1_triosy_lz;
  output [9:0] in_f_d_rsc_adr;
  output [63:0] in_f_d_rsc_d;
  output in_f_d_rsc_we;
  input [63:0] in_f_d_rsc_q;
  output in_f_d_rsc_en;
  output in_f_d_triosy_lz;
  output [9:0] in_u_rsc_adr;
  output [15:0] in_u_rsc_d;
  output in_u_rsc_we;
  input [15:0] in_u_rsc_q;
  output in_u_rsc_en;
  output in_u_triosy_lz;
  output [9:0] out_f_d_rsc_adr;
  output [63:0] out_f_d_rsc_d;
  output out_f_d_rsc_we;
  input [63:0] out_f_d_rsc_q;
  output out_f_d_rsc_en;
  output out_f_d_triosy_lz;
  output [9:0] out_u_rsc_adr;
  output [15:0] out_u_rsc_d;
  output out_u_rsc_we;
  input [15:0] out_u_rsc_q;
  output out_u_rsc_en;
  output out_u_triosy_lz;
  output [15:0] out1_rsc_dat_u;
  output [63:0] out1_rsc_dat_d;
  output out1_rsc_vld;
  input out1_rsc_rdy;
  wire [9:0] in_f_d_rsci_adr_d;
  wire [63:0] in_f_d_rsci_d_d;
  wire in_f_d_rsci_en_d;
  wire [63:0] in_f_d_rsci_q_d;
  wire in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [9:0] in_u_rsci_adr_d;
  wire [15:0] in_u_rsci_d_d;
  wire in_u_rsci_en_d;
  wire [15:0] in_u_rsci_q_d;
  wire in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [9:0] out_f_d_rsci_adr_d;
  wire [63:0] out_f_d_rsci_d_d;
  wire out_f_d_rsci_en_d;
  wire [63:0] out_f_d_rsci_q_d;
  wire out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [9:0] out_u_rsci_adr_d;
  wire [15:0] out_u_rsci_d_d;
  wire out_u_rsci_en_d;
  wire [15:0] out_u_rsci_q_d;
  wire out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [9:0] BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr;
  wire [13:0] BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out;
  wire BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en;
  wire [13:0] BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out;
  wire BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en;
  wire [13:0] BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out;
  wire BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en;
  wire [13:0] BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out;
  wire BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en;
  wire [9:0] r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_addr;
  wire [61:0] r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out;
  wire r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en;
  wire [63:0] BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out;
  wire [79:0] out1_rsc_dat;
  wire in_f_d_rsci_we_d_iff;
  wire in_u_rsci_we_d_iff;
  wire out_f_d_rsci_we_d_iff;
  wire out_u_rsci_we_d_iff;
  stagemgc_rom_sync_regout_14_1024_14_1_0_0_1_0_1_0_0_0_1_60 BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp
      (
      .addr(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .data_out(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out),
      .clk(clk),
      .s_rst(rst),
      .a_rst(arst_n),
      .en(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en)
    );
  stagemgc_rom_sync_regout_13_1024_14_1_0_0_1_0_1_0_0_0_1_60 BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp
      (
      .addr(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .data_out(BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out),
      .clk(clk),
      .s_rst(rst),
      .a_rst(arst_n),
      .en(BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en)
    );
  stagemgc_rom_sync_regout_12_1024_14_1_0_0_1_0_1_0_0_0_1_60 BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp
      (
      .addr(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .data_out(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out),
      .clk(clk),
      .s_rst(rst),
      .a_rst(arst_n),
      .en(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en)
    );
  stagemgc_rom_sync_regout_11_1024_14_1_0_0_1_0_1_0_0_0_1_60 BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp
      (
      .addr(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .data_out(BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out),
      .clk(clk),
      .s_rst(rst),
      .a_rst(arst_n),
      .en(BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en)
    );
  stagemgc_rom_sync_regout_10_1024_62_1_0_0_1_0_1_0_0_0_1_60 r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp
      (
      .addr(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_addr),
      .data_out(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out),
      .clk(clk),
      .s_rst(rst),
      .a_rst(arst_n),
      .en(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en)
    );
  stagemgc_rom_sync_regout_9_1024_64_1_0_0_1_0_1_0_0_0_1_60 BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp
      (
      .addr(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_addr),
      .data_out(BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out),
      .clk(clk),
      .s_rst(rst),
      .a_rst(arst_n),
      .en(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en)
    );
  stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_4_64_10_1024_1024_64_5_gen
      in_f_d_rsci (
      .en(in_f_d_rsc_en),
      .q(in_f_d_rsc_q),
      .we(in_f_d_rsc_we),
      .d(in_f_d_rsc_d),
      .adr(in_f_d_rsc_adr),
      .adr_d(in_f_d_rsci_adr_d),
      .d_d(in_f_d_rsci_d_d),
      .en_d(in_f_d_rsci_en_d),
      .we_d(in_f_d_rsci_we_d_iff),
      .q_d(in_f_d_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(in_f_d_rsci_we_d_iff)
    );
  stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_5_16_10_1024_1024_16_5_gen
      in_u_rsci (
      .en(in_u_rsc_en),
      .q(in_u_rsc_q),
      .we(in_u_rsc_we),
      .d(in_u_rsc_d),
      .adr(in_u_rsc_adr),
      .adr_d(in_u_rsci_adr_d),
      .d_d(in_u_rsci_d_d),
      .en_d(in_u_rsci_en_d),
      .we_d(in_u_rsci_we_d_iff),
      .q_d(in_u_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(in_u_rsci_we_d_iff)
    );
  stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_6_64_10_1024_1024_64_5_gen
      out_f_d_rsci (
      .en(out_f_d_rsc_en),
      .q(out_f_d_rsc_q),
      .we(out_f_d_rsc_we),
      .d(out_f_d_rsc_d),
      .adr(out_f_d_rsc_adr),
      .adr_d(out_f_d_rsci_adr_d),
      .d_d(out_f_d_rsci_d_d),
      .en_d(out_f_d_rsci_en_d),
      .we_d(out_f_d_rsci_we_d_iff),
      .q_d(out_f_d_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(out_f_d_rsci_we_d_iff)
    );
  stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_7_16_10_1024_1024_16_5_gen
      out_u_rsci (
      .en(out_u_rsc_en),
      .q(out_u_rsc_q),
      .we(out_u_rsc_we),
      .d(out_u_rsc_d),
      .adr(out_u_rsc_adr),
      .adr_d(out_u_rsci_adr_d),
      .d_d(out_u_rsci_d_d),
      .en_d(out_u_rsci_en_d),
      .we_d(out_u_rsci_we_d_iff),
      .q_d(out_u_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(out_u_rsci_we_d_iff)
    );
  stage_run stage_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .ap_start_rsc_dat(ap_start_rsc_dat),
      .ap_start_rsc_vld(ap_start_rsc_vld),
      .ap_start_rsc_rdy(ap_start_rsc_rdy),
      .ap_done_rsc_dat(ap_done_rsc_dat),
      .ap_done_rsc_vld(ap_done_rsc_vld),
      .ap_done_rsc_rdy(ap_done_rsc_rdy),
      .mode1_rsc_dat(mode1_rsc_dat),
      .mode1_triosy_lz(mode1_triosy_lz),
      .in_f_d_triosy_lz(in_f_d_triosy_lz),
      .in_u_triosy_lz(in_u_triosy_lz),
      .out_f_d_triosy_lz(out_f_d_triosy_lz),
      .out_u_triosy_lz(out_u_triosy_lz),
      .out1_rsc_dat(out1_rsc_dat),
      .out1_rsc_vld(out1_rsc_vld),
      .out1_rsc_rdy(out1_rsc_rdy),
      .in_f_d_rsci_adr_d(in_f_d_rsci_adr_d),
      .in_f_d_rsci_d_d(in_f_d_rsci_d_d),
      .in_f_d_rsci_en_d(in_f_d_rsci_en_d),
      .in_f_d_rsci_q_d(in_f_d_rsci_q_d),
      .in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .in_u_rsci_adr_d(in_u_rsci_adr_d),
      .in_u_rsci_d_d(in_u_rsci_d_d),
      .in_u_rsci_en_d(in_u_rsci_en_d),
      .in_u_rsci_q_d(in_u_rsci_q_d),
      .in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .out_f_d_rsci_adr_d(out_f_d_rsci_adr_d),
      .out_f_d_rsci_d_d(out_f_d_rsci_d_d),
      .out_f_d_rsci_en_d(out_f_d_rsci_en_d),
      .out_f_d_rsci_q_d(out_f_d_rsci_q_d),
      .out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .out_u_rsci_adr_d(out_u_rsci_adr_d),
      .out_u_rsci_d_d(out_u_rsci_d_d),
      .out_u_rsci_en_d(out_u_rsci_en_d),
      .out_u_rsci_q_d(out_u_rsci_q_d),
      .out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_addr),
      .BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_data_out),
      .BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en(BUTTERFLY_1_else_read_rom_GMb_rom_6_map_1_cmp_en),
      .BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out(BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_data_out),
      .BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en(BUTTERFLY_1_if_read_rom_iGMb_rom_6_map_1_cmp_en),
      .BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_data_out),
      .BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en(BUTTERFLY_else_read_rom_GMb_rom_map_1_cmp_en),
      .BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out(BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_data_out),
      .BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en(BUTTERFLY_if_read_rom_iGMb_rom_map_1_cmp_en),
      .r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_addr(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_addr),
      .r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_data_out),
      .r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en(r_ac_ieee_float_base_read_rom_gm_im_tab_d_rom_map_1_cmp_en),
      .BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out(BUTTERFLY_if_read_rom_gm_re_tab_d_rom_map_1_cmp_data_out),
      .in_f_d_rsci_we_d_pff(in_f_d_rsci_we_d_iff),
      .in_u_rsci_we_d_pff(in_u_rsci_we_d_iff),
      .out_f_d_rsci_we_d_pff(out_f_d_rsci_we_d_iff),
      .out_u_rsci_we_d_pff(out_u_rsci_we_d_iff)
    );
  assign out1_rsc_dat_d = out1_rsc_dat[63:0];
  assign out1_rsc_dat_u = out1_rsc_dat[79:64];
endmodule
module fiFFNTT (
  clk, rst, arst_n, ap_start_rsc_dat, ap_start_rsc_vld, ap_start_rsc_rdy, ap_done_rsc_dat,
      ap_done_rsc_vld, ap_done_rsc_rdy, mode1_rsc_dat, mode1_triosy_lz, in_f_d_rsc_adr,
      in_f_d_rsc_d, in_f_d_rsc_we, in_f_d_rsc_q, in_f_d_rsc_en, in_f_d_triosy_lz,
      in_u_rsc_adr, in_u_rsc_d, in_u_rsc_we, in_u_rsc_q, in_u_rsc_en, in_u_triosy_lz,
      out_f_d_rsc_adr, out_f_d_rsc_d, out_f_d_rsc_we, out_f_d_rsc_q, out_f_d_rsc_en,
      out_f_d_triosy_lz, out_u_rsc_adr, out_u_rsc_d, out_u_rsc_we, out_u_rsc_q, out_u_rsc_en,
      out_u_triosy_lz, out1_rsc_dat, out1_rsc_vld, out1_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input [15:0] mode1_rsc_dat;
  output mode1_triosy_lz;
  output [9:0] in_f_d_rsc_adr;
  output [63:0] in_f_d_rsc_d;
  output in_f_d_rsc_we;
  input [63:0] in_f_d_rsc_q;
  output in_f_d_rsc_en;
  output in_f_d_triosy_lz;
  output [9:0] in_u_rsc_adr;
  output [15:0] in_u_rsc_d;
  output in_u_rsc_we;
  input [15:0] in_u_rsc_q;
  output in_u_rsc_en;
  output in_u_triosy_lz;
  output [9:0] out_f_d_rsc_adr;
  output [63:0] out_f_d_rsc_d;
  output out_f_d_rsc_we;
  input [63:0] out_f_d_rsc_q;
  output out_f_d_rsc_en;
  output out_f_d_triosy_lz;
  output [9:0] out_u_rsc_adr;
  output [15:0] out_u_rsc_d;
  output out_u_rsc_we;
  input [15:0] out_u_rsc_q;
  output out_u_rsc_en;
  output out_u_triosy_lz;
  output [79:0] out1_rsc_dat;
  output out1_rsc_vld;
  input out1_rsc_rdy;
  wire [15:0] out1_rsc_dat_u;
  wire [63:0] out1_rsc_dat_d;
  stage_struct stage_struct_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .ap_start_rsc_dat(ap_start_rsc_dat),
      .ap_start_rsc_vld(ap_start_rsc_vld),
      .ap_start_rsc_rdy(ap_start_rsc_rdy),
      .ap_done_rsc_dat(ap_done_rsc_dat),
      .ap_done_rsc_vld(ap_done_rsc_vld),
      .ap_done_rsc_rdy(ap_done_rsc_rdy),
      .mode1_rsc_dat(mode1_rsc_dat),
      .mode1_triosy_lz(mode1_triosy_lz),
      .in_f_d_rsc_adr(in_f_d_rsc_adr),
      .in_f_d_rsc_d(in_f_d_rsc_d),
      .in_f_d_rsc_we(in_f_d_rsc_we),
      .in_f_d_rsc_q(in_f_d_rsc_q),
      .in_f_d_rsc_en(in_f_d_rsc_en),
      .in_f_d_triosy_lz(in_f_d_triosy_lz),
      .in_u_rsc_adr(in_u_rsc_adr),
      .in_u_rsc_d(in_u_rsc_d),
      .in_u_rsc_we(in_u_rsc_we),
      .in_u_rsc_q(in_u_rsc_q),
      .in_u_rsc_en(in_u_rsc_en),
      .in_u_triosy_lz(in_u_triosy_lz),
      .out_f_d_rsc_adr(out_f_d_rsc_adr),
      .out_f_d_rsc_d(out_f_d_rsc_d),
      .out_f_d_rsc_we(out_f_d_rsc_we),
      .out_f_d_rsc_q(out_f_d_rsc_q),
      .out_f_d_rsc_en(out_f_d_rsc_en),
      .out_f_d_triosy_lz(out_f_d_triosy_lz),
      .out_u_rsc_adr(out_u_rsc_adr),
      .out_u_rsc_d(out_u_rsc_d),
      .out_u_rsc_we(out_u_rsc_we),
      .out_u_rsc_q(out_u_rsc_q),
      .out_u_rsc_en(out_u_rsc_en),
      .out_u_triosy_lz(out_u_triosy_lz),
      .out1_rsc_dat_u(out1_rsc_dat_u),
      .out1_rsc_dat_d(out1_rsc_dat_d),
      .out1_rsc_vld(out1_rsc_vld),
      .out1_rsc_rdy(out1_rsc_rdy)
    );
  assign out1_rsc_dat = {out1_rsc_dat_u , out1_rsc_dat_d};
endmodule
