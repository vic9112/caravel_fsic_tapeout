
//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  localparam stallOff = 0; 
  wire                  stall_ctrl;
  assign stall_ctrl = stallOff;

  assign idat = dat;
  assign rdy = irdy && !stall_ctrl;
  assign ivld = vld && !stall_ctrl;

endmodule


//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  localparam stallOff = 0; 
  wire stall_ctrl;
  assign stall_ctrl = stallOff;

  assign dat = idat;
  assign irdy = rdy && !stall_ctrl;
  assign vld = ivld && !stall_ctrl;

endmodule



//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ../td_ccore_solutions/ROM_1i10_1o14_64308806abd59d677de1cc2043c30c27bd_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Mon May 27 10:58:41 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i10_1o14_64308806abd59d677de1cc2043c30c27bd
// ------------------------------------------------------------------


module ROM_1i10_1o14_64308806abd59d677de1cc2043c30c27bd (
  I_1, O_1
);
  input [9:0] I_1;
  output [13:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_14_1024_2(14'b00111111111011, 14'b01000100110001, 14'b00010000111001,
      14'b00010011001101, 14'b00100111100010, 14'b01011101111110, 14'b01111100001011,
      14'b01010011010001, 14'b00101000010011, 14'b01001010001111, 14'b01100101000000,
      14'b10110110110111, 14'b01101101101111, 14'b00101011111100, 14'b01011100000010,
      14'b10100111001010, 14'b00110000100101, 14'b00100001001101, 14'b00011110101000,
      14'b10101010101101, 14'b10100101101001, 14'b10100010100100, 14'b01000001011101,
      14'b00011101010011, 14'b01011011010111, 14'b10000101100010, 14'b01001000000111,
      14'b01010001000110, 14'b10110000111100, 14'b10100101010010, 14'b01011011111010,
      14'b10101110010011, 14'b10000011100001, 14'b10111111110011, 14'b10100101100111,
      14'b01110100010110, 14'b01011001010111, 14'b00110111110001, 14'b01011101011101,
      14'b10011101111100, 14'b01000101001010, 14'b10000001110010, 14'b10101000000011,
      14'b01001001000111, 14'b10101100101100, 14'b00011000000010, 14'b10111001010001,
      14'b00000001100100, 14'b10000000110111, 14'b01100111100001, 14'b10010111111101,
      14'b01010000011001, 14'b00110101010100, 14'b01111010110010, 14'b01011011000111,
      14'b10010011110100, 14'b01010001100001, 14'b10100111110100, 14'b01111011001010,
      14'b01110101010010, 14'b10111110001100, 14'b10110000011100, 14'b01011110100001,
      14'b00000001001111, 14'b00000000001101, 14'b01101100011010, 14'b10001010110110,
      14'b01010101001101, 14'b01000111101010, 14'b10110010111111, 14'b00101101010111,
      14'b01001001000100, 14'b10011001110011, 14'b01110111000101, 14'b10001001110110,
      14'b10001110010101, 14'b00100000100011, 14'b10000100111011, 14'b10000111101101,
      14'b00110000100110, 14'b01101101100111, 14'b00110011000101, 14'b00010101010111,
      14'b01100011111101, 14'b10100000010011, 14'b10000011110011, 14'b10100100011111,
      14'b10110100100111, 14'b10101101010110, 14'b00100010100011, 14'b00011100010000,
      14'b01110010010111, 14'b00000000110000, 14'b10010101001011, 14'b00101000000000,
      14'b00010011001100, 14'b10010011011110, 14'b10101000100011, 14'b10111000011000,
      14'b00011100011100, 14'b10110010001110, 14'b10001100000110, 14'b01100000001111,
      14'b00101111000100, 14'b01011111011101, 14'b00101011101100, 14'b00100010011011,
      14'b00011001110100, 14'b00001011000111, 14'b01101101011100, 14'b00010000011101,
      14'b10001100001101, 14'b01010001111100, 14'b00010111101101, 14'b10010001101010,
      14'b10110000000101, 14'b00001110000100, 14'b00111100110000, 14'b10101101111101,
      14'b10100111110000, 14'b01001101010101, 14'b01110111000000, 14'b10011011110110,
      14'b01001010001010, 14'b10100000011110, 14'b00000001111110, 14'b00101101101001,
      14'b01101001000000, 14'b01100111101011, 14'b01100110001111, 14'b00011000101110,
      14'b01001100000100, 14'b00000000101010, 14'b00001010100001, 14'b00100011000000,
      14'b01110000110011, 14'b00010100010000, 14'b10111011010101, 14'b01110111111011,
      14'b10000110000010, 14'b10111010101101, 14'b00001111011101, 14'b10100100101101,
      14'b01111000000111, 14'b01101110101101, 14'b10000100100111, 14'b00001111101100,
      14'b10011111111100, 14'b01001001011111, 14'b00000010100011, 14'b10001110110111,
      14'b01000111110101, 14'b01100100011111, 14'b10111100010100, 14'b00101110101111,
      14'b10111010100010, 14'b01001000100111, 14'b00110100100010, 14'b00100000001100,
      14'b10110001011101, 14'b10111011101011, 14'b01101000001000, 14'b01011000010111,
      14'b01110000111001, 14'b01011100011010, 14'b10010001101111, 14'b00111111111100,
      14'b01011011111000, 14'b01101100010100, 14'b00110101001010, 14'b01010000001101,
      14'b10010010110010, 14'b10101111011101, 14'b01010010000100, 14'b10001100110000,
      14'b00011000010100, 14'b01101011111100, 14'b01001010100101, 14'b00111100001101,
      14'b10001001001100, 14'b10100001010101, 14'b01111000111001, 14'b00011011011110,
      14'b01101110111111, 14'b10110001101111, 14'b10111111110001, 14'b10000110011010,
      14'b00110010101011, 14'b01100110001000, 14'b01110110100110, 14'b10000110001111,
      14'b10110100100000, 14'b01011111010101, 14'b00110010110101, 14'b10011011110001,
      14'b10010110101000, 14'b01000110011010, 14'b00111010011000, 14'b01101010101101,
      14'b10101001000110, 14'b10001110101010, 14'b10011011011100, 14'b00110111101110,
      14'b00100001010101, 14'b00111100111101, 14'b01011110010110, 14'b01110010100101,
      14'b01100111010001, 14'b00110110001100, 14'b01001000110011, 14'b00001001110001,
      14'b00101010001100, 14'b01111000111010, 14'b00110101110011, 14'b00101111110100,
      14'b00110100111100, 14'b00110111000110, 14'b01000101000010, 14'b10111010000111,
      14'b01100001011000, 14'b00011011000010, 14'b00100111111110, 14'b10100001100100,
      14'b01010011100000, 14'b01010010100110, 14'b00100010001110, 14'b10110100101010,
      14'b01100000110111, 14'b00100110110010, 14'b10001000110100, 14'b01010100001011,
      14'b01000000000101, 14'b01001000000001, 14'b10000110011101, 14'b10000000100010,
      14'b00000010010000, 14'b01011000011000, 14'b10001000000000, 14'b00101000111101,
      14'b01010100110000, 14'b10101000111100, 14'b00101110001111, 14'b10110001010010,
      14'b01100001101001, 14'b00011010110011, 14'b01001101010111, 14'b10010101000100,
      14'b00011101100000, 14'b00111010110100, 14'b00000000100111, 14'b10000000011011,
      14'b00100000100000, 14'b00100111000110, 14'b00010110111101, 14'b10100100110110,
      14'b10001000000101, 14'b01010111100001, 14'b00010001000101, 14'b00111011001000,
      14'b01001110110001, 14'b00100000001010, 14'b10000011001111, 14'b10110010111000,
      14'b10010110100111, 14'b00100000001011, 14'b10011010010110, 14'b01110011101101,
      14'b00100111000000, 14'b01111011101110, 14'b10110101001010, 14'b00000101110011,
      14'b01111100111001, 14'b00110000000001, 14'b10100001010110, 14'b00000000101000,
      14'b10011100010100, 14'b10010000011101, 14'b01111100110011, 14'b01010111100011,
      14'b00111111010011, 14'b01111011010110, 14'b00001010100100, 14'b10110001110100,
      14'b01110011010011, 14'b01100101100101, 14'b01001101110101, 14'b00101001000100,
      14'b00110110100000, 14'b10101011001100, 14'b01101101101110, 14'b01101001010001,
      14'b10011011001101, 14'b01101111100011, 14'b00100100011010, 14'b00111100101100,
      14'b01010101100001, 14'b01111010111001, 14'b01101100011101, 14'b01011001101001,
      14'b01010111101101, 14'b10010100100001, 14'b10110100110000, 14'b10110000001101,
      14'b00100111001110, 14'b01101000100001, 14'b00000110000010, 14'b01000101101110,
      14'b00000001101001, 14'b00100000011100, 14'b10100011001011, 14'b00000001110111,
      14'b00111101110011, 14'b01000100010010, 14'b10110011110001, 14'b00111001011000,
      14'b10110010101111, 14'b00001011101110, 14'b00110010101000, 14'b00110000111101,
      14'b00001011110010, 14'b00111110101101, 14'b10111010011001, 14'b10001111111010,
      14'b01010100000010, 14'b10111001101001, 14'b10101100001010, 14'b00101100000010,
      14'b00011100111011, 14'b01001101100110, 14'b01111111110101, 14'b00101010000000,
      14'b01100000111101, 14'b01101010011110, 14'b00001110011110, 14'b00101101111000,
      14'b01000011100111, 14'b10011110111111, 14'b01101110110001, 14'b01011110011111,
      14'b10010011000010, 14'b10100011111100, 14'b10001011110110, 14'b00100110101000,
      14'b01100001101111, 14'b00001011011000, 14'b01110110010001, 14'b01011110101000,
      14'b10100011000000, 14'b10101100011100, 14'b00100110010100, 14'b00101011111011,
      14'b00111011001011, 14'b00001110110001, 14'b10001100100110, 14'b00010011011100,
      14'b10001001101111, 14'b10101100001001, 14'b10101111010010, 14'b01011100000110,
      14'b01000011100101, 14'b01001000011111, 14'b00111011101011, 14'b10011001100010,
      14'b01101110010000, 14'b01101010000010, 14'b10000111011110, 14'b01010110100011,
      14'b01111000011011, 14'b00010101010001, 14'b10011001010100, 14'b00101110000101,
      14'b10110000000001, 14'b10100000111101, 14'b10001110010100, 14'b00000111011110,
      14'b01100101011001, 14'b00000001100101, 14'b00011101110111, 14'b10010100001011,
      14'b00111000011000, 14'b10111011011101, 14'b10100100101000, 14'b00001100101100,
      14'b10001011010011, 14'b00001001111101, 14'b01111111011111, 14'b01010010110011,
      14'b10001110101000, 14'b00110110111000, 14'b10000001100010, 14'b01101110011100,
      14'b01111011110010, 14'b00101111011100, 14'b01001010010111, 14'b00100001110011,
      14'b00111101100001, 14'b00111010101011, 14'b10110000101010, 14'b01111000111011,
      14'b01001100111010, 14'b10111010011100, 14'b00000110101000, 14'b01010110100010,
      14'b01100001010100, 14'b10101101111011, 14'b01111001100010, 14'b10111011000110,
      14'b00010001001001, 14'b00101101001010, 14'b10011100101011, 14'b00101000001001,
      14'b00100011001010, 14'b00100100110000, 14'b00001100110101, 14'b00100111110110,
      14'b10101100001000, 14'b01111001011001, 14'b00000010001000, 14'b00001001101001,
      14'b00110001010101, 14'b01011100000001, 14'b10010000000011, 14'b01101011000111,
      14'b00000001111000, 14'b01000100110101, 14'b00011100100001, 14'b10010110100011,
      14'b01110000101110, 14'b10100000010101, 14'b10110010000001, 14'b00100110001001,
      14'b10010101011010, 14'b10101110101000, 14'b00001001010111, 14'b00100000100101,
      14'b10110011001001, 14'b01110001000001, 14'b01100000100001, 14'b01001011000001,
      14'b10011011000110, 14'b10001100110010, 14'b01000110100010, 14'b10010011101111,
      14'b10110001011000, 14'b10110110010110, 14'b01100000011110, 14'b01111100001110,
      14'b10011000100110, 14'b01101011110000, 14'b10110101010011, 14'b00110010001101,
      14'b10000100011001, 14'b10011010010001, 14'b00101100010011, 14'b10100010110110,
      14'b00111010010100, 14'b01111100011001, 14'b00010110110001, 14'b10101001101001,
      14'b01111110000101, 14'b00001101000000, 14'b00011001011100, 14'b00110101010010,
      14'b01001100100100, 14'b10101001100111, 14'b01001111110111, 14'b10010101000111,
      14'b01100010110101, 14'b01110100000111, 14'b00111111110011, 14'b00110000000000,
      14'b10001010001111, 14'b10011001111101, 14'b10011110001010, 14'b01010010001011,
      14'b10110010010101, 14'b01100110011100, 14'b00000100101111, 14'b00010110111001,
      14'b00111100011111, 14'b01001100001001, 14'b01011010110101, 14'b10011100100001,
      14'b01101011110010, 14'b00110011101111, 14'b01011100111011, 14'b10000110111101,
      14'b01011011011100, 14'b00111100010000, 14'b00001110100000, 14'b01001101000101,
      14'b10000101010010, 14'b00011101001111, 14'b00100010001000, 14'b01010111000011,
      14'b01011011110111, 14'b00110110011001, 14'b10110101001101, 14'b10010100100111,
      14'b01111111011001, 14'b00000000100011, 14'b00101000110001, 14'b01011101001011,
      14'b01111110000000, 14'b00010000111000, 14'b10111100000111, 14'b10000011111100,
      14'b00101111101100, 14'b00111011100101, 14'b10101100111001, 14'b01101001010000,
      14'b10000100000110, 14'b00100100100100, 14'b01110111100011, 14'b00011101110110,
      14'b10100111010101, 14'b00100001000101, 14'b10010110100101, 14'b01100100000010,
      14'b01011110001100, 14'b00100001001100, 14'b01111000010101, 14'b00101001110111,
      14'b01010000111111, 14'b01100001111110, 14'b01110100000000, 14'b00101000100101,
      14'b01101010001011, 14'b10010000000110, 14'b10101001010101, 14'b00000100011000,
      14'b10000110000111, 14'b00110011000110, 14'b01101001100001, 14'b00100100110010,
      14'b00111011000011, 14'b01011111010110, 14'b01001001111100, 14'b01011100100110,
      14'b00100111000001, 14'b10000111000000, 14'b10100000110001, 14'b01011111011011,
      14'b10111101011111, 14'b00101110001110, 14'b10111111111111, 14'b10100000110100,
      14'b01111110010110, 14'b00001100110001, 14'b00111110110101, 14'b00101000110010,
      14'b00010110100100, 14'b01011100001011, 14'b10110111001000, 14'b00110011011100,
      14'b00100101111000, 14'b01001111100010, 14'b01110001001010, 14'b01010001010101,
      14'b01010010100001, 14'b10011011100100, 14'b00101010001110, 14'b01101000000000,
      14'b00001011011111, 14'b00100011000011, 14'b10110110001000, 14'b00001101000001,
      14'b00110000100011, 14'b01011101111100, 14'b01101010010001, 14'b00010001100110,
      14'b01100011000011, 14'b01010010000010, 14'b10100010010111, 14'b10010110101010,
      14'b01010010011110, 14'b00110110111001, 14'b10011000101001, 14'b00101111010001,
      14'b00001100001011, 14'b10010011011001, 14'b00110101000000, 14'b01110100001101,
      14'b00001010011100, 14'b10011111001000, 14'b01111110101111, 14'b01100101111111,
      14'b01100110101000, 14'b10101001001111, 14'b01100101010010, 14'b10000001000111,
      14'b01011001001111, 14'b10011000110100, 14'b00000111010011, 14'b01010101010110,
      14'b01000101001001, 14'b10111011011111, 14'b00010010110101, 14'b01001110010111,
      14'b01101100000110, 14'b01001111101000, 14'b00111011110011, 14'b01010110010101,
      14'b10110100111011, 14'b00110110111110, 14'b01001100001011, 14'b01110011011100,
      14'b00011110001011, 14'b01100111010111, 14'b00011000000101, 14'b10001000000100,
      14'b00000100000100, 14'b00110100111001, 14'b01001010111000, 14'b01000100100111,
      14'b01011001000001, 14'b01111011010111, 14'b00100001101011, 14'b01110010101001,
      14'b00000011101100, 14'b10100110001011, 14'b10110100001110, 14'b00011101110010,
      14'b01001010111001, 14'b10010100110111, 14'b01110001000111, 14'b10000010100010,
      14'b01010000000001, 14'b10100110100110, 14'b00100100000111, 14'b00110100010010,
      14'b10000101101100, 14'b00001011000011, 14'b00010001000000, 14'b01001101001000,
      14'b00001010100110, 14'b10100000000101, 14'b00000000010010, 14'b01011000110100,
      14'b00001111000000, 14'b01000101101011, 14'b01111100010101, 14'b00000011100010,
      14'b00100110010011, 14'b00000000000110, 14'b10001010101010, 14'b00000101000000,
      14'b01100010011010, 14'b10001100000011, 14'b10001000011111, 14'b00101100100100,
      14'b00101110100101, 14'b00011010101011, 14'b01010100100000, 14'b01001110011001,
      14'b10011010010100, 14'b10011000111110, 14'b00101110011000, 14'b00011101101011,
      14'b01101001001001, 14'b01000001010111, 14'b01010010101010, 14'b10011101100100,
      14'b01110111111111, 14'b01111100000101, 14'b10001000101000, 14'b01011000111110,
      14'b00110110000101, 14'b01000001001111, 14'b01011001110011, 14'b01010110111001,
      14'b00110100110010, 14'b01010001101011, 14'b00001110111000, 14'b01000011011111,
      14'b10011001010010, 14'b01000100000100, 14'b00110000010000, 14'b10101101101110,
      14'b00001101001000, 14'b01100001110001, 14'b00000111100110, 14'b01011101110000,
      14'b00010100111110, 14'b10100010001110, 14'b01011110000001, 14'b01001010111110,
      14'b01010101110001, 14'b01000110010010, 14'b01000001100001, 14'b00100100000010,
      14'b01100101111001, 14'b00010111000011, 14'b01100011100100, 14'b10001101000101,
      14'b01111101100101, 14'b00011001011001, 14'b01101101101100, 14'b01001010000100,
      14'b01011001100010, 14'b01111100010100, 14'b01100011001111, 14'b01100101011110,
      14'b01101100000101, 14'b10110010001101, 14'b01110100111111, 14'b10011111011010,
      14'b10011110101011, 14'b01110111110010, 14'b01110110000100, 14'b10110011110101,
      14'b00011000001010, 14'b01100110101011, 14'b10011111010111, 14'b00100011011001,
      14'b01110010011111, 14'b01011011000000, 14'b10110010000100, 14'b10110100111101,
      14'b10010111111010, 14'b00100011001011, 14'b10101110111111, 14'b01010011101100,
      14'b01110011110000, 14'b00101100101101, 14'b00111110100011, 14'b10001111111111,
      14'b00000111100100, 14'b01110101100110, 14'b10010011000001, 14'b10111111001011,
      14'b01100000001101, 14'b10001101000001, 14'b00100001001001, 14'b10100000001111,
      14'b00100111010111, 14'b10010100111101, 14'b00111011110000, 14'b10000111100010,
      14'b10110010011011, 14'b10101010001000, 14'b01001010011010, 14'b10110000100111,
      14'b01000000000001, 14'b00100101101110, 14'b01100101100000, 14'b10011011100001,
      14'b10100100111010, 14'b00001100101000, 14'b00101110110111, 14'b00100001010010,
      14'b01000010111110, 14'b10111100101110, 14'b01110100010101, 14'b01010000001100,
      14'b01111011101011, 14'b00000011110101, 14'b01011101010110, 14'b01001100001010,
      14'b01110001111100, 14'b01110110001000, 14'b10100100101011, 14'b10011011100000,
      14'b10001101110011, 14'b00100001000001, 14'b00111010001001, 14'b10100000101101,
      14'b10011100100110, 14'b10010101101010, 14'b10001011100110, 14'b10101101000010,
      14'b10010100011010, 14'b00000100100110, 14'b01001001100111, 14'b00110100111111,
      14'b00010101100001, 14'b10001101110000, 14'b10011111001101, 14'b01000111011001,
      14'b10101010001010, 14'b10011010110101, 14'b01101100001011, 14'b00000000110101,
      14'b01001000101101, 14'b00000110110111, 14'b10100000001101, 14'b01101101110100,
      14'b10011111011111, 14'b10000010010111, 14'b00010001110101, 14'b00100111111100,
      14'b01110110110001, 14'b01111111010110, 14'b10100110000110, 14'b10000111001000,
      14'b10011001101000, 14'b01111100001111, 14'b10101111101101, 14'b00100001010011,
      14'b01011010000101, 14'b10100001100111, 14'b10011000110101, 14'b00101010011110,
      14'b00010110001011, 14'b01000110110011, 14'b00111100000100, 14'b00111111100010,
      14'b01000011000101, 14'b10110110001001, 14'b10110100000101, 14'b10110001011001,
      14'b01000011011001, 14'b01001100000101, 14'b10111110011010, 14'b00011001001011,
      14'b10101010001100, 14'b10110011100001, 14'b10001010000001, 14'b00100101011001,
      14'b00000000001111, 14'b10101001001110, 14'b01001110001011, 14'b00000000010001,
      14'b00001000110101, 14'b01011100000011, 14'b10111110010001, 14'b10101100110010,
      14'b10100010101100, 14'b10001010110101, 14'b00111110000110, 14'b10101011100101,
      14'b01101111011010, 14'b01011011010000, 14'b10100011110010, 14'b10000010010010,
      14'b01011110010011, 14'b01101100110100, 14'b00011000100110, 14'b10101010111000,
      14'b00011111100100, 14'b00100110100001, 14'b01111111111111, 14'b00000110000000,
      14'b00101001010010, 14'b00101010101001, 14'b01010100010111, 14'b00100001111111,
      14'b10010010110100, 14'b10111011010011, 14'b01111101100011, 14'b01000100010111,
      14'b01100111010011, 14'b01001110010010, 14'b10111000100100, 14'b10001110101011,
      14'b10110010100011, 14'b00000001101000, 14'b01100011001100, 14'b10010110101011,
      14'b01101001100101, 14'b10111101001110, 14'b01010111110001, 14'b10101010110111,
      14'b00001000011101, 14'b00000010000111, 14'b00101111100001, 14'b01110000100000,
      14'b01100101111110, 14'b01001111011101, 14'b10111101101000, 14'b00001101001010,
      14'b01000000100001, 14'b01111000000101, 14'b10101101000111, 14'b10000011101010,
      14'b00001111110000, 14'b00101010100101, 14'b10110111111100, 14'b01011110101010,
      14'b00010001001101, 14'b00011110011110, 14'b10000011101000, 14'b01011000111000,
      14'b01101011011100, 14'b10111011100101, 14'b10011101011111, 14'b01010011010111,
      14'b00001110011111, 14'b00011011101010, 14'b00000100010001, 14'b10000010111001,
      14'b00100011011111, 14'b01010001101001, 14'b10100000101011, 14'b00000001110100,
      14'b10111000011111, 14'b00000001011011, 14'b10110110110011, 14'b00001011110101,
      14'b00010100011000, 14'b01110101100100, 14'b01100100110011, 14'b01111101100000,
      14'b01111111011010, 14'b01110100100000, 14'b01000001011111, 14'b00000100110101,
      14'b00100100001110, 14'b00100011110100, 14'b10100010011001, 14'b10110101110111,
      14'b10010100001001, 14'b10111111001110, 14'b10100101100010, 14'b10010101100001,
      14'b01111011101000, 14'b10100010000000, 14'b10011010100001, 14'b10111111010100,
      14'b01110000001011, 14'b00111101010100, 14'b00110001110100, 14'b00000101101111,
      14'b00100000011101, 14'b00000101010000, 14'b01010100001000, 14'b01010111111111,
      14'b10000110010100, 14'b01001000001101, 14'b00011011101111, 14'b10001010100010,
      14'b00000111000011, 14'b01011111011100, 14'b00010100100101, 14'b01100001100110,
      14'b10001001011011, 14'b01011100001000, 14'b01110001110011, 14'b00110000111100,
      14'b10110100101100, 14'b01001101110001, 14'b10111110000001, 14'b01110011001011,
      14'b00010101010110, 14'b10111101100010, 14'b10100101111011, 14'b00111011100001,
      14'b01010000011101, 14'b01100010011100, 14'b00101001001110, 14'b01000001100101,
      14'b00010110001010, 14'b10011101010001, 14'b01000000111100, 14'b10000010110101,
      14'b10000111000100, 14'b10100011001101, 14'b00001101110010, 14'b01111111011110,
      14'b10011110111101, 14'b10011000100011, 14'b10111110011111, 14'b00000111001011,
      14'b00101110010110, 14'b00110001011110, 14'b00000110010101, 14'b01001110001000,
      14'b10010001011111, 14'b01100100000100, 14'b10001100011010, 14'b00011000001111,
      14'b01111111101111, 14'b00111000101110, 14'b10101000001110, 14'b10010000110001,
      14'b00001010111100, 14'b10000101111101, 14'b10010100100100, 14'b01100111100110,
      14'b10110010101101, 14'b10110101001011, 14'b01011011011010, 14'b00111101101110,
      14'b01001010100111, 14'b10111010100101, 14'b00010110100110, 14'b01011110000010,
      14'b00110100111010, 14'b10110011001110, 14'b01010010111110, 14'b01010101100100,
      14'b00001000101001, 14'b10010100000010, 14'b00101000011010, 14'b00010110010111,
      14'b00101010110101, 14'b00000111011001, 14'b10110001110111, 14'b01001010001001,
      14'b00001101000100, 14'b00111111011110, 14'b10100110101010, 14'b01111000101111,
      14'b10110111101000, 14'b01010110011110, 14'b00000100111000, 14'b01000011010011,
      14'b01000011111111, 14'b01011010000100, 14'b10000111100111, 14'b10000010111101,
      14'b01111111111011, 14'b00000000000101, 14'b01110011100011, 14'b01000100001011,
      14'b00010010000000, 14'b01010100101101, 14'b01010001101111, 14'b01100101001001,
      14'b00000110110100, 14'b01110110001111, 14'b10000110011011, 14'b01100001010101,
      14'b10000000100110, I_1);

  function automatic [13:0] MUX_v_14_1024_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [13:0] input_2;
    input [13:0] input_3;
    input [13:0] input_4;
    input [13:0] input_5;
    input [13:0] input_6;
    input [13:0] input_7;
    input [13:0] input_8;
    input [13:0] input_9;
    input [13:0] input_10;
    input [13:0] input_11;
    input [13:0] input_12;
    input [13:0] input_13;
    input [13:0] input_14;
    input [13:0] input_15;
    input [13:0] input_16;
    input [13:0] input_17;
    input [13:0] input_18;
    input [13:0] input_19;
    input [13:0] input_20;
    input [13:0] input_21;
    input [13:0] input_22;
    input [13:0] input_23;
    input [13:0] input_24;
    input [13:0] input_25;
    input [13:0] input_26;
    input [13:0] input_27;
    input [13:0] input_28;
    input [13:0] input_29;
    input [13:0] input_30;
    input [13:0] input_31;
    input [13:0] input_32;
    input [13:0] input_33;
    input [13:0] input_34;
    input [13:0] input_35;
    input [13:0] input_36;
    input [13:0] input_37;
    input [13:0] input_38;
    input [13:0] input_39;
    input [13:0] input_40;
    input [13:0] input_41;
    input [13:0] input_42;
    input [13:0] input_43;
    input [13:0] input_44;
    input [13:0] input_45;
    input [13:0] input_46;
    input [13:0] input_47;
    input [13:0] input_48;
    input [13:0] input_49;
    input [13:0] input_50;
    input [13:0] input_51;
    input [13:0] input_52;
    input [13:0] input_53;
    input [13:0] input_54;
    input [13:0] input_55;
    input [13:0] input_56;
    input [13:0] input_57;
    input [13:0] input_58;
    input [13:0] input_59;
    input [13:0] input_60;
    input [13:0] input_61;
    input [13:0] input_62;
    input [13:0] input_63;
    input [13:0] input_64;
    input [13:0] input_65;
    input [13:0] input_66;
    input [13:0] input_67;
    input [13:0] input_68;
    input [13:0] input_69;
    input [13:0] input_70;
    input [13:0] input_71;
    input [13:0] input_72;
    input [13:0] input_73;
    input [13:0] input_74;
    input [13:0] input_75;
    input [13:0] input_76;
    input [13:0] input_77;
    input [13:0] input_78;
    input [13:0] input_79;
    input [13:0] input_80;
    input [13:0] input_81;
    input [13:0] input_82;
    input [13:0] input_83;
    input [13:0] input_84;
    input [13:0] input_85;
    input [13:0] input_86;
    input [13:0] input_87;
    input [13:0] input_88;
    input [13:0] input_89;
    input [13:0] input_90;
    input [13:0] input_91;
    input [13:0] input_92;
    input [13:0] input_93;
    input [13:0] input_94;
    input [13:0] input_95;
    input [13:0] input_96;
    input [13:0] input_97;
    input [13:0] input_98;
    input [13:0] input_99;
    input [13:0] input_100;
    input [13:0] input_101;
    input [13:0] input_102;
    input [13:0] input_103;
    input [13:0] input_104;
    input [13:0] input_105;
    input [13:0] input_106;
    input [13:0] input_107;
    input [13:0] input_108;
    input [13:0] input_109;
    input [13:0] input_110;
    input [13:0] input_111;
    input [13:0] input_112;
    input [13:0] input_113;
    input [13:0] input_114;
    input [13:0] input_115;
    input [13:0] input_116;
    input [13:0] input_117;
    input [13:0] input_118;
    input [13:0] input_119;
    input [13:0] input_120;
    input [13:0] input_121;
    input [13:0] input_122;
    input [13:0] input_123;
    input [13:0] input_124;
    input [13:0] input_125;
    input [13:0] input_126;
    input [13:0] input_127;
    input [13:0] input_128;
    input [13:0] input_129;
    input [13:0] input_130;
    input [13:0] input_131;
    input [13:0] input_132;
    input [13:0] input_133;
    input [13:0] input_134;
    input [13:0] input_135;
    input [13:0] input_136;
    input [13:0] input_137;
    input [13:0] input_138;
    input [13:0] input_139;
    input [13:0] input_140;
    input [13:0] input_141;
    input [13:0] input_142;
    input [13:0] input_143;
    input [13:0] input_144;
    input [13:0] input_145;
    input [13:0] input_146;
    input [13:0] input_147;
    input [13:0] input_148;
    input [13:0] input_149;
    input [13:0] input_150;
    input [13:0] input_151;
    input [13:0] input_152;
    input [13:0] input_153;
    input [13:0] input_154;
    input [13:0] input_155;
    input [13:0] input_156;
    input [13:0] input_157;
    input [13:0] input_158;
    input [13:0] input_159;
    input [13:0] input_160;
    input [13:0] input_161;
    input [13:0] input_162;
    input [13:0] input_163;
    input [13:0] input_164;
    input [13:0] input_165;
    input [13:0] input_166;
    input [13:0] input_167;
    input [13:0] input_168;
    input [13:0] input_169;
    input [13:0] input_170;
    input [13:0] input_171;
    input [13:0] input_172;
    input [13:0] input_173;
    input [13:0] input_174;
    input [13:0] input_175;
    input [13:0] input_176;
    input [13:0] input_177;
    input [13:0] input_178;
    input [13:0] input_179;
    input [13:0] input_180;
    input [13:0] input_181;
    input [13:0] input_182;
    input [13:0] input_183;
    input [13:0] input_184;
    input [13:0] input_185;
    input [13:0] input_186;
    input [13:0] input_187;
    input [13:0] input_188;
    input [13:0] input_189;
    input [13:0] input_190;
    input [13:0] input_191;
    input [13:0] input_192;
    input [13:0] input_193;
    input [13:0] input_194;
    input [13:0] input_195;
    input [13:0] input_196;
    input [13:0] input_197;
    input [13:0] input_198;
    input [13:0] input_199;
    input [13:0] input_200;
    input [13:0] input_201;
    input [13:0] input_202;
    input [13:0] input_203;
    input [13:0] input_204;
    input [13:0] input_205;
    input [13:0] input_206;
    input [13:0] input_207;
    input [13:0] input_208;
    input [13:0] input_209;
    input [13:0] input_210;
    input [13:0] input_211;
    input [13:0] input_212;
    input [13:0] input_213;
    input [13:0] input_214;
    input [13:0] input_215;
    input [13:0] input_216;
    input [13:0] input_217;
    input [13:0] input_218;
    input [13:0] input_219;
    input [13:0] input_220;
    input [13:0] input_221;
    input [13:0] input_222;
    input [13:0] input_223;
    input [13:0] input_224;
    input [13:0] input_225;
    input [13:0] input_226;
    input [13:0] input_227;
    input [13:0] input_228;
    input [13:0] input_229;
    input [13:0] input_230;
    input [13:0] input_231;
    input [13:0] input_232;
    input [13:0] input_233;
    input [13:0] input_234;
    input [13:0] input_235;
    input [13:0] input_236;
    input [13:0] input_237;
    input [13:0] input_238;
    input [13:0] input_239;
    input [13:0] input_240;
    input [13:0] input_241;
    input [13:0] input_242;
    input [13:0] input_243;
    input [13:0] input_244;
    input [13:0] input_245;
    input [13:0] input_246;
    input [13:0] input_247;
    input [13:0] input_248;
    input [13:0] input_249;
    input [13:0] input_250;
    input [13:0] input_251;
    input [13:0] input_252;
    input [13:0] input_253;
    input [13:0] input_254;
    input [13:0] input_255;
    input [13:0] input_256;
    input [13:0] input_257;
    input [13:0] input_258;
    input [13:0] input_259;
    input [13:0] input_260;
    input [13:0] input_261;
    input [13:0] input_262;
    input [13:0] input_263;
    input [13:0] input_264;
    input [13:0] input_265;
    input [13:0] input_266;
    input [13:0] input_267;
    input [13:0] input_268;
    input [13:0] input_269;
    input [13:0] input_270;
    input [13:0] input_271;
    input [13:0] input_272;
    input [13:0] input_273;
    input [13:0] input_274;
    input [13:0] input_275;
    input [13:0] input_276;
    input [13:0] input_277;
    input [13:0] input_278;
    input [13:0] input_279;
    input [13:0] input_280;
    input [13:0] input_281;
    input [13:0] input_282;
    input [13:0] input_283;
    input [13:0] input_284;
    input [13:0] input_285;
    input [13:0] input_286;
    input [13:0] input_287;
    input [13:0] input_288;
    input [13:0] input_289;
    input [13:0] input_290;
    input [13:0] input_291;
    input [13:0] input_292;
    input [13:0] input_293;
    input [13:0] input_294;
    input [13:0] input_295;
    input [13:0] input_296;
    input [13:0] input_297;
    input [13:0] input_298;
    input [13:0] input_299;
    input [13:0] input_300;
    input [13:0] input_301;
    input [13:0] input_302;
    input [13:0] input_303;
    input [13:0] input_304;
    input [13:0] input_305;
    input [13:0] input_306;
    input [13:0] input_307;
    input [13:0] input_308;
    input [13:0] input_309;
    input [13:0] input_310;
    input [13:0] input_311;
    input [13:0] input_312;
    input [13:0] input_313;
    input [13:0] input_314;
    input [13:0] input_315;
    input [13:0] input_316;
    input [13:0] input_317;
    input [13:0] input_318;
    input [13:0] input_319;
    input [13:0] input_320;
    input [13:0] input_321;
    input [13:0] input_322;
    input [13:0] input_323;
    input [13:0] input_324;
    input [13:0] input_325;
    input [13:0] input_326;
    input [13:0] input_327;
    input [13:0] input_328;
    input [13:0] input_329;
    input [13:0] input_330;
    input [13:0] input_331;
    input [13:0] input_332;
    input [13:0] input_333;
    input [13:0] input_334;
    input [13:0] input_335;
    input [13:0] input_336;
    input [13:0] input_337;
    input [13:0] input_338;
    input [13:0] input_339;
    input [13:0] input_340;
    input [13:0] input_341;
    input [13:0] input_342;
    input [13:0] input_343;
    input [13:0] input_344;
    input [13:0] input_345;
    input [13:0] input_346;
    input [13:0] input_347;
    input [13:0] input_348;
    input [13:0] input_349;
    input [13:0] input_350;
    input [13:0] input_351;
    input [13:0] input_352;
    input [13:0] input_353;
    input [13:0] input_354;
    input [13:0] input_355;
    input [13:0] input_356;
    input [13:0] input_357;
    input [13:0] input_358;
    input [13:0] input_359;
    input [13:0] input_360;
    input [13:0] input_361;
    input [13:0] input_362;
    input [13:0] input_363;
    input [13:0] input_364;
    input [13:0] input_365;
    input [13:0] input_366;
    input [13:0] input_367;
    input [13:0] input_368;
    input [13:0] input_369;
    input [13:0] input_370;
    input [13:0] input_371;
    input [13:0] input_372;
    input [13:0] input_373;
    input [13:0] input_374;
    input [13:0] input_375;
    input [13:0] input_376;
    input [13:0] input_377;
    input [13:0] input_378;
    input [13:0] input_379;
    input [13:0] input_380;
    input [13:0] input_381;
    input [13:0] input_382;
    input [13:0] input_383;
    input [13:0] input_384;
    input [13:0] input_385;
    input [13:0] input_386;
    input [13:0] input_387;
    input [13:0] input_388;
    input [13:0] input_389;
    input [13:0] input_390;
    input [13:0] input_391;
    input [13:0] input_392;
    input [13:0] input_393;
    input [13:0] input_394;
    input [13:0] input_395;
    input [13:0] input_396;
    input [13:0] input_397;
    input [13:0] input_398;
    input [13:0] input_399;
    input [13:0] input_400;
    input [13:0] input_401;
    input [13:0] input_402;
    input [13:0] input_403;
    input [13:0] input_404;
    input [13:0] input_405;
    input [13:0] input_406;
    input [13:0] input_407;
    input [13:0] input_408;
    input [13:0] input_409;
    input [13:0] input_410;
    input [13:0] input_411;
    input [13:0] input_412;
    input [13:0] input_413;
    input [13:0] input_414;
    input [13:0] input_415;
    input [13:0] input_416;
    input [13:0] input_417;
    input [13:0] input_418;
    input [13:0] input_419;
    input [13:0] input_420;
    input [13:0] input_421;
    input [13:0] input_422;
    input [13:0] input_423;
    input [13:0] input_424;
    input [13:0] input_425;
    input [13:0] input_426;
    input [13:0] input_427;
    input [13:0] input_428;
    input [13:0] input_429;
    input [13:0] input_430;
    input [13:0] input_431;
    input [13:0] input_432;
    input [13:0] input_433;
    input [13:0] input_434;
    input [13:0] input_435;
    input [13:0] input_436;
    input [13:0] input_437;
    input [13:0] input_438;
    input [13:0] input_439;
    input [13:0] input_440;
    input [13:0] input_441;
    input [13:0] input_442;
    input [13:0] input_443;
    input [13:0] input_444;
    input [13:0] input_445;
    input [13:0] input_446;
    input [13:0] input_447;
    input [13:0] input_448;
    input [13:0] input_449;
    input [13:0] input_450;
    input [13:0] input_451;
    input [13:0] input_452;
    input [13:0] input_453;
    input [13:0] input_454;
    input [13:0] input_455;
    input [13:0] input_456;
    input [13:0] input_457;
    input [13:0] input_458;
    input [13:0] input_459;
    input [13:0] input_460;
    input [13:0] input_461;
    input [13:0] input_462;
    input [13:0] input_463;
    input [13:0] input_464;
    input [13:0] input_465;
    input [13:0] input_466;
    input [13:0] input_467;
    input [13:0] input_468;
    input [13:0] input_469;
    input [13:0] input_470;
    input [13:0] input_471;
    input [13:0] input_472;
    input [13:0] input_473;
    input [13:0] input_474;
    input [13:0] input_475;
    input [13:0] input_476;
    input [13:0] input_477;
    input [13:0] input_478;
    input [13:0] input_479;
    input [13:0] input_480;
    input [13:0] input_481;
    input [13:0] input_482;
    input [13:0] input_483;
    input [13:0] input_484;
    input [13:0] input_485;
    input [13:0] input_486;
    input [13:0] input_487;
    input [13:0] input_488;
    input [13:0] input_489;
    input [13:0] input_490;
    input [13:0] input_491;
    input [13:0] input_492;
    input [13:0] input_493;
    input [13:0] input_494;
    input [13:0] input_495;
    input [13:0] input_496;
    input [13:0] input_497;
    input [13:0] input_498;
    input [13:0] input_499;
    input [13:0] input_500;
    input [13:0] input_501;
    input [13:0] input_502;
    input [13:0] input_503;
    input [13:0] input_504;
    input [13:0] input_505;
    input [13:0] input_506;
    input [13:0] input_507;
    input [13:0] input_508;
    input [13:0] input_509;
    input [13:0] input_510;
    input [13:0] input_511;
    input [13:0] input_512;
    input [13:0] input_513;
    input [13:0] input_514;
    input [13:0] input_515;
    input [13:0] input_516;
    input [13:0] input_517;
    input [13:0] input_518;
    input [13:0] input_519;
    input [13:0] input_520;
    input [13:0] input_521;
    input [13:0] input_522;
    input [13:0] input_523;
    input [13:0] input_524;
    input [13:0] input_525;
    input [13:0] input_526;
    input [13:0] input_527;
    input [13:0] input_528;
    input [13:0] input_529;
    input [13:0] input_530;
    input [13:0] input_531;
    input [13:0] input_532;
    input [13:0] input_533;
    input [13:0] input_534;
    input [13:0] input_535;
    input [13:0] input_536;
    input [13:0] input_537;
    input [13:0] input_538;
    input [13:0] input_539;
    input [13:0] input_540;
    input [13:0] input_541;
    input [13:0] input_542;
    input [13:0] input_543;
    input [13:0] input_544;
    input [13:0] input_545;
    input [13:0] input_546;
    input [13:0] input_547;
    input [13:0] input_548;
    input [13:0] input_549;
    input [13:0] input_550;
    input [13:0] input_551;
    input [13:0] input_552;
    input [13:0] input_553;
    input [13:0] input_554;
    input [13:0] input_555;
    input [13:0] input_556;
    input [13:0] input_557;
    input [13:0] input_558;
    input [13:0] input_559;
    input [13:0] input_560;
    input [13:0] input_561;
    input [13:0] input_562;
    input [13:0] input_563;
    input [13:0] input_564;
    input [13:0] input_565;
    input [13:0] input_566;
    input [13:0] input_567;
    input [13:0] input_568;
    input [13:0] input_569;
    input [13:0] input_570;
    input [13:0] input_571;
    input [13:0] input_572;
    input [13:0] input_573;
    input [13:0] input_574;
    input [13:0] input_575;
    input [13:0] input_576;
    input [13:0] input_577;
    input [13:0] input_578;
    input [13:0] input_579;
    input [13:0] input_580;
    input [13:0] input_581;
    input [13:0] input_582;
    input [13:0] input_583;
    input [13:0] input_584;
    input [13:0] input_585;
    input [13:0] input_586;
    input [13:0] input_587;
    input [13:0] input_588;
    input [13:0] input_589;
    input [13:0] input_590;
    input [13:0] input_591;
    input [13:0] input_592;
    input [13:0] input_593;
    input [13:0] input_594;
    input [13:0] input_595;
    input [13:0] input_596;
    input [13:0] input_597;
    input [13:0] input_598;
    input [13:0] input_599;
    input [13:0] input_600;
    input [13:0] input_601;
    input [13:0] input_602;
    input [13:0] input_603;
    input [13:0] input_604;
    input [13:0] input_605;
    input [13:0] input_606;
    input [13:0] input_607;
    input [13:0] input_608;
    input [13:0] input_609;
    input [13:0] input_610;
    input [13:0] input_611;
    input [13:0] input_612;
    input [13:0] input_613;
    input [13:0] input_614;
    input [13:0] input_615;
    input [13:0] input_616;
    input [13:0] input_617;
    input [13:0] input_618;
    input [13:0] input_619;
    input [13:0] input_620;
    input [13:0] input_621;
    input [13:0] input_622;
    input [13:0] input_623;
    input [13:0] input_624;
    input [13:0] input_625;
    input [13:0] input_626;
    input [13:0] input_627;
    input [13:0] input_628;
    input [13:0] input_629;
    input [13:0] input_630;
    input [13:0] input_631;
    input [13:0] input_632;
    input [13:0] input_633;
    input [13:0] input_634;
    input [13:0] input_635;
    input [13:0] input_636;
    input [13:0] input_637;
    input [13:0] input_638;
    input [13:0] input_639;
    input [13:0] input_640;
    input [13:0] input_641;
    input [13:0] input_642;
    input [13:0] input_643;
    input [13:0] input_644;
    input [13:0] input_645;
    input [13:0] input_646;
    input [13:0] input_647;
    input [13:0] input_648;
    input [13:0] input_649;
    input [13:0] input_650;
    input [13:0] input_651;
    input [13:0] input_652;
    input [13:0] input_653;
    input [13:0] input_654;
    input [13:0] input_655;
    input [13:0] input_656;
    input [13:0] input_657;
    input [13:0] input_658;
    input [13:0] input_659;
    input [13:0] input_660;
    input [13:0] input_661;
    input [13:0] input_662;
    input [13:0] input_663;
    input [13:0] input_664;
    input [13:0] input_665;
    input [13:0] input_666;
    input [13:0] input_667;
    input [13:0] input_668;
    input [13:0] input_669;
    input [13:0] input_670;
    input [13:0] input_671;
    input [13:0] input_672;
    input [13:0] input_673;
    input [13:0] input_674;
    input [13:0] input_675;
    input [13:0] input_676;
    input [13:0] input_677;
    input [13:0] input_678;
    input [13:0] input_679;
    input [13:0] input_680;
    input [13:0] input_681;
    input [13:0] input_682;
    input [13:0] input_683;
    input [13:0] input_684;
    input [13:0] input_685;
    input [13:0] input_686;
    input [13:0] input_687;
    input [13:0] input_688;
    input [13:0] input_689;
    input [13:0] input_690;
    input [13:0] input_691;
    input [13:0] input_692;
    input [13:0] input_693;
    input [13:0] input_694;
    input [13:0] input_695;
    input [13:0] input_696;
    input [13:0] input_697;
    input [13:0] input_698;
    input [13:0] input_699;
    input [13:0] input_700;
    input [13:0] input_701;
    input [13:0] input_702;
    input [13:0] input_703;
    input [13:0] input_704;
    input [13:0] input_705;
    input [13:0] input_706;
    input [13:0] input_707;
    input [13:0] input_708;
    input [13:0] input_709;
    input [13:0] input_710;
    input [13:0] input_711;
    input [13:0] input_712;
    input [13:0] input_713;
    input [13:0] input_714;
    input [13:0] input_715;
    input [13:0] input_716;
    input [13:0] input_717;
    input [13:0] input_718;
    input [13:0] input_719;
    input [13:0] input_720;
    input [13:0] input_721;
    input [13:0] input_722;
    input [13:0] input_723;
    input [13:0] input_724;
    input [13:0] input_725;
    input [13:0] input_726;
    input [13:0] input_727;
    input [13:0] input_728;
    input [13:0] input_729;
    input [13:0] input_730;
    input [13:0] input_731;
    input [13:0] input_732;
    input [13:0] input_733;
    input [13:0] input_734;
    input [13:0] input_735;
    input [13:0] input_736;
    input [13:0] input_737;
    input [13:0] input_738;
    input [13:0] input_739;
    input [13:0] input_740;
    input [13:0] input_741;
    input [13:0] input_742;
    input [13:0] input_743;
    input [13:0] input_744;
    input [13:0] input_745;
    input [13:0] input_746;
    input [13:0] input_747;
    input [13:0] input_748;
    input [13:0] input_749;
    input [13:0] input_750;
    input [13:0] input_751;
    input [13:0] input_752;
    input [13:0] input_753;
    input [13:0] input_754;
    input [13:0] input_755;
    input [13:0] input_756;
    input [13:0] input_757;
    input [13:0] input_758;
    input [13:0] input_759;
    input [13:0] input_760;
    input [13:0] input_761;
    input [13:0] input_762;
    input [13:0] input_763;
    input [13:0] input_764;
    input [13:0] input_765;
    input [13:0] input_766;
    input [13:0] input_767;
    input [13:0] input_768;
    input [13:0] input_769;
    input [13:0] input_770;
    input [13:0] input_771;
    input [13:0] input_772;
    input [13:0] input_773;
    input [13:0] input_774;
    input [13:0] input_775;
    input [13:0] input_776;
    input [13:0] input_777;
    input [13:0] input_778;
    input [13:0] input_779;
    input [13:0] input_780;
    input [13:0] input_781;
    input [13:0] input_782;
    input [13:0] input_783;
    input [13:0] input_784;
    input [13:0] input_785;
    input [13:0] input_786;
    input [13:0] input_787;
    input [13:0] input_788;
    input [13:0] input_789;
    input [13:0] input_790;
    input [13:0] input_791;
    input [13:0] input_792;
    input [13:0] input_793;
    input [13:0] input_794;
    input [13:0] input_795;
    input [13:0] input_796;
    input [13:0] input_797;
    input [13:0] input_798;
    input [13:0] input_799;
    input [13:0] input_800;
    input [13:0] input_801;
    input [13:0] input_802;
    input [13:0] input_803;
    input [13:0] input_804;
    input [13:0] input_805;
    input [13:0] input_806;
    input [13:0] input_807;
    input [13:0] input_808;
    input [13:0] input_809;
    input [13:0] input_810;
    input [13:0] input_811;
    input [13:0] input_812;
    input [13:0] input_813;
    input [13:0] input_814;
    input [13:0] input_815;
    input [13:0] input_816;
    input [13:0] input_817;
    input [13:0] input_818;
    input [13:0] input_819;
    input [13:0] input_820;
    input [13:0] input_821;
    input [13:0] input_822;
    input [13:0] input_823;
    input [13:0] input_824;
    input [13:0] input_825;
    input [13:0] input_826;
    input [13:0] input_827;
    input [13:0] input_828;
    input [13:0] input_829;
    input [13:0] input_830;
    input [13:0] input_831;
    input [13:0] input_832;
    input [13:0] input_833;
    input [13:0] input_834;
    input [13:0] input_835;
    input [13:0] input_836;
    input [13:0] input_837;
    input [13:0] input_838;
    input [13:0] input_839;
    input [13:0] input_840;
    input [13:0] input_841;
    input [13:0] input_842;
    input [13:0] input_843;
    input [13:0] input_844;
    input [13:0] input_845;
    input [13:0] input_846;
    input [13:0] input_847;
    input [13:0] input_848;
    input [13:0] input_849;
    input [13:0] input_850;
    input [13:0] input_851;
    input [13:0] input_852;
    input [13:0] input_853;
    input [13:0] input_854;
    input [13:0] input_855;
    input [13:0] input_856;
    input [13:0] input_857;
    input [13:0] input_858;
    input [13:0] input_859;
    input [13:0] input_860;
    input [13:0] input_861;
    input [13:0] input_862;
    input [13:0] input_863;
    input [13:0] input_864;
    input [13:0] input_865;
    input [13:0] input_866;
    input [13:0] input_867;
    input [13:0] input_868;
    input [13:0] input_869;
    input [13:0] input_870;
    input [13:0] input_871;
    input [13:0] input_872;
    input [13:0] input_873;
    input [13:0] input_874;
    input [13:0] input_875;
    input [13:0] input_876;
    input [13:0] input_877;
    input [13:0] input_878;
    input [13:0] input_879;
    input [13:0] input_880;
    input [13:0] input_881;
    input [13:0] input_882;
    input [13:0] input_883;
    input [13:0] input_884;
    input [13:0] input_885;
    input [13:0] input_886;
    input [13:0] input_887;
    input [13:0] input_888;
    input [13:0] input_889;
    input [13:0] input_890;
    input [13:0] input_891;
    input [13:0] input_892;
    input [13:0] input_893;
    input [13:0] input_894;
    input [13:0] input_895;
    input [13:0] input_896;
    input [13:0] input_897;
    input [13:0] input_898;
    input [13:0] input_899;
    input [13:0] input_900;
    input [13:0] input_901;
    input [13:0] input_902;
    input [13:0] input_903;
    input [13:0] input_904;
    input [13:0] input_905;
    input [13:0] input_906;
    input [13:0] input_907;
    input [13:0] input_908;
    input [13:0] input_909;
    input [13:0] input_910;
    input [13:0] input_911;
    input [13:0] input_912;
    input [13:0] input_913;
    input [13:0] input_914;
    input [13:0] input_915;
    input [13:0] input_916;
    input [13:0] input_917;
    input [13:0] input_918;
    input [13:0] input_919;
    input [13:0] input_920;
    input [13:0] input_921;
    input [13:0] input_922;
    input [13:0] input_923;
    input [13:0] input_924;
    input [13:0] input_925;
    input [13:0] input_926;
    input [13:0] input_927;
    input [13:0] input_928;
    input [13:0] input_929;
    input [13:0] input_930;
    input [13:0] input_931;
    input [13:0] input_932;
    input [13:0] input_933;
    input [13:0] input_934;
    input [13:0] input_935;
    input [13:0] input_936;
    input [13:0] input_937;
    input [13:0] input_938;
    input [13:0] input_939;
    input [13:0] input_940;
    input [13:0] input_941;
    input [13:0] input_942;
    input [13:0] input_943;
    input [13:0] input_944;
    input [13:0] input_945;
    input [13:0] input_946;
    input [13:0] input_947;
    input [13:0] input_948;
    input [13:0] input_949;
    input [13:0] input_950;
    input [13:0] input_951;
    input [13:0] input_952;
    input [13:0] input_953;
    input [13:0] input_954;
    input [13:0] input_955;
    input [13:0] input_956;
    input [13:0] input_957;
    input [13:0] input_958;
    input [13:0] input_959;
    input [13:0] input_960;
    input [13:0] input_961;
    input [13:0] input_962;
    input [13:0] input_963;
    input [13:0] input_964;
    input [13:0] input_965;
    input [13:0] input_966;
    input [13:0] input_967;
    input [13:0] input_968;
    input [13:0] input_969;
    input [13:0] input_970;
    input [13:0] input_971;
    input [13:0] input_972;
    input [13:0] input_973;
    input [13:0] input_974;
    input [13:0] input_975;
    input [13:0] input_976;
    input [13:0] input_977;
    input [13:0] input_978;
    input [13:0] input_979;
    input [13:0] input_980;
    input [13:0] input_981;
    input [13:0] input_982;
    input [13:0] input_983;
    input [13:0] input_984;
    input [13:0] input_985;
    input [13:0] input_986;
    input [13:0] input_987;
    input [13:0] input_988;
    input [13:0] input_989;
    input [13:0] input_990;
    input [13:0] input_991;
    input [13:0] input_992;
    input [13:0] input_993;
    input [13:0] input_994;
    input [13:0] input_995;
    input [13:0] input_996;
    input [13:0] input_997;
    input [13:0] input_998;
    input [13:0] input_999;
    input [13:0] input_1000;
    input [13:0] input_1001;
    input [13:0] input_1002;
    input [13:0] input_1003;
    input [13:0] input_1004;
    input [13:0] input_1005;
    input [13:0] input_1006;
    input [13:0] input_1007;
    input [13:0] input_1008;
    input [13:0] input_1009;
    input [13:0] input_1010;
    input [13:0] input_1011;
    input [13:0] input_1012;
    input [13:0] input_1013;
    input [13:0] input_1014;
    input [13:0] input_1015;
    input [13:0] input_1016;
    input [13:0] input_1017;
    input [13:0] input_1018;
    input [13:0] input_1019;
    input [13:0] input_1020;
    input [13:0] input_1021;
    input [13:0] input_1022;
    input [13:0] input_1023;
    input [9:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      10'b0000000000 : begin
        result = input_0;
      end
      10'b0000000001 : begin
        result = input_1;
      end
      10'b0000000010 : begin
        result = input_2;
      end
      10'b0000000011 : begin
        result = input_3;
      end
      10'b0000000100 : begin
        result = input_4;
      end
      10'b0000000101 : begin
        result = input_5;
      end
      10'b0000000110 : begin
        result = input_6;
      end
      10'b0000000111 : begin
        result = input_7;
      end
      10'b0000001000 : begin
        result = input_8;
      end
      10'b0000001001 : begin
        result = input_9;
      end
      10'b0000001010 : begin
        result = input_10;
      end
      10'b0000001011 : begin
        result = input_11;
      end
      10'b0000001100 : begin
        result = input_12;
      end
      10'b0000001101 : begin
        result = input_13;
      end
      10'b0000001110 : begin
        result = input_14;
      end
      10'b0000001111 : begin
        result = input_15;
      end
      10'b0000010000 : begin
        result = input_16;
      end
      10'b0000010001 : begin
        result = input_17;
      end
      10'b0000010010 : begin
        result = input_18;
      end
      10'b0000010011 : begin
        result = input_19;
      end
      10'b0000010100 : begin
        result = input_20;
      end
      10'b0000010101 : begin
        result = input_21;
      end
      10'b0000010110 : begin
        result = input_22;
      end
      10'b0000010111 : begin
        result = input_23;
      end
      10'b0000011000 : begin
        result = input_24;
      end
      10'b0000011001 : begin
        result = input_25;
      end
      10'b0000011010 : begin
        result = input_26;
      end
      10'b0000011011 : begin
        result = input_27;
      end
      10'b0000011100 : begin
        result = input_28;
      end
      10'b0000011101 : begin
        result = input_29;
      end
      10'b0000011110 : begin
        result = input_30;
      end
      10'b0000011111 : begin
        result = input_31;
      end
      10'b0000100000 : begin
        result = input_32;
      end
      10'b0000100001 : begin
        result = input_33;
      end
      10'b0000100010 : begin
        result = input_34;
      end
      10'b0000100011 : begin
        result = input_35;
      end
      10'b0000100100 : begin
        result = input_36;
      end
      10'b0000100101 : begin
        result = input_37;
      end
      10'b0000100110 : begin
        result = input_38;
      end
      10'b0000100111 : begin
        result = input_39;
      end
      10'b0000101000 : begin
        result = input_40;
      end
      10'b0000101001 : begin
        result = input_41;
      end
      10'b0000101010 : begin
        result = input_42;
      end
      10'b0000101011 : begin
        result = input_43;
      end
      10'b0000101100 : begin
        result = input_44;
      end
      10'b0000101101 : begin
        result = input_45;
      end
      10'b0000101110 : begin
        result = input_46;
      end
      10'b0000101111 : begin
        result = input_47;
      end
      10'b0000110000 : begin
        result = input_48;
      end
      10'b0000110001 : begin
        result = input_49;
      end
      10'b0000110010 : begin
        result = input_50;
      end
      10'b0000110011 : begin
        result = input_51;
      end
      10'b0000110100 : begin
        result = input_52;
      end
      10'b0000110101 : begin
        result = input_53;
      end
      10'b0000110110 : begin
        result = input_54;
      end
      10'b0000110111 : begin
        result = input_55;
      end
      10'b0000111000 : begin
        result = input_56;
      end
      10'b0000111001 : begin
        result = input_57;
      end
      10'b0000111010 : begin
        result = input_58;
      end
      10'b0000111011 : begin
        result = input_59;
      end
      10'b0000111100 : begin
        result = input_60;
      end
      10'b0000111101 : begin
        result = input_61;
      end
      10'b0000111110 : begin
        result = input_62;
      end
      10'b0000111111 : begin
        result = input_63;
      end
      10'b0001000000 : begin
        result = input_64;
      end
      10'b0001000001 : begin
        result = input_65;
      end
      10'b0001000010 : begin
        result = input_66;
      end
      10'b0001000011 : begin
        result = input_67;
      end
      10'b0001000100 : begin
        result = input_68;
      end
      10'b0001000101 : begin
        result = input_69;
      end
      10'b0001000110 : begin
        result = input_70;
      end
      10'b0001000111 : begin
        result = input_71;
      end
      10'b0001001000 : begin
        result = input_72;
      end
      10'b0001001001 : begin
        result = input_73;
      end
      10'b0001001010 : begin
        result = input_74;
      end
      10'b0001001011 : begin
        result = input_75;
      end
      10'b0001001100 : begin
        result = input_76;
      end
      10'b0001001101 : begin
        result = input_77;
      end
      10'b0001001110 : begin
        result = input_78;
      end
      10'b0001001111 : begin
        result = input_79;
      end
      10'b0001010000 : begin
        result = input_80;
      end
      10'b0001010001 : begin
        result = input_81;
      end
      10'b0001010010 : begin
        result = input_82;
      end
      10'b0001010011 : begin
        result = input_83;
      end
      10'b0001010100 : begin
        result = input_84;
      end
      10'b0001010101 : begin
        result = input_85;
      end
      10'b0001010110 : begin
        result = input_86;
      end
      10'b0001010111 : begin
        result = input_87;
      end
      10'b0001011000 : begin
        result = input_88;
      end
      10'b0001011001 : begin
        result = input_89;
      end
      10'b0001011010 : begin
        result = input_90;
      end
      10'b0001011011 : begin
        result = input_91;
      end
      10'b0001011100 : begin
        result = input_92;
      end
      10'b0001011101 : begin
        result = input_93;
      end
      10'b0001011110 : begin
        result = input_94;
      end
      10'b0001011111 : begin
        result = input_95;
      end
      10'b0001100000 : begin
        result = input_96;
      end
      10'b0001100001 : begin
        result = input_97;
      end
      10'b0001100010 : begin
        result = input_98;
      end
      10'b0001100011 : begin
        result = input_99;
      end
      10'b0001100100 : begin
        result = input_100;
      end
      10'b0001100101 : begin
        result = input_101;
      end
      10'b0001100110 : begin
        result = input_102;
      end
      10'b0001100111 : begin
        result = input_103;
      end
      10'b0001101000 : begin
        result = input_104;
      end
      10'b0001101001 : begin
        result = input_105;
      end
      10'b0001101010 : begin
        result = input_106;
      end
      10'b0001101011 : begin
        result = input_107;
      end
      10'b0001101100 : begin
        result = input_108;
      end
      10'b0001101101 : begin
        result = input_109;
      end
      10'b0001101110 : begin
        result = input_110;
      end
      10'b0001101111 : begin
        result = input_111;
      end
      10'b0001110000 : begin
        result = input_112;
      end
      10'b0001110001 : begin
        result = input_113;
      end
      10'b0001110010 : begin
        result = input_114;
      end
      10'b0001110011 : begin
        result = input_115;
      end
      10'b0001110100 : begin
        result = input_116;
      end
      10'b0001110101 : begin
        result = input_117;
      end
      10'b0001110110 : begin
        result = input_118;
      end
      10'b0001110111 : begin
        result = input_119;
      end
      10'b0001111000 : begin
        result = input_120;
      end
      10'b0001111001 : begin
        result = input_121;
      end
      10'b0001111010 : begin
        result = input_122;
      end
      10'b0001111011 : begin
        result = input_123;
      end
      10'b0001111100 : begin
        result = input_124;
      end
      10'b0001111101 : begin
        result = input_125;
      end
      10'b0001111110 : begin
        result = input_126;
      end
      10'b0001111111 : begin
        result = input_127;
      end
      10'b0010000000 : begin
        result = input_128;
      end
      10'b0010000001 : begin
        result = input_129;
      end
      10'b0010000010 : begin
        result = input_130;
      end
      10'b0010000011 : begin
        result = input_131;
      end
      10'b0010000100 : begin
        result = input_132;
      end
      10'b0010000101 : begin
        result = input_133;
      end
      10'b0010000110 : begin
        result = input_134;
      end
      10'b0010000111 : begin
        result = input_135;
      end
      10'b0010001000 : begin
        result = input_136;
      end
      10'b0010001001 : begin
        result = input_137;
      end
      10'b0010001010 : begin
        result = input_138;
      end
      10'b0010001011 : begin
        result = input_139;
      end
      10'b0010001100 : begin
        result = input_140;
      end
      10'b0010001101 : begin
        result = input_141;
      end
      10'b0010001110 : begin
        result = input_142;
      end
      10'b0010001111 : begin
        result = input_143;
      end
      10'b0010010000 : begin
        result = input_144;
      end
      10'b0010010001 : begin
        result = input_145;
      end
      10'b0010010010 : begin
        result = input_146;
      end
      10'b0010010011 : begin
        result = input_147;
      end
      10'b0010010100 : begin
        result = input_148;
      end
      10'b0010010101 : begin
        result = input_149;
      end
      10'b0010010110 : begin
        result = input_150;
      end
      10'b0010010111 : begin
        result = input_151;
      end
      10'b0010011000 : begin
        result = input_152;
      end
      10'b0010011001 : begin
        result = input_153;
      end
      10'b0010011010 : begin
        result = input_154;
      end
      10'b0010011011 : begin
        result = input_155;
      end
      10'b0010011100 : begin
        result = input_156;
      end
      10'b0010011101 : begin
        result = input_157;
      end
      10'b0010011110 : begin
        result = input_158;
      end
      10'b0010011111 : begin
        result = input_159;
      end
      10'b0010100000 : begin
        result = input_160;
      end
      10'b0010100001 : begin
        result = input_161;
      end
      10'b0010100010 : begin
        result = input_162;
      end
      10'b0010100011 : begin
        result = input_163;
      end
      10'b0010100100 : begin
        result = input_164;
      end
      10'b0010100101 : begin
        result = input_165;
      end
      10'b0010100110 : begin
        result = input_166;
      end
      10'b0010100111 : begin
        result = input_167;
      end
      10'b0010101000 : begin
        result = input_168;
      end
      10'b0010101001 : begin
        result = input_169;
      end
      10'b0010101010 : begin
        result = input_170;
      end
      10'b0010101011 : begin
        result = input_171;
      end
      10'b0010101100 : begin
        result = input_172;
      end
      10'b0010101101 : begin
        result = input_173;
      end
      10'b0010101110 : begin
        result = input_174;
      end
      10'b0010101111 : begin
        result = input_175;
      end
      10'b0010110000 : begin
        result = input_176;
      end
      10'b0010110001 : begin
        result = input_177;
      end
      10'b0010110010 : begin
        result = input_178;
      end
      10'b0010110011 : begin
        result = input_179;
      end
      10'b0010110100 : begin
        result = input_180;
      end
      10'b0010110101 : begin
        result = input_181;
      end
      10'b0010110110 : begin
        result = input_182;
      end
      10'b0010110111 : begin
        result = input_183;
      end
      10'b0010111000 : begin
        result = input_184;
      end
      10'b0010111001 : begin
        result = input_185;
      end
      10'b0010111010 : begin
        result = input_186;
      end
      10'b0010111011 : begin
        result = input_187;
      end
      10'b0010111100 : begin
        result = input_188;
      end
      10'b0010111101 : begin
        result = input_189;
      end
      10'b0010111110 : begin
        result = input_190;
      end
      10'b0010111111 : begin
        result = input_191;
      end
      10'b0011000000 : begin
        result = input_192;
      end
      10'b0011000001 : begin
        result = input_193;
      end
      10'b0011000010 : begin
        result = input_194;
      end
      10'b0011000011 : begin
        result = input_195;
      end
      10'b0011000100 : begin
        result = input_196;
      end
      10'b0011000101 : begin
        result = input_197;
      end
      10'b0011000110 : begin
        result = input_198;
      end
      10'b0011000111 : begin
        result = input_199;
      end
      10'b0011001000 : begin
        result = input_200;
      end
      10'b0011001001 : begin
        result = input_201;
      end
      10'b0011001010 : begin
        result = input_202;
      end
      10'b0011001011 : begin
        result = input_203;
      end
      10'b0011001100 : begin
        result = input_204;
      end
      10'b0011001101 : begin
        result = input_205;
      end
      10'b0011001110 : begin
        result = input_206;
      end
      10'b0011001111 : begin
        result = input_207;
      end
      10'b0011010000 : begin
        result = input_208;
      end
      10'b0011010001 : begin
        result = input_209;
      end
      10'b0011010010 : begin
        result = input_210;
      end
      10'b0011010011 : begin
        result = input_211;
      end
      10'b0011010100 : begin
        result = input_212;
      end
      10'b0011010101 : begin
        result = input_213;
      end
      10'b0011010110 : begin
        result = input_214;
      end
      10'b0011010111 : begin
        result = input_215;
      end
      10'b0011011000 : begin
        result = input_216;
      end
      10'b0011011001 : begin
        result = input_217;
      end
      10'b0011011010 : begin
        result = input_218;
      end
      10'b0011011011 : begin
        result = input_219;
      end
      10'b0011011100 : begin
        result = input_220;
      end
      10'b0011011101 : begin
        result = input_221;
      end
      10'b0011011110 : begin
        result = input_222;
      end
      10'b0011011111 : begin
        result = input_223;
      end
      10'b0011100000 : begin
        result = input_224;
      end
      10'b0011100001 : begin
        result = input_225;
      end
      10'b0011100010 : begin
        result = input_226;
      end
      10'b0011100011 : begin
        result = input_227;
      end
      10'b0011100100 : begin
        result = input_228;
      end
      10'b0011100101 : begin
        result = input_229;
      end
      10'b0011100110 : begin
        result = input_230;
      end
      10'b0011100111 : begin
        result = input_231;
      end
      10'b0011101000 : begin
        result = input_232;
      end
      10'b0011101001 : begin
        result = input_233;
      end
      10'b0011101010 : begin
        result = input_234;
      end
      10'b0011101011 : begin
        result = input_235;
      end
      10'b0011101100 : begin
        result = input_236;
      end
      10'b0011101101 : begin
        result = input_237;
      end
      10'b0011101110 : begin
        result = input_238;
      end
      10'b0011101111 : begin
        result = input_239;
      end
      10'b0011110000 : begin
        result = input_240;
      end
      10'b0011110001 : begin
        result = input_241;
      end
      10'b0011110010 : begin
        result = input_242;
      end
      10'b0011110011 : begin
        result = input_243;
      end
      10'b0011110100 : begin
        result = input_244;
      end
      10'b0011110101 : begin
        result = input_245;
      end
      10'b0011110110 : begin
        result = input_246;
      end
      10'b0011110111 : begin
        result = input_247;
      end
      10'b0011111000 : begin
        result = input_248;
      end
      10'b0011111001 : begin
        result = input_249;
      end
      10'b0011111010 : begin
        result = input_250;
      end
      10'b0011111011 : begin
        result = input_251;
      end
      10'b0011111100 : begin
        result = input_252;
      end
      10'b0011111101 : begin
        result = input_253;
      end
      10'b0011111110 : begin
        result = input_254;
      end
      10'b0011111111 : begin
        result = input_255;
      end
      10'b0100000000 : begin
        result = input_256;
      end
      10'b0100000001 : begin
        result = input_257;
      end
      10'b0100000010 : begin
        result = input_258;
      end
      10'b0100000011 : begin
        result = input_259;
      end
      10'b0100000100 : begin
        result = input_260;
      end
      10'b0100000101 : begin
        result = input_261;
      end
      10'b0100000110 : begin
        result = input_262;
      end
      10'b0100000111 : begin
        result = input_263;
      end
      10'b0100001000 : begin
        result = input_264;
      end
      10'b0100001001 : begin
        result = input_265;
      end
      10'b0100001010 : begin
        result = input_266;
      end
      10'b0100001011 : begin
        result = input_267;
      end
      10'b0100001100 : begin
        result = input_268;
      end
      10'b0100001101 : begin
        result = input_269;
      end
      10'b0100001110 : begin
        result = input_270;
      end
      10'b0100001111 : begin
        result = input_271;
      end
      10'b0100010000 : begin
        result = input_272;
      end
      10'b0100010001 : begin
        result = input_273;
      end
      10'b0100010010 : begin
        result = input_274;
      end
      10'b0100010011 : begin
        result = input_275;
      end
      10'b0100010100 : begin
        result = input_276;
      end
      10'b0100010101 : begin
        result = input_277;
      end
      10'b0100010110 : begin
        result = input_278;
      end
      10'b0100010111 : begin
        result = input_279;
      end
      10'b0100011000 : begin
        result = input_280;
      end
      10'b0100011001 : begin
        result = input_281;
      end
      10'b0100011010 : begin
        result = input_282;
      end
      10'b0100011011 : begin
        result = input_283;
      end
      10'b0100011100 : begin
        result = input_284;
      end
      10'b0100011101 : begin
        result = input_285;
      end
      10'b0100011110 : begin
        result = input_286;
      end
      10'b0100011111 : begin
        result = input_287;
      end
      10'b0100100000 : begin
        result = input_288;
      end
      10'b0100100001 : begin
        result = input_289;
      end
      10'b0100100010 : begin
        result = input_290;
      end
      10'b0100100011 : begin
        result = input_291;
      end
      10'b0100100100 : begin
        result = input_292;
      end
      10'b0100100101 : begin
        result = input_293;
      end
      10'b0100100110 : begin
        result = input_294;
      end
      10'b0100100111 : begin
        result = input_295;
      end
      10'b0100101000 : begin
        result = input_296;
      end
      10'b0100101001 : begin
        result = input_297;
      end
      10'b0100101010 : begin
        result = input_298;
      end
      10'b0100101011 : begin
        result = input_299;
      end
      10'b0100101100 : begin
        result = input_300;
      end
      10'b0100101101 : begin
        result = input_301;
      end
      10'b0100101110 : begin
        result = input_302;
      end
      10'b0100101111 : begin
        result = input_303;
      end
      10'b0100110000 : begin
        result = input_304;
      end
      10'b0100110001 : begin
        result = input_305;
      end
      10'b0100110010 : begin
        result = input_306;
      end
      10'b0100110011 : begin
        result = input_307;
      end
      10'b0100110100 : begin
        result = input_308;
      end
      10'b0100110101 : begin
        result = input_309;
      end
      10'b0100110110 : begin
        result = input_310;
      end
      10'b0100110111 : begin
        result = input_311;
      end
      10'b0100111000 : begin
        result = input_312;
      end
      10'b0100111001 : begin
        result = input_313;
      end
      10'b0100111010 : begin
        result = input_314;
      end
      10'b0100111011 : begin
        result = input_315;
      end
      10'b0100111100 : begin
        result = input_316;
      end
      10'b0100111101 : begin
        result = input_317;
      end
      10'b0100111110 : begin
        result = input_318;
      end
      10'b0100111111 : begin
        result = input_319;
      end
      10'b0101000000 : begin
        result = input_320;
      end
      10'b0101000001 : begin
        result = input_321;
      end
      10'b0101000010 : begin
        result = input_322;
      end
      10'b0101000011 : begin
        result = input_323;
      end
      10'b0101000100 : begin
        result = input_324;
      end
      10'b0101000101 : begin
        result = input_325;
      end
      10'b0101000110 : begin
        result = input_326;
      end
      10'b0101000111 : begin
        result = input_327;
      end
      10'b0101001000 : begin
        result = input_328;
      end
      10'b0101001001 : begin
        result = input_329;
      end
      10'b0101001010 : begin
        result = input_330;
      end
      10'b0101001011 : begin
        result = input_331;
      end
      10'b0101001100 : begin
        result = input_332;
      end
      10'b0101001101 : begin
        result = input_333;
      end
      10'b0101001110 : begin
        result = input_334;
      end
      10'b0101001111 : begin
        result = input_335;
      end
      10'b0101010000 : begin
        result = input_336;
      end
      10'b0101010001 : begin
        result = input_337;
      end
      10'b0101010010 : begin
        result = input_338;
      end
      10'b0101010011 : begin
        result = input_339;
      end
      10'b0101010100 : begin
        result = input_340;
      end
      10'b0101010101 : begin
        result = input_341;
      end
      10'b0101010110 : begin
        result = input_342;
      end
      10'b0101010111 : begin
        result = input_343;
      end
      10'b0101011000 : begin
        result = input_344;
      end
      10'b0101011001 : begin
        result = input_345;
      end
      10'b0101011010 : begin
        result = input_346;
      end
      10'b0101011011 : begin
        result = input_347;
      end
      10'b0101011100 : begin
        result = input_348;
      end
      10'b0101011101 : begin
        result = input_349;
      end
      10'b0101011110 : begin
        result = input_350;
      end
      10'b0101011111 : begin
        result = input_351;
      end
      10'b0101100000 : begin
        result = input_352;
      end
      10'b0101100001 : begin
        result = input_353;
      end
      10'b0101100010 : begin
        result = input_354;
      end
      10'b0101100011 : begin
        result = input_355;
      end
      10'b0101100100 : begin
        result = input_356;
      end
      10'b0101100101 : begin
        result = input_357;
      end
      10'b0101100110 : begin
        result = input_358;
      end
      10'b0101100111 : begin
        result = input_359;
      end
      10'b0101101000 : begin
        result = input_360;
      end
      10'b0101101001 : begin
        result = input_361;
      end
      10'b0101101010 : begin
        result = input_362;
      end
      10'b0101101011 : begin
        result = input_363;
      end
      10'b0101101100 : begin
        result = input_364;
      end
      10'b0101101101 : begin
        result = input_365;
      end
      10'b0101101110 : begin
        result = input_366;
      end
      10'b0101101111 : begin
        result = input_367;
      end
      10'b0101110000 : begin
        result = input_368;
      end
      10'b0101110001 : begin
        result = input_369;
      end
      10'b0101110010 : begin
        result = input_370;
      end
      10'b0101110011 : begin
        result = input_371;
      end
      10'b0101110100 : begin
        result = input_372;
      end
      10'b0101110101 : begin
        result = input_373;
      end
      10'b0101110110 : begin
        result = input_374;
      end
      10'b0101110111 : begin
        result = input_375;
      end
      10'b0101111000 : begin
        result = input_376;
      end
      10'b0101111001 : begin
        result = input_377;
      end
      10'b0101111010 : begin
        result = input_378;
      end
      10'b0101111011 : begin
        result = input_379;
      end
      10'b0101111100 : begin
        result = input_380;
      end
      10'b0101111101 : begin
        result = input_381;
      end
      10'b0101111110 : begin
        result = input_382;
      end
      10'b0101111111 : begin
        result = input_383;
      end
      10'b0110000000 : begin
        result = input_384;
      end
      10'b0110000001 : begin
        result = input_385;
      end
      10'b0110000010 : begin
        result = input_386;
      end
      10'b0110000011 : begin
        result = input_387;
      end
      10'b0110000100 : begin
        result = input_388;
      end
      10'b0110000101 : begin
        result = input_389;
      end
      10'b0110000110 : begin
        result = input_390;
      end
      10'b0110000111 : begin
        result = input_391;
      end
      10'b0110001000 : begin
        result = input_392;
      end
      10'b0110001001 : begin
        result = input_393;
      end
      10'b0110001010 : begin
        result = input_394;
      end
      10'b0110001011 : begin
        result = input_395;
      end
      10'b0110001100 : begin
        result = input_396;
      end
      10'b0110001101 : begin
        result = input_397;
      end
      10'b0110001110 : begin
        result = input_398;
      end
      10'b0110001111 : begin
        result = input_399;
      end
      10'b0110010000 : begin
        result = input_400;
      end
      10'b0110010001 : begin
        result = input_401;
      end
      10'b0110010010 : begin
        result = input_402;
      end
      10'b0110010011 : begin
        result = input_403;
      end
      10'b0110010100 : begin
        result = input_404;
      end
      10'b0110010101 : begin
        result = input_405;
      end
      10'b0110010110 : begin
        result = input_406;
      end
      10'b0110010111 : begin
        result = input_407;
      end
      10'b0110011000 : begin
        result = input_408;
      end
      10'b0110011001 : begin
        result = input_409;
      end
      10'b0110011010 : begin
        result = input_410;
      end
      10'b0110011011 : begin
        result = input_411;
      end
      10'b0110011100 : begin
        result = input_412;
      end
      10'b0110011101 : begin
        result = input_413;
      end
      10'b0110011110 : begin
        result = input_414;
      end
      10'b0110011111 : begin
        result = input_415;
      end
      10'b0110100000 : begin
        result = input_416;
      end
      10'b0110100001 : begin
        result = input_417;
      end
      10'b0110100010 : begin
        result = input_418;
      end
      10'b0110100011 : begin
        result = input_419;
      end
      10'b0110100100 : begin
        result = input_420;
      end
      10'b0110100101 : begin
        result = input_421;
      end
      10'b0110100110 : begin
        result = input_422;
      end
      10'b0110100111 : begin
        result = input_423;
      end
      10'b0110101000 : begin
        result = input_424;
      end
      10'b0110101001 : begin
        result = input_425;
      end
      10'b0110101010 : begin
        result = input_426;
      end
      10'b0110101011 : begin
        result = input_427;
      end
      10'b0110101100 : begin
        result = input_428;
      end
      10'b0110101101 : begin
        result = input_429;
      end
      10'b0110101110 : begin
        result = input_430;
      end
      10'b0110101111 : begin
        result = input_431;
      end
      10'b0110110000 : begin
        result = input_432;
      end
      10'b0110110001 : begin
        result = input_433;
      end
      10'b0110110010 : begin
        result = input_434;
      end
      10'b0110110011 : begin
        result = input_435;
      end
      10'b0110110100 : begin
        result = input_436;
      end
      10'b0110110101 : begin
        result = input_437;
      end
      10'b0110110110 : begin
        result = input_438;
      end
      10'b0110110111 : begin
        result = input_439;
      end
      10'b0110111000 : begin
        result = input_440;
      end
      10'b0110111001 : begin
        result = input_441;
      end
      10'b0110111010 : begin
        result = input_442;
      end
      10'b0110111011 : begin
        result = input_443;
      end
      10'b0110111100 : begin
        result = input_444;
      end
      10'b0110111101 : begin
        result = input_445;
      end
      10'b0110111110 : begin
        result = input_446;
      end
      10'b0110111111 : begin
        result = input_447;
      end
      10'b0111000000 : begin
        result = input_448;
      end
      10'b0111000001 : begin
        result = input_449;
      end
      10'b0111000010 : begin
        result = input_450;
      end
      10'b0111000011 : begin
        result = input_451;
      end
      10'b0111000100 : begin
        result = input_452;
      end
      10'b0111000101 : begin
        result = input_453;
      end
      10'b0111000110 : begin
        result = input_454;
      end
      10'b0111000111 : begin
        result = input_455;
      end
      10'b0111001000 : begin
        result = input_456;
      end
      10'b0111001001 : begin
        result = input_457;
      end
      10'b0111001010 : begin
        result = input_458;
      end
      10'b0111001011 : begin
        result = input_459;
      end
      10'b0111001100 : begin
        result = input_460;
      end
      10'b0111001101 : begin
        result = input_461;
      end
      10'b0111001110 : begin
        result = input_462;
      end
      10'b0111001111 : begin
        result = input_463;
      end
      10'b0111010000 : begin
        result = input_464;
      end
      10'b0111010001 : begin
        result = input_465;
      end
      10'b0111010010 : begin
        result = input_466;
      end
      10'b0111010011 : begin
        result = input_467;
      end
      10'b0111010100 : begin
        result = input_468;
      end
      10'b0111010101 : begin
        result = input_469;
      end
      10'b0111010110 : begin
        result = input_470;
      end
      10'b0111010111 : begin
        result = input_471;
      end
      10'b0111011000 : begin
        result = input_472;
      end
      10'b0111011001 : begin
        result = input_473;
      end
      10'b0111011010 : begin
        result = input_474;
      end
      10'b0111011011 : begin
        result = input_475;
      end
      10'b0111011100 : begin
        result = input_476;
      end
      10'b0111011101 : begin
        result = input_477;
      end
      10'b0111011110 : begin
        result = input_478;
      end
      10'b0111011111 : begin
        result = input_479;
      end
      10'b0111100000 : begin
        result = input_480;
      end
      10'b0111100001 : begin
        result = input_481;
      end
      10'b0111100010 : begin
        result = input_482;
      end
      10'b0111100011 : begin
        result = input_483;
      end
      10'b0111100100 : begin
        result = input_484;
      end
      10'b0111100101 : begin
        result = input_485;
      end
      10'b0111100110 : begin
        result = input_486;
      end
      10'b0111100111 : begin
        result = input_487;
      end
      10'b0111101000 : begin
        result = input_488;
      end
      10'b0111101001 : begin
        result = input_489;
      end
      10'b0111101010 : begin
        result = input_490;
      end
      10'b0111101011 : begin
        result = input_491;
      end
      10'b0111101100 : begin
        result = input_492;
      end
      10'b0111101101 : begin
        result = input_493;
      end
      10'b0111101110 : begin
        result = input_494;
      end
      10'b0111101111 : begin
        result = input_495;
      end
      10'b0111110000 : begin
        result = input_496;
      end
      10'b0111110001 : begin
        result = input_497;
      end
      10'b0111110010 : begin
        result = input_498;
      end
      10'b0111110011 : begin
        result = input_499;
      end
      10'b0111110100 : begin
        result = input_500;
      end
      10'b0111110101 : begin
        result = input_501;
      end
      10'b0111110110 : begin
        result = input_502;
      end
      10'b0111110111 : begin
        result = input_503;
      end
      10'b0111111000 : begin
        result = input_504;
      end
      10'b0111111001 : begin
        result = input_505;
      end
      10'b0111111010 : begin
        result = input_506;
      end
      10'b0111111011 : begin
        result = input_507;
      end
      10'b0111111100 : begin
        result = input_508;
      end
      10'b0111111101 : begin
        result = input_509;
      end
      10'b0111111110 : begin
        result = input_510;
      end
      10'b0111111111 : begin
        result = input_511;
      end
      10'b1000000000 : begin
        result = input_512;
      end
      10'b1000000001 : begin
        result = input_513;
      end
      10'b1000000010 : begin
        result = input_514;
      end
      10'b1000000011 : begin
        result = input_515;
      end
      10'b1000000100 : begin
        result = input_516;
      end
      10'b1000000101 : begin
        result = input_517;
      end
      10'b1000000110 : begin
        result = input_518;
      end
      10'b1000000111 : begin
        result = input_519;
      end
      10'b1000001000 : begin
        result = input_520;
      end
      10'b1000001001 : begin
        result = input_521;
      end
      10'b1000001010 : begin
        result = input_522;
      end
      10'b1000001011 : begin
        result = input_523;
      end
      10'b1000001100 : begin
        result = input_524;
      end
      10'b1000001101 : begin
        result = input_525;
      end
      10'b1000001110 : begin
        result = input_526;
      end
      10'b1000001111 : begin
        result = input_527;
      end
      10'b1000010000 : begin
        result = input_528;
      end
      10'b1000010001 : begin
        result = input_529;
      end
      10'b1000010010 : begin
        result = input_530;
      end
      10'b1000010011 : begin
        result = input_531;
      end
      10'b1000010100 : begin
        result = input_532;
      end
      10'b1000010101 : begin
        result = input_533;
      end
      10'b1000010110 : begin
        result = input_534;
      end
      10'b1000010111 : begin
        result = input_535;
      end
      10'b1000011000 : begin
        result = input_536;
      end
      10'b1000011001 : begin
        result = input_537;
      end
      10'b1000011010 : begin
        result = input_538;
      end
      10'b1000011011 : begin
        result = input_539;
      end
      10'b1000011100 : begin
        result = input_540;
      end
      10'b1000011101 : begin
        result = input_541;
      end
      10'b1000011110 : begin
        result = input_542;
      end
      10'b1000011111 : begin
        result = input_543;
      end
      10'b1000100000 : begin
        result = input_544;
      end
      10'b1000100001 : begin
        result = input_545;
      end
      10'b1000100010 : begin
        result = input_546;
      end
      10'b1000100011 : begin
        result = input_547;
      end
      10'b1000100100 : begin
        result = input_548;
      end
      10'b1000100101 : begin
        result = input_549;
      end
      10'b1000100110 : begin
        result = input_550;
      end
      10'b1000100111 : begin
        result = input_551;
      end
      10'b1000101000 : begin
        result = input_552;
      end
      10'b1000101001 : begin
        result = input_553;
      end
      10'b1000101010 : begin
        result = input_554;
      end
      10'b1000101011 : begin
        result = input_555;
      end
      10'b1000101100 : begin
        result = input_556;
      end
      10'b1000101101 : begin
        result = input_557;
      end
      10'b1000101110 : begin
        result = input_558;
      end
      10'b1000101111 : begin
        result = input_559;
      end
      10'b1000110000 : begin
        result = input_560;
      end
      10'b1000110001 : begin
        result = input_561;
      end
      10'b1000110010 : begin
        result = input_562;
      end
      10'b1000110011 : begin
        result = input_563;
      end
      10'b1000110100 : begin
        result = input_564;
      end
      10'b1000110101 : begin
        result = input_565;
      end
      10'b1000110110 : begin
        result = input_566;
      end
      10'b1000110111 : begin
        result = input_567;
      end
      10'b1000111000 : begin
        result = input_568;
      end
      10'b1000111001 : begin
        result = input_569;
      end
      10'b1000111010 : begin
        result = input_570;
      end
      10'b1000111011 : begin
        result = input_571;
      end
      10'b1000111100 : begin
        result = input_572;
      end
      10'b1000111101 : begin
        result = input_573;
      end
      10'b1000111110 : begin
        result = input_574;
      end
      10'b1000111111 : begin
        result = input_575;
      end
      10'b1001000000 : begin
        result = input_576;
      end
      10'b1001000001 : begin
        result = input_577;
      end
      10'b1001000010 : begin
        result = input_578;
      end
      10'b1001000011 : begin
        result = input_579;
      end
      10'b1001000100 : begin
        result = input_580;
      end
      10'b1001000101 : begin
        result = input_581;
      end
      10'b1001000110 : begin
        result = input_582;
      end
      10'b1001000111 : begin
        result = input_583;
      end
      10'b1001001000 : begin
        result = input_584;
      end
      10'b1001001001 : begin
        result = input_585;
      end
      10'b1001001010 : begin
        result = input_586;
      end
      10'b1001001011 : begin
        result = input_587;
      end
      10'b1001001100 : begin
        result = input_588;
      end
      10'b1001001101 : begin
        result = input_589;
      end
      10'b1001001110 : begin
        result = input_590;
      end
      10'b1001001111 : begin
        result = input_591;
      end
      10'b1001010000 : begin
        result = input_592;
      end
      10'b1001010001 : begin
        result = input_593;
      end
      10'b1001010010 : begin
        result = input_594;
      end
      10'b1001010011 : begin
        result = input_595;
      end
      10'b1001010100 : begin
        result = input_596;
      end
      10'b1001010101 : begin
        result = input_597;
      end
      10'b1001010110 : begin
        result = input_598;
      end
      10'b1001010111 : begin
        result = input_599;
      end
      10'b1001011000 : begin
        result = input_600;
      end
      10'b1001011001 : begin
        result = input_601;
      end
      10'b1001011010 : begin
        result = input_602;
      end
      10'b1001011011 : begin
        result = input_603;
      end
      10'b1001011100 : begin
        result = input_604;
      end
      10'b1001011101 : begin
        result = input_605;
      end
      10'b1001011110 : begin
        result = input_606;
      end
      10'b1001011111 : begin
        result = input_607;
      end
      10'b1001100000 : begin
        result = input_608;
      end
      10'b1001100001 : begin
        result = input_609;
      end
      10'b1001100010 : begin
        result = input_610;
      end
      10'b1001100011 : begin
        result = input_611;
      end
      10'b1001100100 : begin
        result = input_612;
      end
      10'b1001100101 : begin
        result = input_613;
      end
      10'b1001100110 : begin
        result = input_614;
      end
      10'b1001100111 : begin
        result = input_615;
      end
      10'b1001101000 : begin
        result = input_616;
      end
      10'b1001101001 : begin
        result = input_617;
      end
      10'b1001101010 : begin
        result = input_618;
      end
      10'b1001101011 : begin
        result = input_619;
      end
      10'b1001101100 : begin
        result = input_620;
      end
      10'b1001101101 : begin
        result = input_621;
      end
      10'b1001101110 : begin
        result = input_622;
      end
      10'b1001101111 : begin
        result = input_623;
      end
      10'b1001110000 : begin
        result = input_624;
      end
      10'b1001110001 : begin
        result = input_625;
      end
      10'b1001110010 : begin
        result = input_626;
      end
      10'b1001110011 : begin
        result = input_627;
      end
      10'b1001110100 : begin
        result = input_628;
      end
      10'b1001110101 : begin
        result = input_629;
      end
      10'b1001110110 : begin
        result = input_630;
      end
      10'b1001110111 : begin
        result = input_631;
      end
      10'b1001111000 : begin
        result = input_632;
      end
      10'b1001111001 : begin
        result = input_633;
      end
      10'b1001111010 : begin
        result = input_634;
      end
      10'b1001111011 : begin
        result = input_635;
      end
      10'b1001111100 : begin
        result = input_636;
      end
      10'b1001111101 : begin
        result = input_637;
      end
      10'b1001111110 : begin
        result = input_638;
      end
      10'b1001111111 : begin
        result = input_639;
      end
      10'b1010000000 : begin
        result = input_640;
      end
      10'b1010000001 : begin
        result = input_641;
      end
      10'b1010000010 : begin
        result = input_642;
      end
      10'b1010000011 : begin
        result = input_643;
      end
      10'b1010000100 : begin
        result = input_644;
      end
      10'b1010000101 : begin
        result = input_645;
      end
      10'b1010000110 : begin
        result = input_646;
      end
      10'b1010000111 : begin
        result = input_647;
      end
      10'b1010001000 : begin
        result = input_648;
      end
      10'b1010001001 : begin
        result = input_649;
      end
      10'b1010001010 : begin
        result = input_650;
      end
      10'b1010001011 : begin
        result = input_651;
      end
      10'b1010001100 : begin
        result = input_652;
      end
      10'b1010001101 : begin
        result = input_653;
      end
      10'b1010001110 : begin
        result = input_654;
      end
      10'b1010001111 : begin
        result = input_655;
      end
      10'b1010010000 : begin
        result = input_656;
      end
      10'b1010010001 : begin
        result = input_657;
      end
      10'b1010010010 : begin
        result = input_658;
      end
      10'b1010010011 : begin
        result = input_659;
      end
      10'b1010010100 : begin
        result = input_660;
      end
      10'b1010010101 : begin
        result = input_661;
      end
      10'b1010010110 : begin
        result = input_662;
      end
      10'b1010010111 : begin
        result = input_663;
      end
      10'b1010011000 : begin
        result = input_664;
      end
      10'b1010011001 : begin
        result = input_665;
      end
      10'b1010011010 : begin
        result = input_666;
      end
      10'b1010011011 : begin
        result = input_667;
      end
      10'b1010011100 : begin
        result = input_668;
      end
      10'b1010011101 : begin
        result = input_669;
      end
      10'b1010011110 : begin
        result = input_670;
      end
      10'b1010011111 : begin
        result = input_671;
      end
      10'b1010100000 : begin
        result = input_672;
      end
      10'b1010100001 : begin
        result = input_673;
      end
      10'b1010100010 : begin
        result = input_674;
      end
      10'b1010100011 : begin
        result = input_675;
      end
      10'b1010100100 : begin
        result = input_676;
      end
      10'b1010100101 : begin
        result = input_677;
      end
      10'b1010100110 : begin
        result = input_678;
      end
      10'b1010100111 : begin
        result = input_679;
      end
      10'b1010101000 : begin
        result = input_680;
      end
      10'b1010101001 : begin
        result = input_681;
      end
      10'b1010101010 : begin
        result = input_682;
      end
      10'b1010101011 : begin
        result = input_683;
      end
      10'b1010101100 : begin
        result = input_684;
      end
      10'b1010101101 : begin
        result = input_685;
      end
      10'b1010101110 : begin
        result = input_686;
      end
      10'b1010101111 : begin
        result = input_687;
      end
      10'b1010110000 : begin
        result = input_688;
      end
      10'b1010110001 : begin
        result = input_689;
      end
      10'b1010110010 : begin
        result = input_690;
      end
      10'b1010110011 : begin
        result = input_691;
      end
      10'b1010110100 : begin
        result = input_692;
      end
      10'b1010110101 : begin
        result = input_693;
      end
      10'b1010110110 : begin
        result = input_694;
      end
      10'b1010110111 : begin
        result = input_695;
      end
      10'b1010111000 : begin
        result = input_696;
      end
      10'b1010111001 : begin
        result = input_697;
      end
      10'b1010111010 : begin
        result = input_698;
      end
      10'b1010111011 : begin
        result = input_699;
      end
      10'b1010111100 : begin
        result = input_700;
      end
      10'b1010111101 : begin
        result = input_701;
      end
      10'b1010111110 : begin
        result = input_702;
      end
      10'b1010111111 : begin
        result = input_703;
      end
      10'b1011000000 : begin
        result = input_704;
      end
      10'b1011000001 : begin
        result = input_705;
      end
      10'b1011000010 : begin
        result = input_706;
      end
      10'b1011000011 : begin
        result = input_707;
      end
      10'b1011000100 : begin
        result = input_708;
      end
      10'b1011000101 : begin
        result = input_709;
      end
      10'b1011000110 : begin
        result = input_710;
      end
      10'b1011000111 : begin
        result = input_711;
      end
      10'b1011001000 : begin
        result = input_712;
      end
      10'b1011001001 : begin
        result = input_713;
      end
      10'b1011001010 : begin
        result = input_714;
      end
      10'b1011001011 : begin
        result = input_715;
      end
      10'b1011001100 : begin
        result = input_716;
      end
      10'b1011001101 : begin
        result = input_717;
      end
      10'b1011001110 : begin
        result = input_718;
      end
      10'b1011001111 : begin
        result = input_719;
      end
      10'b1011010000 : begin
        result = input_720;
      end
      10'b1011010001 : begin
        result = input_721;
      end
      10'b1011010010 : begin
        result = input_722;
      end
      10'b1011010011 : begin
        result = input_723;
      end
      10'b1011010100 : begin
        result = input_724;
      end
      10'b1011010101 : begin
        result = input_725;
      end
      10'b1011010110 : begin
        result = input_726;
      end
      10'b1011010111 : begin
        result = input_727;
      end
      10'b1011011000 : begin
        result = input_728;
      end
      10'b1011011001 : begin
        result = input_729;
      end
      10'b1011011010 : begin
        result = input_730;
      end
      10'b1011011011 : begin
        result = input_731;
      end
      10'b1011011100 : begin
        result = input_732;
      end
      10'b1011011101 : begin
        result = input_733;
      end
      10'b1011011110 : begin
        result = input_734;
      end
      10'b1011011111 : begin
        result = input_735;
      end
      10'b1011100000 : begin
        result = input_736;
      end
      10'b1011100001 : begin
        result = input_737;
      end
      10'b1011100010 : begin
        result = input_738;
      end
      10'b1011100011 : begin
        result = input_739;
      end
      10'b1011100100 : begin
        result = input_740;
      end
      10'b1011100101 : begin
        result = input_741;
      end
      10'b1011100110 : begin
        result = input_742;
      end
      10'b1011100111 : begin
        result = input_743;
      end
      10'b1011101000 : begin
        result = input_744;
      end
      10'b1011101001 : begin
        result = input_745;
      end
      10'b1011101010 : begin
        result = input_746;
      end
      10'b1011101011 : begin
        result = input_747;
      end
      10'b1011101100 : begin
        result = input_748;
      end
      10'b1011101101 : begin
        result = input_749;
      end
      10'b1011101110 : begin
        result = input_750;
      end
      10'b1011101111 : begin
        result = input_751;
      end
      10'b1011110000 : begin
        result = input_752;
      end
      10'b1011110001 : begin
        result = input_753;
      end
      10'b1011110010 : begin
        result = input_754;
      end
      10'b1011110011 : begin
        result = input_755;
      end
      10'b1011110100 : begin
        result = input_756;
      end
      10'b1011110101 : begin
        result = input_757;
      end
      10'b1011110110 : begin
        result = input_758;
      end
      10'b1011110111 : begin
        result = input_759;
      end
      10'b1011111000 : begin
        result = input_760;
      end
      10'b1011111001 : begin
        result = input_761;
      end
      10'b1011111010 : begin
        result = input_762;
      end
      10'b1011111011 : begin
        result = input_763;
      end
      10'b1011111100 : begin
        result = input_764;
      end
      10'b1011111101 : begin
        result = input_765;
      end
      10'b1011111110 : begin
        result = input_766;
      end
      10'b1011111111 : begin
        result = input_767;
      end
      10'b1100000000 : begin
        result = input_768;
      end
      10'b1100000001 : begin
        result = input_769;
      end
      10'b1100000010 : begin
        result = input_770;
      end
      10'b1100000011 : begin
        result = input_771;
      end
      10'b1100000100 : begin
        result = input_772;
      end
      10'b1100000101 : begin
        result = input_773;
      end
      10'b1100000110 : begin
        result = input_774;
      end
      10'b1100000111 : begin
        result = input_775;
      end
      10'b1100001000 : begin
        result = input_776;
      end
      10'b1100001001 : begin
        result = input_777;
      end
      10'b1100001010 : begin
        result = input_778;
      end
      10'b1100001011 : begin
        result = input_779;
      end
      10'b1100001100 : begin
        result = input_780;
      end
      10'b1100001101 : begin
        result = input_781;
      end
      10'b1100001110 : begin
        result = input_782;
      end
      10'b1100001111 : begin
        result = input_783;
      end
      10'b1100010000 : begin
        result = input_784;
      end
      10'b1100010001 : begin
        result = input_785;
      end
      10'b1100010010 : begin
        result = input_786;
      end
      10'b1100010011 : begin
        result = input_787;
      end
      10'b1100010100 : begin
        result = input_788;
      end
      10'b1100010101 : begin
        result = input_789;
      end
      10'b1100010110 : begin
        result = input_790;
      end
      10'b1100010111 : begin
        result = input_791;
      end
      10'b1100011000 : begin
        result = input_792;
      end
      10'b1100011001 : begin
        result = input_793;
      end
      10'b1100011010 : begin
        result = input_794;
      end
      10'b1100011011 : begin
        result = input_795;
      end
      10'b1100011100 : begin
        result = input_796;
      end
      10'b1100011101 : begin
        result = input_797;
      end
      10'b1100011110 : begin
        result = input_798;
      end
      10'b1100011111 : begin
        result = input_799;
      end
      10'b1100100000 : begin
        result = input_800;
      end
      10'b1100100001 : begin
        result = input_801;
      end
      10'b1100100010 : begin
        result = input_802;
      end
      10'b1100100011 : begin
        result = input_803;
      end
      10'b1100100100 : begin
        result = input_804;
      end
      10'b1100100101 : begin
        result = input_805;
      end
      10'b1100100110 : begin
        result = input_806;
      end
      10'b1100100111 : begin
        result = input_807;
      end
      10'b1100101000 : begin
        result = input_808;
      end
      10'b1100101001 : begin
        result = input_809;
      end
      10'b1100101010 : begin
        result = input_810;
      end
      10'b1100101011 : begin
        result = input_811;
      end
      10'b1100101100 : begin
        result = input_812;
      end
      10'b1100101101 : begin
        result = input_813;
      end
      10'b1100101110 : begin
        result = input_814;
      end
      10'b1100101111 : begin
        result = input_815;
      end
      10'b1100110000 : begin
        result = input_816;
      end
      10'b1100110001 : begin
        result = input_817;
      end
      10'b1100110010 : begin
        result = input_818;
      end
      10'b1100110011 : begin
        result = input_819;
      end
      10'b1100110100 : begin
        result = input_820;
      end
      10'b1100110101 : begin
        result = input_821;
      end
      10'b1100110110 : begin
        result = input_822;
      end
      10'b1100110111 : begin
        result = input_823;
      end
      10'b1100111000 : begin
        result = input_824;
      end
      10'b1100111001 : begin
        result = input_825;
      end
      10'b1100111010 : begin
        result = input_826;
      end
      10'b1100111011 : begin
        result = input_827;
      end
      10'b1100111100 : begin
        result = input_828;
      end
      10'b1100111101 : begin
        result = input_829;
      end
      10'b1100111110 : begin
        result = input_830;
      end
      10'b1100111111 : begin
        result = input_831;
      end
      10'b1101000000 : begin
        result = input_832;
      end
      10'b1101000001 : begin
        result = input_833;
      end
      10'b1101000010 : begin
        result = input_834;
      end
      10'b1101000011 : begin
        result = input_835;
      end
      10'b1101000100 : begin
        result = input_836;
      end
      10'b1101000101 : begin
        result = input_837;
      end
      10'b1101000110 : begin
        result = input_838;
      end
      10'b1101000111 : begin
        result = input_839;
      end
      10'b1101001000 : begin
        result = input_840;
      end
      10'b1101001001 : begin
        result = input_841;
      end
      10'b1101001010 : begin
        result = input_842;
      end
      10'b1101001011 : begin
        result = input_843;
      end
      10'b1101001100 : begin
        result = input_844;
      end
      10'b1101001101 : begin
        result = input_845;
      end
      10'b1101001110 : begin
        result = input_846;
      end
      10'b1101001111 : begin
        result = input_847;
      end
      10'b1101010000 : begin
        result = input_848;
      end
      10'b1101010001 : begin
        result = input_849;
      end
      10'b1101010010 : begin
        result = input_850;
      end
      10'b1101010011 : begin
        result = input_851;
      end
      10'b1101010100 : begin
        result = input_852;
      end
      10'b1101010101 : begin
        result = input_853;
      end
      10'b1101010110 : begin
        result = input_854;
      end
      10'b1101010111 : begin
        result = input_855;
      end
      10'b1101011000 : begin
        result = input_856;
      end
      10'b1101011001 : begin
        result = input_857;
      end
      10'b1101011010 : begin
        result = input_858;
      end
      10'b1101011011 : begin
        result = input_859;
      end
      10'b1101011100 : begin
        result = input_860;
      end
      10'b1101011101 : begin
        result = input_861;
      end
      10'b1101011110 : begin
        result = input_862;
      end
      10'b1101011111 : begin
        result = input_863;
      end
      10'b1101100000 : begin
        result = input_864;
      end
      10'b1101100001 : begin
        result = input_865;
      end
      10'b1101100010 : begin
        result = input_866;
      end
      10'b1101100011 : begin
        result = input_867;
      end
      10'b1101100100 : begin
        result = input_868;
      end
      10'b1101100101 : begin
        result = input_869;
      end
      10'b1101100110 : begin
        result = input_870;
      end
      10'b1101100111 : begin
        result = input_871;
      end
      10'b1101101000 : begin
        result = input_872;
      end
      10'b1101101001 : begin
        result = input_873;
      end
      10'b1101101010 : begin
        result = input_874;
      end
      10'b1101101011 : begin
        result = input_875;
      end
      10'b1101101100 : begin
        result = input_876;
      end
      10'b1101101101 : begin
        result = input_877;
      end
      10'b1101101110 : begin
        result = input_878;
      end
      10'b1101101111 : begin
        result = input_879;
      end
      10'b1101110000 : begin
        result = input_880;
      end
      10'b1101110001 : begin
        result = input_881;
      end
      10'b1101110010 : begin
        result = input_882;
      end
      10'b1101110011 : begin
        result = input_883;
      end
      10'b1101110100 : begin
        result = input_884;
      end
      10'b1101110101 : begin
        result = input_885;
      end
      10'b1101110110 : begin
        result = input_886;
      end
      10'b1101110111 : begin
        result = input_887;
      end
      10'b1101111000 : begin
        result = input_888;
      end
      10'b1101111001 : begin
        result = input_889;
      end
      10'b1101111010 : begin
        result = input_890;
      end
      10'b1101111011 : begin
        result = input_891;
      end
      10'b1101111100 : begin
        result = input_892;
      end
      10'b1101111101 : begin
        result = input_893;
      end
      10'b1101111110 : begin
        result = input_894;
      end
      10'b1101111111 : begin
        result = input_895;
      end
      10'b1110000000 : begin
        result = input_896;
      end
      10'b1110000001 : begin
        result = input_897;
      end
      10'b1110000010 : begin
        result = input_898;
      end
      10'b1110000011 : begin
        result = input_899;
      end
      10'b1110000100 : begin
        result = input_900;
      end
      10'b1110000101 : begin
        result = input_901;
      end
      10'b1110000110 : begin
        result = input_902;
      end
      10'b1110000111 : begin
        result = input_903;
      end
      10'b1110001000 : begin
        result = input_904;
      end
      10'b1110001001 : begin
        result = input_905;
      end
      10'b1110001010 : begin
        result = input_906;
      end
      10'b1110001011 : begin
        result = input_907;
      end
      10'b1110001100 : begin
        result = input_908;
      end
      10'b1110001101 : begin
        result = input_909;
      end
      10'b1110001110 : begin
        result = input_910;
      end
      10'b1110001111 : begin
        result = input_911;
      end
      10'b1110010000 : begin
        result = input_912;
      end
      10'b1110010001 : begin
        result = input_913;
      end
      10'b1110010010 : begin
        result = input_914;
      end
      10'b1110010011 : begin
        result = input_915;
      end
      10'b1110010100 : begin
        result = input_916;
      end
      10'b1110010101 : begin
        result = input_917;
      end
      10'b1110010110 : begin
        result = input_918;
      end
      10'b1110010111 : begin
        result = input_919;
      end
      10'b1110011000 : begin
        result = input_920;
      end
      10'b1110011001 : begin
        result = input_921;
      end
      10'b1110011010 : begin
        result = input_922;
      end
      10'b1110011011 : begin
        result = input_923;
      end
      10'b1110011100 : begin
        result = input_924;
      end
      10'b1110011101 : begin
        result = input_925;
      end
      10'b1110011110 : begin
        result = input_926;
      end
      10'b1110011111 : begin
        result = input_927;
      end
      10'b1110100000 : begin
        result = input_928;
      end
      10'b1110100001 : begin
        result = input_929;
      end
      10'b1110100010 : begin
        result = input_930;
      end
      10'b1110100011 : begin
        result = input_931;
      end
      10'b1110100100 : begin
        result = input_932;
      end
      10'b1110100101 : begin
        result = input_933;
      end
      10'b1110100110 : begin
        result = input_934;
      end
      10'b1110100111 : begin
        result = input_935;
      end
      10'b1110101000 : begin
        result = input_936;
      end
      10'b1110101001 : begin
        result = input_937;
      end
      10'b1110101010 : begin
        result = input_938;
      end
      10'b1110101011 : begin
        result = input_939;
      end
      10'b1110101100 : begin
        result = input_940;
      end
      10'b1110101101 : begin
        result = input_941;
      end
      10'b1110101110 : begin
        result = input_942;
      end
      10'b1110101111 : begin
        result = input_943;
      end
      10'b1110110000 : begin
        result = input_944;
      end
      10'b1110110001 : begin
        result = input_945;
      end
      10'b1110110010 : begin
        result = input_946;
      end
      10'b1110110011 : begin
        result = input_947;
      end
      10'b1110110100 : begin
        result = input_948;
      end
      10'b1110110101 : begin
        result = input_949;
      end
      10'b1110110110 : begin
        result = input_950;
      end
      10'b1110110111 : begin
        result = input_951;
      end
      10'b1110111000 : begin
        result = input_952;
      end
      10'b1110111001 : begin
        result = input_953;
      end
      10'b1110111010 : begin
        result = input_954;
      end
      10'b1110111011 : begin
        result = input_955;
      end
      10'b1110111100 : begin
        result = input_956;
      end
      10'b1110111101 : begin
        result = input_957;
      end
      10'b1110111110 : begin
        result = input_958;
      end
      10'b1110111111 : begin
        result = input_959;
      end
      10'b1111000000 : begin
        result = input_960;
      end
      10'b1111000001 : begin
        result = input_961;
      end
      10'b1111000010 : begin
        result = input_962;
      end
      10'b1111000011 : begin
        result = input_963;
      end
      10'b1111000100 : begin
        result = input_964;
      end
      10'b1111000101 : begin
        result = input_965;
      end
      10'b1111000110 : begin
        result = input_966;
      end
      10'b1111000111 : begin
        result = input_967;
      end
      10'b1111001000 : begin
        result = input_968;
      end
      10'b1111001001 : begin
        result = input_969;
      end
      10'b1111001010 : begin
        result = input_970;
      end
      10'b1111001011 : begin
        result = input_971;
      end
      10'b1111001100 : begin
        result = input_972;
      end
      10'b1111001101 : begin
        result = input_973;
      end
      10'b1111001110 : begin
        result = input_974;
      end
      10'b1111001111 : begin
        result = input_975;
      end
      10'b1111010000 : begin
        result = input_976;
      end
      10'b1111010001 : begin
        result = input_977;
      end
      10'b1111010010 : begin
        result = input_978;
      end
      10'b1111010011 : begin
        result = input_979;
      end
      10'b1111010100 : begin
        result = input_980;
      end
      10'b1111010101 : begin
        result = input_981;
      end
      10'b1111010110 : begin
        result = input_982;
      end
      10'b1111010111 : begin
        result = input_983;
      end
      10'b1111011000 : begin
        result = input_984;
      end
      10'b1111011001 : begin
        result = input_985;
      end
      10'b1111011010 : begin
        result = input_986;
      end
      10'b1111011011 : begin
        result = input_987;
      end
      10'b1111011100 : begin
        result = input_988;
      end
      10'b1111011101 : begin
        result = input_989;
      end
      10'b1111011110 : begin
        result = input_990;
      end
      10'b1111011111 : begin
        result = input_991;
      end
      10'b1111100000 : begin
        result = input_992;
      end
      10'b1111100001 : begin
        result = input_993;
      end
      10'b1111100010 : begin
        result = input_994;
      end
      10'b1111100011 : begin
        result = input_995;
      end
      10'b1111100100 : begin
        result = input_996;
      end
      10'b1111100101 : begin
        result = input_997;
      end
      10'b1111100110 : begin
        result = input_998;
      end
      10'b1111100111 : begin
        result = input_999;
      end
      10'b1111101000 : begin
        result = input_1000;
      end
      10'b1111101001 : begin
        result = input_1001;
      end
      10'b1111101010 : begin
        result = input_1002;
      end
      10'b1111101011 : begin
        result = input_1003;
      end
      10'b1111101100 : begin
        result = input_1004;
      end
      10'b1111101101 : begin
        result = input_1005;
      end
      10'b1111101110 : begin
        result = input_1006;
      end
      10'b1111101111 : begin
        result = input_1007;
      end
      10'b1111110000 : begin
        result = input_1008;
      end
      10'b1111110001 : begin
        result = input_1009;
      end
      10'b1111110010 : begin
        result = input_1010;
      end
      10'b1111110011 : begin
        result = input_1011;
      end
      10'b1111110100 : begin
        result = input_1012;
      end
      10'b1111110101 : begin
        result = input_1013;
      end
      10'b1111110110 : begin
        result = input_1014;
      end
      10'b1111110111 : begin
        result = input_1015;
      end
      10'b1111111000 : begin
        result = input_1016;
      end
      10'b1111111001 : begin
        result = input_1017;
      end
      10'b1111111010 : begin
        result = input_1018;
      end
      10'b1111111011 : begin
        result = input_1019;
      end
      10'b1111111100 : begin
        result = input_1020;
      end
      10'b1111111101 : begin
        result = input_1021;
      end
      10'b1111111110 : begin
        result = input_1022;
      end
      default : begin
        result = input_1023;
      end
    endcase
    MUX_v_14_1024_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i10_1o14_281e23127cb7ddaedd69e0bbd10d0137bd_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Mon May 27 10:59:03 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i10_1o14_281e23127cb7ddaedd69e0bbd10d0137bd
// ------------------------------------------------------------------


module ROM_1i10_1o14_281e23127cb7ddaedd69e0bbd10d0137bd (
  I_1, O_1
);
  input [9:0] I_1;
  output [13:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_14_1024_2(14'b00111111111011, 14'b01111011010000, 14'b10101100110100,
      14'b10101111001000, 14'b01101100110000, 14'b01000011110110, 14'b01100010000011,
      14'b10011000011111, 14'b00011000110111, 14'b01100011111111, 14'b10010100000101,
      14'b01010010010010, 14'b00001001001010, 14'b01011011000001, 14'b01110101110010,
      14'b10010111101110, 14'b00010001101110, 14'b01100100000111, 14'b00011010101111,
      14'b00001111000101, 14'b01101110111011, 14'b01110111111010, 14'b00111010011111,
      14'b01100100101010, 14'b10100010101110, 14'b01111110100100, 14'b00011101011101,
      14'b00011010011000, 14'b00010101010100, 14'b10100001011001, 14'b10011110110100,
      14'b10001111011100, 14'b10111110110010, 14'b01100001100000, 14'b00001111100101,
      14'b00000001110101, 14'b01001010101111, 14'b01000100110111, 14'b00011000001101,
      14'b01101110100000, 14'b00101100001101, 14'b01100100111010, 14'b01000101001111,
      14'b10001010101101, 14'b01101111101000, 14'b00101000000100, 14'b01011000100000,
      14'b00111111001010, 14'b10111110011101, 14'b00000110110000, 14'b10100111111111,
      14'b00010011010101, 14'b01110110111010, 14'b00010111111110, 14'b00111110001111,
      14'b01111010110111, 14'b00100010000101, 14'b01100010100100, 14'b10001000010000,
      14'b01100110101010, 14'b01001011101011, 14'b00011010011010, 14'b00000000001110,
      14'b00111100100000, 14'b01010111000001, 14'b10010010011000, 14'b10111110000011,
      14'b00011111100011, 14'b01110101110111, 14'b00100100001011, 14'b01001001000001,
      14'b01110010101100, 14'b00011000010001, 14'b00010010000100, 14'b10000011010001,
      14'b10110001111101, 14'b00001111111100, 14'b00101110010111, 14'b10101000010100,
      14'b01101110000101, 14'b00110011110100, 14'b10101111100100, 14'b01010010100101,
      14'b10110100111010, 14'b10100110001101, 14'b10011101100110, 14'b10010100010101,
      14'b01100000100100, 14'b10010000111101, 14'b01011111110010, 14'b00110011111011,
      14'b00001101110011, 14'b10100011100101, 14'b00000111101001, 14'b00010111011110,
      14'b00101100100011, 14'b10101100110101, 14'b10011000000001, 14'b00101010110110,
      14'b10111111010001, 14'b01001101101010, 14'b10100011110001, 14'b10011101011110,
      14'b00010010101011, 14'b00001011011010, 14'b00011011100010, 14'b00111100001110,
      14'b00011111101110, 14'b01011100000100, 14'b10101010101010, 14'b10001100111100,
      14'b01010010011010, 14'b10001111011011, 14'b00111000010100, 14'b00111011000110,
      14'b10011111011110, 14'b00110001101100, 14'b00110110001011, 14'b01001000111100,
      14'b00100110001110, 14'b01110110111101, 14'b10010010101010, 14'b00001101000010,
      14'b01111000010111, 14'b01101010110100, 14'b00110101001011, 14'b01010011100111,
      14'b10111111110100, 14'b00110111111100, 14'b00011011001011, 14'b10101001000100,
      14'b10011000111011, 14'b10011111100001, 14'b00111111100110, 14'b10111111011010,
      14'b10000101001101, 14'b10100010100001, 14'b00101010111101, 14'b01110010101010,
      14'b10100101001110, 14'b01011110011000, 14'b00001110101111, 14'b10010001110010,
      14'b00010111000101, 14'b01101011010001, 14'b10010111000100, 14'b00111000000001,
      14'b01100111101001, 14'b10111101110001, 14'b00111111011111, 14'b00111001100100,
      14'b01111000000000, 14'b01111111111100, 14'b01101011110110, 14'b00110111001101,
      14'b10011001001111, 14'b01011111001010, 14'b00001011010111, 14'b10011101110011,
      14'b01101101011011, 14'b01101100100001, 14'b00011110011101, 14'b10011000000011,
      14'b10100100111111, 14'b01011110101001, 14'b00000101111010, 14'b01111010111111,
      14'b10001000111011, 14'b10001011000101, 14'b10010000001101, 14'b10001010001110,
      14'b01000111000111, 14'b10010101110101, 14'b10110110010000, 14'b01110111001110,
      14'b10001001110101, 14'b01011000110000, 14'b01001101011100, 14'b01100001101011,
      14'b10000011000100, 14'b10011110101100, 14'b10001000010011, 14'b00100100100101,
      14'b00110001010111, 14'b00010110111011, 14'b01010101010100, 14'b10000101101001,
      14'b01111001100111, 14'b00101001011001, 14'b00100100010000, 14'b10001101001100,
      14'b01100000101100, 14'b00001011100001, 14'b00111001110010, 14'b01001001011011,
      14'b01011001111001, 14'b10001101010110, 14'b00111001100111, 14'b00000000010000,
      14'b00001110010010, 14'b01010001000010, 14'b10100100100011, 14'b01000111001000,
      14'b00011110101100, 14'b00110110110101, 14'b10000011110100, 14'b01110101011100,
      14'b01010100000101, 14'b10100111101101, 14'b00110011010001, 14'b01101101111101,
      14'b00010000100100, 14'b00101101001111, 14'b01101111110100, 14'b10001010110111,
      14'b01010011101101, 14'b01100100001001, 14'b10000000000101, 14'b00101110010010,
      14'b01100011100111, 14'b01001111001000, 14'b01100111101010, 14'b01010111111001,
      14'b00000100010110, 14'b00001110100100, 14'b10011111110101, 14'b10001011011111,
      14'b01110111011010, 14'b00000101011111, 14'b10010001010010, 14'b00000011101101,
      14'b01011011100010, 14'b01111000001100, 14'b00110001001010, 14'b10111101011110,
      14'b01110110100010, 14'b00100000000101, 14'b10110000010101, 14'b00111011011010,
      14'b01010001010100, 14'b01000111111010, 14'b00011011010100, 14'b10110000100100,
      14'b00000101010100, 14'b00111001111111, 14'b01001000000110, 14'b00000100101100,
      14'b10101011110001, 14'b01001111001110, 14'b10011101000001, 14'b10110101100000,
      14'b10111111010111, 14'b01110011111101, 14'b10100111010011, 14'b01011001110010,
      14'b01011000010110, 14'b00111011111011, 14'b01010110110001, 14'b00010011001000,
      14'b10000100011100, 14'b10010000010101, 14'b00111100000101, 14'b00000011111010,
      14'b10101111001001, 14'b01000010000001, 14'b01100010110110, 14'b10010111010000,
      14'b10111111011110, 14'b01000000101000, 14'b00101011011010, 14'b00001010110100,
      14'b10001001101000, 14'b01100100001010, 14'b01101000111110, 14'b10011101111001,
      14'b10100010110010, 14'b00111010101111, 14'b01110010111100, 14'b10110001100001,
      14'b10000011110001, 14'b01100100100101, 14'b00111001000100, 14'b01100011000110,
      14'b10001100010010, 14'b01010100001111, 14'b00100011100000, 14'b01100101001100,
      14'b01110011111000, 14'b10000011100010, 14'b10101001001000, 14'b10111011010010,
      14'b01011001100101, 14'b00001101101100, 14'b01101101110110, 14'b00100001110111,
      14'b00100110000100, 14'b00110101110010, 14'b10010000000001, 14'b10000000001110,
      14'b01001011111010, 14'b01011101001100, 14'b00101010111010, 14'b01110000001010,
      14'b00010110011010, 14'b01110011011101, 14'b10001010101111, 14'b10100110100101,
      14'b10110011000001, 14'b01000001111100, 14'b00010110011000, 14'b10101001010000,
      14'b01000011101000, 14'b10000101101101, 14'b00011101001011, 14'b10010011101110,
      14'b00100101110000, 14'b00111011101000, 14'b10001101110100, 14'b00001010101110,
      14'b01010100010001, 14'b00100111011011, 14'b01000011110011, 14'b01011111100011,
      14'b00001001101011, 14'b00001110101001, 14'b00101100010010, 14'b01111001011111,
      14'b00110011001111, 14'b00100100111011, 14'b01110101000000, 14'b01011111100000,
      14'b01001111000000, 14'b00001100111000, 14'b10011111011100, 14'b10110110101010,
      14'b00010001011001, 14'b00101010100111, 14'b10011001111000, 14'b00001110000000,
      14'b00011111101100, 14'b01001111010011, 14'b00101001011110, 14'b10100011100000,
      14'b01111011001100, 14'b10111110001001, 14'b01010100111010, 14'b00101111111110,
      14'b01100100000000, 14'b10001110101100, 14'b10110110011000, 14'b10111101111001,
      14'b01000110101000, 14'b00010011111001, 14'b10011000001011, 14'b10110011001100,
      14'b10011011010001, 14'b10011100110111, 14'b10010111111000, 14'b00100011010110,
      14'b10010010110111, 14'b10101110111000, 14'b00000100111011, 14'b01000110011111,
      14'b00010010000110, 14'b01011110101101, 14'b01101001011111, 14'b10111001011001,
      14'b00000101100101, 14'b01110011000111, 14'b01000111000110, 14'b00001111010111,
      14'b10000101010110, 14'b10000010100000, 14'b10011110001110, 14'b01110101101010,
      14'b10010000100101, 14'b01000100001111, 14'b01010001100101, 14'b00111110011111,
      14'b10001001001001, 14'b00110001011001, 14'b01101101001110, 14'b01000000100010,
      14'b10110110000100, 14'b00110100101110, 14'b10110011010101, 14'b00011011011001,
      14'b00000100100100, 14'b10000111101001, 14'b00101011110110, 14'b10100010001010,
      14'b10111110011100, 14'b01011010101000, 14'b10111000100011, 14'b00110001101101,
      14'b00011111000100, 14'b00010000000000, 14'b10010001111100, 14'b00100110101101,
      14'b10101010110000, 14'b01000111100110, 14'b01101001011110, 14'b00111000100011,
      14'b01010101111111, 14'b01010001110001, 14'b00100110011111, 14'b10000100010110,
      14'b01110111100010, 14'b01111100011100, 14'b01100011111011, 14'b00010000101111,
      14'b00010011111000, 14'b00110110010010, 14'b10101100100101, 14'b00110011011011,
      14'b10110001010000, 14'b10000100110110, 14'b10010100000110, 14'b10011001101101,
      14'b00010011100101, 14'b00011101000001, 14'b01100001011001, 14'b01001001110000,
      14'b10110100101001, 14'b01011110010010, 14'b10011001011001, 14'b00110100001011,
      14'b00011100000101, 14'b00101100111111, 14'b01100001100010, 14'b01010001010000,
      14'b00100001000010, 14'b01111100011010, 14'b10010010001001, 14'b10110001100011,
      14'b01010101100011, 14'b01011111000100, 14'b10010110000001, 14'b01000000001100,
      14'b01110010011011, 14'b10100011000110, 14'b10010011111111, 14'b00010011110111,
      14'b00000110011000, 14'b01101011111111, 14'b00110000000111, 14'b00000101101000,
      14'b10000001010100, 14'b10110100001111, 14'b10001111000100, 14'b10001101011001,
      14'b10110100010011, 14'b00001101010010, 14'b10000110101001, 14'b00001100010000,
      14'b01111011101111, 14'b10000010001110, 14'b10111110001010, 14'b00011100110110,
      14'b10011111100101, 14'b10111110011000, 14'b01111010010011, 14'b10111001111111,
      14'b01010111100000, 14'b10011000110011, 14'b00001111110100, 14'b00001011010001,
      14'b00101011100000, 14'b01101000010100, 14'b01100110011000, 14'b01010011100100,
      14'b01000101001000, 14'b01101010100000, 14'b10000011010101, 14'b10011011100111,
      14'b01010000011110, 14'b00100100110100, 14'b01010110110000, 14'b01010010010011,
      14'b00010100110101, 14'b10001001100001, 14'b10010110111101, 14'b01110010001100,
      14'b01011010011100, 14'b01001100101110, 14'b00001110001101, 14'b10110101011101,
      14'b01000100101011, 14'b10000000101110, 14'b01101000011110, 14'b01000011001110,
      14'b00101111100100, 14'b00100011101101, 14'b10111111011001, 14'b00011110101011,
      14'b10010000000000, 14'b01000011001000, 14'b10111010001110, 14'b00001010110111,
      14'b01000100010011, 14'b10011001000001, 14'b01001100010100, 14'b00100101101011,
      14'b10011111110110, 14'b00101001011010, 14'b00001101001001, 14'b00111100110010,
      14'b10011111110111, 14'b01110001010000, 14'b10000100111001, 14'b10101110111100,
      14'b01101000100000, 14'b00111111011011, 14'b01011110101100, 14'b00111001100110,
      14'b01001001110010, 14'b10111001001101, 14'b01011010111000, 14'b01101110010010,
      14'b01101011010100, 14'b10101110000001, 14'b01111011110110, 14'b01001100011110,
      14'b10111111111100, 14'b01000000000110, 14'b00111101000100, 14'b00111000011010,
      14'b01100101111101, 14'b01111100000010, 14'b01111100101110, 14'b10111011001001,
      14'b01101001100011, 14'b00001000011001, 14'b01000111010010, 14'b00011001010111,
      14'b10000000100011, 14'b10110010111101, 14'b01110101111000, 14'b00001110001010,
      14'b10111000101000, 14'b10010101001100, 14'b10101001101010, 14'b10010111100111,
      14'b00101011111111, 14'b10110111011000, 14'b01101010011101, 14'b01101101000011,
      14'b00001100110011, 14'b10001011000111, 14'b01100001111111, 14'b10101001011011,
      14'b00000101011100, 14'b01110101011010, 14'b10000010010011, 14'b01100100100111,
      14'b00001010110110, 14'b00001101010100, 14'b01011000011011, 14'b00101011011101,
      14'b00111010000100, 14'b10110101000101, 14'b00101111010000, 14'b00010111110011,
      14'b10000111010011, 14'b01000000010010, 14'b10100111110010, 14'b00110011100111,
      14'b01011011111101, 14'b00101110100010, 14'b01110001111001, 14'b10111001101100,
      14'b10001110100011, 14'b10010001101011, 14'b10111000110110, 14'b00000001100010,
      14'b00100111011110, 14'b00100001000100, 14'b01000000100011, 14'b10110010001111,
      14'b00011100110100, 14'b00111000111101, 14'b00111101001100, 14'b01111111000101,
      14'b00100010110000, 14'b10101001110111, 14'b01111110011100, 14'b10010110110011,
      14'b01011101100101, 14'b01101111100100, 14'b10000100100000, 14'b00011010000110,
      14'b00000010011111, 14'b10101010101011, 14'b01001100110110, 14'b00000010000000,
      14'b01110010010000, 14'b00001011010101, 14'b10001111000101, 14'b01001110001110,
      14'b01100011111001, 14'b00110110100110, 14'b01011110011011, 14'b10101011011100,
      14'b01100000100101, 14'b10111000111110, 14'b00110101011111, 14'b10100100010010,
      14'b01110111110100, 14'b00111001101101, 14'b01101000000010, 14'b01101011111001,
      14'b10111010110001, 14'b10011111100100, 14'b10111010010010, 14'b10001110001101,
      14'b10000010101101, 14'b01001111110110, 14'b00000000101101, 14'b00100101100000,
      14'b00011110000001, 14'b01000100011001, 14'b00101010100000, 14'b00011010011111,
      14'b00000000110011, 14'b00101011111000, 14'b00001010001010, 14'b00011101101000,
      14'b10011100001101, 14'b10011011110011, 14'b10111011001100, 14'b01111110100010,
      14'b01001011100001, 14'b01000000100111, 14'b01000010100001, 14'b01011011001110,
      14'b01001010011101, 14'b10101011101001, 14'b10110100001100, 14'b00001001001110,
      14'b10111110100110, 14'b00000111100010, 14'b10111110001101, 14'b00011111010110,
      14'b01101110011000, 14'b10011100100010, 14'b00111101001000, 14'b10111011110000,
      14'b10100100010111, 14'b10110001100010, 14'b01101100101010, 14'b00100010100010,
      14'b00000100011100, 14'b01010100100101, 14'b01100111001001, 14'b00111100011001,
      14'b10100001100011, 14'b10101110110100, 14'b01100001010111, 14'b00001000000101,
      14'b10010101011100, 14'b10110000010001, 14'b00111100010111, 14'b00010010111010,
      14'b01000111111100, 14'b01111111100000, 14'b10110010110111, 14'b00000010011001,
      14'b01110000100100, 14'b01011010000011, 14'b01001111100001, 14'b10010000100000,
      14'b10111101111010, 14'b10110111100100, 14'b00010101001010, 14'b01101000010000,
      14'b00000010110011, 14'b01010110011100, 14'b00101001010110, 14'b01011100110101,
      14'b10111110011001, 14'b00001101011110, 14'b00110001010110, 14'b00000111011101,
      14'b01110001101111, 14'b01011000101110, 14'b01111011101010, 14'b01000010011110,
      14'b00000100101110, 14'b00101101001101, 14'b10011110000010, 14'b01101011101010,
      14'b10010101011000, 14'b10010110101111, 14'b10111010000001, 14'b01000000000010,
      14'b10011001100000, 14'b10100000011101, 14'b00010101001001, 14'b10100111011011,
      14'b01010011001101, 14'b01100001101110, 14'b00111101101111, 14'b00011100001111,
      14'b01100100110001, 14'b01010000100111, 14'b00010100011100, 14'b10000001111011,
      14'b00110101001100, 14'b00011101010101, 14'b00010011001111, 14'b00000001110000,
      14'b01100011111110, 14'b10110111001100, 14'b10111111110000, 14'b01110001110110,
      14'b00010110110011, 14'b10111111110010, 14'b10011010101000, 14'b00110110000000,
      14'b00001100100000, 14'b00010101110101, 14'b10100110110110, 14'b00000001100111,
      14'b01110011111100, 14'b01111100101000, 14'b00001110101000, 14'b00001011111100,
      14'b00001001111000, 14'b01111100111100, 14'b10000000011111, 14'b10000011111101,
      14'b01111001001110, 14'b10101001110110, 14'b10010101100011, 14'b00100111001100,
      14'b00011110011010, 14'b01100101111100, 14'b10011110101110, 14'b00010000010100,
      14'b01000011110010, 14'b00100110011001, 14'b00111000111001, 14'b00011001111011,
      14'b01000000101011, 14'b01001001010000, 14'b10011000000101, 14'b10101110001100,
      14'b00111101101010, 14'b00100000100010, 14'b01010010001101, 14'b00011111110100,
      14'b10111001001010, 14'b01110111010100, 14'b10111111001100, 14'b01010011110110,
      14'b00100101001100, 14'b00010101110111, 14'b01111000101000, 14'b00100000110100,
      14'b00110010010001, 14'b10101010100000, 14'b10001011000010, 14'b01110110011010,
      14'b10111011011011, 14'b00101011100111, 14'b00010010111111, 14'b00110100011011,
      14'b00101010010111, 14'b00100011011011, 14'b00011111010100, 14'b10000101111000,
      14'b10011111000000, 14'b00110010001110, 14'b00100100100001, 14'b00011011010110,
      14'b01001001111001, 14'b01001110000101, 14'b01110011110111, 14'b01100010101011,
      14'b10111100001100, 14'b01000100010110, 14'b01101111110101, 14'b01001011101100,
      14'b00000011010011, 14'b01111101000011, 14'b10011110101111, 14'b10010001001010,
      14'b10110011011001, 14'b00011011000111, 14'b00100100100000, 14'b01011010100001,
      14'b10011010010011, 14'b10000000000000, 14'b00001111011010, 14'b01110101100111,
      14'b00010101111001, 14'b00001101100110, 14'b00111000011111, 14'b10000100010001,
      14'b00101011000100, 14'b10011000101010, 14'b00011111110010, 14'b10011110111000,
      14'b00110011000000, 14'b01011111110100, 14'b00000000110110, 14'b00101101000000,
      14'b01001010011011, 14'b10111000011101, 14'b00110000000010, 14'b10000001011110,
      14'b10010011010100, 14'b01001100010001, 14'b01101100010101, 14'b00010001000010,
      14'b10011100110110, 14'b00101000000111, 14'b00001011000100, 14'b00001101111101,
      14'b01100101000001, 14'b01001101100010, 14'b10011100101000, 14'b00100000101010,
      14'b01011001010110, 14'b10100111110111, 14'b00001100001100, 14'b01001001111101,
      14'b01001000001111, 14'b00100001010110, 14'b00100000100111, 14'b01001011000010,
      14'b00001101110100, 14'b01010011111100, 14'b01011010100011, 14'b01011100110010,
      14'b01000011101101, 14'b01100110011111, 14'b01110101111101, 14'b01010010010101,
      14'b10100110101000, 14'b01000010011100, 14'b00110010111100, 14'b01011100011101,
      14'b10101000111110, 14'b01011010001000, 14'b10011011111111, 14'b01111110100000,
      14'b01111001101111, 14'b01101010010000, 14'b01110101000011, 14'b01100010000000,
      14'b00011101110011, 14'b10101011000011, 14'b01100010010001, 14'b10111000011011,
      14'b01011110010000, 14'b10110010111001, 14'b00010010010011, 14'b10001111110001,
      14'b01111011111101, 14'b00100110101111, 14'b01111100100010, 14'b10110001001001,
      14'b01101110010110, 14'b10001011001111, 14'b01101001001000, 14'b01100110001110,
      14'b01111110110010, 14'b10001001111100, 14'b01100111000011, 14'b00110111011001,
      14'b01000011111100, 14'b01001000000010, 14'b00100010011101, 14'b01101101010111,
      14'b01111110101010, 14'b01010110111000, 14'b10100010010110, 14'b10010001101001,
      14'b00100111000011, 14'b00100101101101, 14'b01110001101000, 14'b01101011100001,
      14'b10100101010110, 14'b10010001011100, 14'b10010011011101, 14'b00110111100010,
      14'b00110011111110, 14'b01011101100111, 14'b10111011000001, 14'b00110101010111,
      14'b10111111111011, 14'b10011001101110, 14'b10111100011111, 14'b01000011101100,
      14'b01111010010110, 14'b10110001000001, 14'b01100111001101, 14'b10111111101111,
      14'b00011111111100, 14'b10110101011011, 14'b01110010111001, 14'b10101111000001,
      14'b10110100111110, 14'b00111010010101, 14'b10001011101111, 14'b10011011111010,
      14'b00011001011011, 14'b01110000000000, 14'b00111101011111, 14'b01001110111010,
      14'b00101011001010, 14'b01110101001000, 14'b10100010001111, 14'b00001011110011,
      14'b00011001110110, 14'b10111100010101, 14'b01001101011000, 14'b10011110010110,
      14'b01000100101010, 14'b01100111000000, 14'b01111011011010, 14'b01110101001001,
      14'b10001011001000, 14'b10111011111101, 14'b00110111111101, 14'b10100111111100,
      14'b01011000101010, 14'b10100001110110, 14'b01001100100101, 14'b01110011110110,
      14'b10001001000011, 14'b00001011000110, 14'b01101001101100, 14'b10000100001110,
      14'b01110000011001, 14'b01010011111011, 14'b01110001101010, 14'b10101101001100,
      14'b00000100100010, 14'b01111010111000, 14'b01101010101011, 14'b10111000101110,
      14'b00100111001101, 14'b01100110110010, 14'b00111110111010, 14'b01011010101111,
      14'b00010110110010, 14'b01011001011001, 14'b01011010000010, 14'b01000001010010,
      14'b00100000111001, 14'b10110101100101, 14'b01001011110100, 14'b10001011000001,
      14'b00101100101000, 14'b10110011110110, 14'b10010000110000, 14'b00100111011000,
      14'b10001001001000, 14'b01101101100011, 14'b00101001010111, 14'b00011101101010,
      14'b01101101111111, 14'b01011100111110, 14'b10101110011011, 14'b01010101110000,
      14'b01100010000101, 14'b10001111011110, 14'b10110011000000, 14'b00001001111001,
      14'b10011100111110, 14'b10110100100010, 14'b01011000000001, 14'b10010101110011,
      14'b00100100011101, 14'b01101101100000, 14'b01101110101100, 14'b01001110110111,
      14'b01110000011111, 14'b10011010001001, 14'b10001100100101, 14'b00001000111001,
      14'b01100011110110, 14'b10101001011101, 14'b10010111001111, 14'b10000001001100,
      14'b10110011010000, 14'b01000001101011, 14'b00011111001101, 14'b00000000000010,
      14'b10010001110011, 14'b00000010100010, 14'b01100000100110, 14'b00011111010000,
      14'b00111001000001, 14'b10011001000000, 14'b01100011011011, 14'b01110110000101,
      14'b01100000101011, 14'b10000100111110, 14'b10011011001111, 14'b01010110100000,
      14'b10001100111011, 14'b00111001111010, 14'b10111011101001, 14'b00010110101100,
      14'b00101111111011, 14'b01010101110110, 14'b10010111011100, 14'b01001100000001,
      14'b01011110000011, 14'b01101111000010, 14'b10010110001010, 14'b01000111101100,
      14'b10011110110101, 14'b01100001110101, 14'b01011011111111, 14'b00101001011100,
      14'b10011110111100, 14'b00011000101100, 14'b10100010001011, 14'b01001000011110,
      14'b10011011011101, I_1);

  function automatic [13:0] MUX_v_14_1024_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [13:0] input_2;
    input [13:0] input_3;
    input [13:0] input_4;
    input [13:0] input_5;
    input [13:0] input_6;
    input [13:0] input_7;
    input [13:0] input_8;
    input [13:0] input_9;
    input [13:0] input_10;
    input [13:0] input_11;
    input [13:0] input_12;
    input [13:0] input_13;
    input [13:0] input_14;
    input [13:0] input_15;
    input [13:0] input_16;
    input [13:0] input_17;
    input [13:0] input_18;
    input [13:0] input_19;
    input [13:0] input_20;
    input [13:0] input_21;
    input [13:0] input_22;
    input [13:0] input_23;
    input [13:0] input_24;
    input [13:0] input_25;
    input [13:0] input_26;
    input [13:0] input_27;
    input [13:0] input_28;
    input [13:0] input_29;
    input [13:0] input_30;
    input [13:0] input_31;
    input [13:0] input_32;
    input [13:0] input_33;
    input [13:0] input_34;
    input [13:0] input_35;
    input [13:0] input_36;
    input [13:0] input_37;
    input [13:0] input_38;
    input [13:0] input_39;
    input [13:0] input_40;
    input [13:0] input_41;
    input [13:0] input_42;
    input [13:0] input_43;
    input [13:0] input_44;
    input [13:0] input_45;
    input [13:0] input_46;
    input [13:0] input_47;
    input [13:0] input_48;
    input [13:0] input_49;
    input [13:0] input_50;
    input [13:0] input_51;
    input [13:0] input_52;
    input [13:0] input_53;
    input [13:0] input_54;
    input [13:0] input_55;
    input [13:0] input_56;
    input [13:0] input_57;
    input [13:0] input_58;
    input [13:0] input_59;
    input [13:0] input_60;
    input [13:0] input_61;
    input [13:0] input_62;
    input [13:0] input_63;
    input [13:0] input_64;
    input [13:0] input_65;
    input [13:0] input_66;
    input [13:0] input_67;
    input [13:0] input_68;
    input [13:0] input_69;
    input [13:0] input_70;
    input [13:0] input_71;
    input [13:0] input_72;
    input [13:0] input_73;
    input [13:0] input_74;
    input [13:0] input_75;
    input [13:0] input_76;
    input [13:0] input_77;
    input [13:0] input_78;
    input [13:0] input_79;
    input [13:0] input_80;
    input [13:0] input_81;
    input [13:0] input_82;
    input [13:0] input_83;
    input [13:0] input_84;
    input [13:0] input_85;
    input [13:0] input_86;
    input [13:0] input_87;
    input [13:0] input_88;
    input [13:0] input_89;
    input [13:0] input_90;
    input [13:0] input_91;
    input [13:0] input_92;
    input [13:0] input_93;
    input [13:0] input_94;
    input [13:0] input_95;
    input [13:0] input_96;
    input [13:0] input_97;
    input [13:0] input_98;
    input [13:0] input_99;
    input [13:0] input_100;
    input [13:0] input_101;
    input [13:0] input_102;
    input [13:0] input_103;
    input [13:0] input_104;
    input [13:0] input_105;
    input [13:0] input_106;
    input [13:0] input_107;
    input [13:0] input_108;
    input [13:0] input_109;
    input [13:0] input_110;
    input [13:0] input_111;
    input [13:0] input_112;
    input [13:0] input_113;
    input [13:0] input_114;
    input [13:0] input_115;
    input [13:0] input_116;
    input [13:0] input_117;
    input [13:0] input_118;
    input [13:0] input_119;
    input [13:0] input_120;
    input [13:0] input_121;
    input [13:0] input_122;
    input [13:0] input_123;
    input [13:0] input_124;
    input [13:0] input_125;
    input [13:0] input_126;
    input [13:0] input_127;
    input [13:0] input_128;
    input [13:0] input_129;
    input [13:0] input_130;
    input [13:0] input_131;
    input [13:0] input_132;
    input [13:0] input_133;
    input [13:0] input_134;
    input [13:0] input_135;
    input [13:0] input_136;
    input [13:0] input_137;
    input [13:0] input_138;
    input [13:0] input_139;
    input [13:0] input_140;
    input [13:0] input_141;
    input [13:0] input_142;
    input [13:0] input_143;
    input [13:0] input_144;
    input [13:0] input_145;
    input [13:0] input_146;
    input [13:0] input_147;
    input [13:0] input_148;
    input [13:0] input_149;
    input [13:0] input_150;
    input [13:0] input_151;
    input [13:0] input_152;
    input [13:0] input_153;
    input [13:0] input_154;
    input [13:0] input_155;
    input [13:0] input_156;
    input [13:0] input_157;
    input [13:0] input_158;
    input [13:0] input_159;
    input [13:0] input_160;
    input [13:0] input_161;
    input [13:0] input_162;
    input [13:0] input_163;
    input [13:0] input_164;
    input [13:0] input_165;
    input [13:0] input_166;
    input [13:0] input_167;
    input [13:0] input_168;
    input [13:0] input_169;
    input [13:0] input_170;
    input [13:0] input_171;
    input [13:0] input_172;
    input [13:0] input_173;
    input [13:0] input_174;
    input [13:0] input_175;
    input [13:0] input_176;
    input [13:0] input_177;
    input [13:0] input_178;
    input [13:0] input_179;
    input [13:0] input_180;
    input [13:0] input_181;
    input [13:0] input_182;
    input [13:0] input_183;
    input [13:0] input_184;
    input [13:0] input_185;
    input [13:0] input_186;
    input [13:0] input_187;
    input [13:0] input_188;
    input [13:0] input_189;
    input [13:0] input_190;
    input [13:0] input_191;
    input [13:0] input_192;
    input [13:0] input_193;
    input [13:0] input_194;
    input [13:0] input_195;
    input [13:0] input_196;
    input [13:0] input_197;
    input [13:0] input_198;
    input [13:0] input_199;
    input [13:0] input_200;
    input [13:0] input_201;
    input [13:0] input_202;
    input [13:0] input_203;
    input [13:0] input_204;
    input [13:0] input_205;
    input [13:0] input_206;
    input [13:0] input_207;
    input [13:0] input_208;
    input [13:0] input_209;
    input [13:0] input_210;
    input [13:0] input_211;
    input [13:0] input_212;
    input [13:0] input_213;
    input [13:0] input_214;
    input [13:0] input_215;
    input [13:0] input_216;
    input [13:0] input_217;
    input [13:0] input_218;
    input [13:0] input_219;
    input [13:0] input_220;
    input [13:0] input_221;
    input [13:0] input_222;
    input [13:0] input_223;
    input [13:0] input_224;
    input [13:0] input_225;
    input [13:0] input_226;
    input [13:0] input_227;
    input [13:0] input_228;
    input [13:0] input_229;
    input [13:0] input_230;
    input [13:0] input_231;
    input [13:0] input_232;
    input [13:0] input_233;
    input [13:0] input_234;
    input [13:0] input_235;
    input [13:0] input_236;
    input [13:0] input_237;
    input [13:0] input_238;
    input [13:0] input_239;
    input [13:0] input_240;
    input [13:0] input_241;
    input [13:0] input_242;
    input [13:0] input_243;
    input [13:0] input_244;
    input [13:0] input_245;
    input [13:0] input_246;
    input [13:0] input_247;
    input [13:0] input_248;
    input [13:0] input_249;
    input [13:0] input_250;
    input [13:0] input_251;
    input [13:0] input_252;
    input [13:0] input_253;
    input [13:0] input_254;
    input [13:0] input_255;
    input [13:0] input_256;
    input [13:0] input_257;
    input [13:0] input_258;
    input [13:0] input_259;
    input [13:0] input_260;
    input [13:0] input_261;
    input [13:0] input_262;
    input [13:0] input_263;
    input [13:0] input_264;
    input [13:0] input_265;
    input [13:0] input_266;
    input [13:0] input_267;
    input [13:0] input_268;
    input [13:0] input_269;
    input [13:0] input_270;
    input [13:0] input_271;
    input [13:0] input_272;
    input [13:0] input_273;
    input [13:0] input_274;
    input [13:0] input_275;
    input [13:0] input_276;
    input [13:0] input_277;
    input [13:0] input_278;
    input [13:0] input_279;
    input [13:0] input_280;
    input [13:0] input_281;
    input [13:0] input_282;
    input [13:0] input_283;
    input [13:0] input_284;
    input [13:0] input_285;
    input [13:0] input_286;
    input [13:0] input_287;
    input [13:0] input_288;
    input [13:0] input_289;
    input [13:0] input_290;
    input [13:0] input_291;
    input [13:0] input_292;
    input [13:0] input_293;
    input [13:0] input_294;
    input [13:0] input_295;
    input [13:0] input_296;
    input [13:0] input_297;
    input [13:0] input_298;
    input [13:0] input_299;
    input [13:0] input_300;
    input [13:0] input_301;
    input [13:0] input_302;
    input [13:0] input_303;
    input [13:0] input_304;
    input [13:0] input_305;
    input [13:0] input_306;
    input [13:0] input_307;
    input [13:0] input_308;
    input [13:0] input_309;
    input [13:0] input_310;
    input [13:0] input_311;
    input [13:0] input_312;
    input [13:0] input_313;
    input [13:0] input_314;
    input [13:0] input_315;
    input [13:0] input_316;
    input [13:0] input_317;
    input [13:0] input_318;
    input [13:0] input_319;
    input [13:0] input_320;
    input [13:0] input_321;
    input [13:0] input_322;
    input [13:0] input_323;
    input [13:0] input_324;
    input [13:0] input_325;
    input [13:0] input_326;
    input [13:0] input_327;
    input [13:0] input_328;
    input [13:0] input_329;
    input [13:0] input_330;
    input [13:0] input_331;
    input [13:0] input_332;
    input [13:0] input_333;
    input [13:0] input_334;
    input [13:0] input_335;
    input [13:0] input_336;
    input [13:0] input_337;
    input [13:0] input_338;
    input [13:0] input_339;
    input [13:0] input_340;
    input [13:0] input_341;
    input [13:0] input_342;
    input [13:0] input_343;
    input [13:0] input_344;
    input [13:0] input_345;
    input [13:0] input_346;
    input [13:0] input_347;
    input [13:0] input_348;
    input [13:0] input_349;
    input [13:0] input_350;
    input [13:0] input_351;
    input [13:0] input_352;
    input [13:0] input_353;
    input [13:0] input_354;
    input [13:0] input_355;
    input [13:0] input_356;
    input [13:0] input_357;
    input [13:0] input_358;
    input [13:0] input_359;
    input [13:0] input_360;
    input [13:0] input_361;
    input [13:0] input_362;
    input [13:0] input_363;
    input [13:0] input_364;
    input [13:0] input_365;
    input [13:0] input_366;
    input [13:0] input_367;
    input [13:0] input_368;
    input [13:0] input_369;
    input [13:0] input_370;
    input [13:0] input_371;
    input [13:0] input_372;
    input [13:0] input_373;
    input [13:0] input_374;
    input [13:0] input_375;
    input [13:0] input_376;
    input [13:0] input_377;
    input [13:0] input_378;
    input [13:0] input_379;
    input [13:0] input_380;
    input [13:0] input_381;
    input [13:0] input_382;
    input [13:0] input_383;
    input [13:0] input_384;
    input [13:0] input_385;
    input [13:0] input_386;
    input [13:0] input_387;
    input [13:0] input_388;
    input [13:0] input_389;
    input [13:0] input_390;
    input [13:0] input_391;
    input [13:0] input_392;
    input [13:0] input_393;
    input [13:0] input_394;
    input [13:0] input_395;
    input [13:0] input_396;
    input [13:0] input_397;
    input [13:0] input_398;
    input [13:0] input_399;
    input [13:0] input_400;
    input [13:0] input_401;
    input [13:0] input_402;
    input [13:0] input_403;
    input [13:0] input_404;
    input [13:0] input_405;
    input [13:0] input_406;
    input [13:0] input_407;
    input [13:0] input_408;
    input [13:0] input_409;
    input [13:0] input_410;
    input [13:0] input_411;
    input [13:0] input_412;
    input [13:0] input_413;
    input [13:0] input_414;
    input [13:0] input_415;
    input [13:0] input_416;
    input [13:0] input_417;
    input [13:0] input_418;
    input [13:0] input_419;
    input [13:0] input_420;
    input [13:0] input_421;
    input [13:0] input_422;
    input [13:0] input_423;
    input [13:0] input_424;
    input [13:0] input_425;
    input [13:0] input_426;
    input [13:0] input_427;
    input [13:0] input_428;
    input [13:0] input_429;
    input [13:0] input_430;
    input [13:0] input_431;
    input [13:0] input_432;
    input [13:0] input_433;
    input [13:0] input_434;
    input [13:0] input_435;
    input [13:0] input_436;
    input [13:0] input_437;
    input [13:0] input_438;
    input [13:0] input_439;
    input [13:0] input_440;
    input [13:0] input_441;
    input [13:0] input_442;
    input [13:0] input_443;
    input [13:0] input_444;
    input [13:0] input_445;
    input [13:0] input_446;
    input [13:0] input_447;
    input [13:0] input_448;
    input [13:0] input_449;
    input [13:0] input_450;
    input [13:0] input_451;
    input [13:0] input_452;
    input [13:0] input_453;
    input [13:0] input_454;
    input [13:0] input_455;
    input [13:0] input_456;
    input [13:0] input_457;
    input [13:0] input_458;
    input [13:0] input_459;
    input [13:0] input_460;
    input [13:0] input_461;
    input [13:0] input_462;
    input [13:0] input_463;
    input [13:0] input_464;
    input [13:0] input_465;
    input [13:0] input_466;
    input [13:0] input_467;
    input [13:0] input_468;
    input [13:0] input_469;
    input [13:0] input_470;
    input [13:0] input_471;
    input [13:0] input_472;
    input [13:0] input_473;
    input [13:0] input_474;
    input [13:0] input_475;
    input [13:0] input_476;
    input [13:0] input_477;
    input [13:0] input_478;
    input [13:0] input_479;
    input [13:0] input_480;
    input [13:0] input_481;
    input [13:0] input_482;
    input [13:0] input_483;
    input [13:0] input_484;
    input [13:0] input_485;
    input [13:0] input_486;
    input [13:0] input_487;
    input [13:0] input_488;
    input [13:0] input_489;
    input [13:0] input_490;
    input [13:0] input_491;
    input [13:0] input_492;
    input [13:0] input_493;
    input [13:0] input_494;
    input [13:0] input_495;
    input [13:0] input_496;
    input [13:0] input_497;
    input [13:0] input_498;
    input [13:0] input_499;
    input [13:0] input_500;
    input [13:0] input_501;
    input [13:0] input_502;
    input [13:0] input_503;
    input [13:0] input_504;
    input [13:0] input_505;
    input [13:0] input_506;
    input [13:0] input_507;
    input [13:0] input_508;
    input [13:0] input_509;
    input [13:0] input_510;
    input [13:0] input_511;
    input [13:0] input_512;
    input [13:0] input_513;
    input [13:0] input_514;
    input [13:0] input_515;
    input [13:0] input_516;
    input [13:0] input_517;
    input [13:0] input_518;
    input [13:0] input_519;
    input [13:0] input_520;
    input [13:0] input_521;
    input [13:0] input_522;
    input [13:0] input_523;
    input [13:0] input_524;
    input [13:0] input_525;
    input [13:0] input_526;
    input [13:0] input_527;
    input [13:0] input_528;
    input [13:0] input_529;
    input [13:0] input_530;
    input [13:0] input_531;
    input [13:0] input_532;
    input [13:0] input_533;
    input [13:0] input_534;
    input [13:0] input_535;
    input [13:0] input_536;
    input [13:0] input_537;
    input [13:0] input_538;
    input [13:0] input_539;
    input [13:0] input_540;
    input [13:0] input_541;
    input [13:0] input_542;
    input [13:0] input_543;
    input [13:0] input_544;
    input [13:0] input_545;
    input [13:0] input_546;
    input [13:0] input_547;
    input [13:0] input_548;
    input [13:0] input_549;
    input [13:0] input_550;
    input [13:0] input_551;
    input [13:0] input_552;
    input [13:0] input_553;
    input [13:0] input_554;
    input [13:0] input_555;
    input [13:0] input_556;
    input [13:0] input_557;
    input [13:0] input_558;
    input [13:0] input_559;
    input [13:0] input_560;
    input [13:0] input_561;
    input [13:0] input_562;
    input [13:0] input_563;
    input [13:0] input_564;
    input [13:0] input_565;
    input [13:0] input_566;
    input [13:0] input_567;
    input [13:0] input_568;
    input [13:0] input_569;
    input [13:0] input_570;
    input [13:0] input_571;
    input [13:0] input_572;
    input [13:0] input_573;
    input [13:0] input_574;
    input [13:0] input_575;
    input [13:0] input_576;
    input [13:0] input_577;
    input [13:0] input_578;
    input [13:0] input_579;
    input [13:0] input_580;
    input [13:0] input_581;
    input [13:0] input_582;
    input [13:0] input_583;
    input [13:0] input_584;
    input [13:0] input_585;
    input [13:0] input_586;
    input [13:0] input_587;
    input [13:0] input_588;
    input [13:0] input_589;
    input [13:0] input_590;
    input [13:0] input_591;
    input [13:0] input_592;
    input [13:0] input_593;
    input [13:0] input_594;
    input [13:0] input_595;
    input [13:0] input_596;
    input [13:0] input_597;
    input [13:0] input_598;
    input [13:0] input_599;
    input [13:0] input_600;
    input [13:0] input_601;
    input [13:0] input_602;
    input [13:0] input_603;
    input [13:0] input_604;
    input [13:0] input_605;
    input [13:0] input_606;
    input [13:0] input_607;
    input [13:0] input_608;
    input [13:0] input_609;
    input [13:0] input_610;
    input [13:0] input_611;
    input [13:0] input_612;
    input [13:0] input_613;
    input [13:0] input_614;
    input [13:0] input_615;
    input [13:0] input_616;
    input [13:0] input_617;
    input [13:0] input_618;
    input [13:0] input_619;
    input [13:0] input_620;
    input [13:0] input_621;
    input [13:0] input_622;
    input [13:0] input_623;
    input [13:0] input_624;
    input [13:0] input_625;
    input [13:0] input_626;
    input [13:0] input_627;
    input [13:0] input_628;
    input [13:0] input_629;
    input [13:0] input_630;
    input [13:0] input_631;
    input [13:0] input_632;
    input [13:0] input_633;
    input [13:0] input_634;
    input [13:0] input_635;
    input [13:0] input_636;
    input [13:0] input_637;
    input [13:0] input_638;
    input [13:0] input_639;
    input [13:0] input_640;
    input [13:0] input_641;
    input [13:0] input_642;
    input [13:0] input_643;
    input [13:0] input_644;
    input [13:0] input_645;
    input [13:0] input_646;
    input [13:0] input_647;
    input [13:0] input_648;
    input [13:0] input_649;
    input [13:0] input_650;
    input [13:0] input_651;
    input [13:0] input_652;
    input [13:0] input_653;
    input [13:0] input_654;
    input [13:0] input_655;
    input [13:0] input_656;
    input [13:0] input_657;
    input [13:0] input_658;
    input [13:0] input_659;
    input [13:0] input_660;
    input [13:0] input_661;
    input [13:0] input_662;
    input [13:0] input_663;
    input [13:0] input_664;
    input [13:0] input_665;
    input [13:0] input_666;
    input [13:0] input_667;
    input [13:0] input_668;
    input [13:0] input_669;
    input [13:0] input_670;
    input [13:0] input_671;
    input [13:0] input_672;
    input [13:0] input_673;
    input [13:0] input_674;
    input [13:0] input_675;
    input [13:0] input_676;
    input [13:0] input_677;
    input [13:0] input_678;
    input [13:0] input_679;
    input [13:0] input_680;
    input [13:0] input_681;
    input [13:0] input_682;
    input [13:0] input_683;
    input [13:0] input_684;
    input [13:0] input_685;
    input [13:0] input_686;
    input [13:0] input_687;
    input [13:0] input_688;
    input [13:0] input_689;
    input [13:0] input_690;
    input [13:0] input_691;
    input [13:0] input_692;
    input [13:0] input_693;
    input [13:0] input_694;
    input [13:0] input_695;
    input [13:0] input_696;
    input [13:0] input_697;
    input [13:0] input_698;
    input [13:0] input_699;
    input [13:0] input_700;
    input [13:0] input_701;
    input [13:0] input_702;
    input [13:0] input_703;
    input [13:0] input_704;
    input [13:0] input_705;
    input [13:0] input_706;
    input [13:0] input_707;
    input [13:0] input_708;
    input [13:0] input_709;
    input [13:0] input_710;
    input [13:0] input_711;
    input [13:0] input_712;
    input [13:0] input_713;
    input [13:0] input_714;
    input [13:0] input_715;
    input [13:0] input_716;
    input [13:0] input_717;
    input [13:0] input_718;
    input [13:0] input_719;
    input [13:0] input_720;
    input [13:0] input_721;
    input [13:0] input_722;
    input [13:0] input_723;
    input [13:0] input_724;
    input [13:0] input_725;
    input [13:0] input_726;
    input [13:0] input_727;
    input [13:0] input_728;
    input [13:0] input_729;
    input [13:0] input_730;
    input [13:0] input_731;
    input [13:0] input_732;
    input [13:0] input_733;
    input [13:0] input_734;
    input [13:0] input_735;
    input [13:0] input_736;
    input [13:0] input_737;
    input [13:0] input_738;
    input [13:0] input_739;
    input [13:0] input_740;
    input [13:0] input_741;
    input [13:0] input_742;
    input [13:0] input_743;
    input [13:0] input_744;
    input [13:0] input_745;
    input [13:0] input_746;
    input [13:0] input_747;
    input [13:0] input_748;
    input [13:0] input_749;
    input [13:0] input_750;
    input [13:0] input_751;
    input [13:0] input_752;
    input [13:0] input_753;
    input [13:0] input_754;
    input [13:0] input_755;
    input [13:0] input_756;
    input [13:0] input_757;
    input [13:0] input_758;
    input [13:0] input_759;
    input [13:0] input_760;
    input [13:0] input_761;
    input [13:0] input_762;
    input [13:0] input_763;
    input [13:0] input_764;
    input [13:0] input_765;
    input [13:0] input_766;
    input [13:0] input_767;
    input [13:0] input_768;
    input [13:0] input_769;
    input [13:0] input_770;
    input [13:0] input_771;
    input [13:0] input_772;
    input [13:0] input_773;
    input [13:0] input_774;
    input [13:0] input_775;
    input [13:0] input_776;
    input [13:0] input_777;
    input [13:0] input_778;
    input [13:0] input_779;
    input [13:0] input_780;
    input [13:0] input_781;
    input [13:0] input_782;
    input [13:0] input_783;
    input [13:0] input_784;
    input [13:0] input_785;
    input [13:0] input_786;
    input [13:0] input_787;
    input [13:0] input_788;
    input [13:0] input_789;
    input [13:0] input_790;
    input [13:0] input_791;
    input [13:0] input_792;
    input [13:0] input_793;
    input [13:0] input_794;
    input [13:0] input_795;
    input [13:0] input_796;
    input [13:0] input_797;
    input [13:0] input_798;
    input [13:0] input_799;
    input [13:0] input_800;
    input [13:0] input_801;
    input [13:0] input_802;
    input [13:0] input_803;
    input [13:0] input_804;
    input [13:0] input_805;
    input [13:0] input_806;
    input [13:0] input_807;
    input [13:0] input_808;
    input [13:0] input_809;
    input [13:0] input_810;
    input [13:0] input_811;
    input [13:0] input_812;
    input [13:0] input_813;
    input [13:0] input_814;
    input [13:0] input_815;
    input [13:0] input_816;
    input [13:0] input_817;
    input [13:0] input_818;
    input [13:0] input_819;
    input [13:0] input_820;
    input [13:0] input_821;
    input [13:0] input_822;
    input [13:0] input_823;
    input [13:0] input_824;
    input [13:0] input_825;
    input [13:0] input_826;
    input [13:0] input_827;
    input [13:0] input_828;
    input [13:0] input_829;
    input [13:0] input_830;
    input [13:0] input_831;
    input [13:0] input_832;
    input [13:0] input_833;
    input [13:0] input_834;
    input [13:0] input_835;
    input [13:0] input_836;
    input [13:0] input_837;
    input [13:0] input_838;
    input [13:0] input_839;
    input [13:0] input_840;
    input [13:0] input_841;
    input [13:0] input_842;
    input [13:0] input_843;
    input [13:0] input_844;
    input [13:0] input_845;
    input [13:0] input_846;
    input [13:0] input_847;
    input [13:0] input_848;
    input [13:0] input_849;
    input [13:0] input_850;
    input [13:0] input_851;
    input [13:0] input_852;
    input [13:0] input_853;
    input [13:0] input_854;
    input [13:0] input_855;
    input [13:0] input_856;
    input [13:0] input_857;
    input [13:0] input_858;
    input [13:0] input_859;
    input [13:0] input_860;
    input [13:0] input_861;
    input [13:0] input_862;
    input [13:0] input_863;
    input [13:0] input_864;
    input [13:0] input_865;
    input [13:0] input_866;
    input [13:0] input_867;
    input [13:0] input_868;
    input [13:0] input_869;
    input [13:0] input_870;
    input [13:0] input_871;
    input [13:0] input_872;
    input [13:0] input_873;
    input [13:0] input_874;
    input [13:0] input_875;
    input [13:0] input_876;
    input [13:0] input_877;
    input [13:0] input_878;
    input [13:0] input_879;
    input [13:0] input_880;
    input [13:0] input_881;
    input [13:0] input_882;
    input [13:0] input_883;
    input [13:0] input_884;
    input [13:0] input_885;
    input [13:0] input_886;
    input [13:0] input_887;
    input [13:0] input_888;
    input [13:0] input_889;
    input [13:0] input_890;
    input [13:0] input_891;
    input [13:0] input_892;
    input [13:0] input_893;
    input [13:0] input_894;
    input [13:0] input_895;
    input [13:0] input_896;
    input [13:0] input_897;
    input [13:0] input_898;
    input [13:0] input_899;
    input [13:0] input_900;
    input [13:0] input_901;
    input [13:0] input_902;
    input [13:0] input_903;
    input [13:0] input_904;
    input [13:0] input_905;
    input [13:0] input_906;
    input [13:0] input_907;
    input [13:0] input_908;
    input [13:0] input_909;
    input [13:0] input_910;
    input [13:0] input_911;
    input [13:0] input_912;
    input [13:0] input_913;
    input [13:0] input_914;
    input [13:0] input_915;
    input [13:0] input_916;
    input [13:0] input_917;
    input [13:0] input_918;
    input [13:0] input_919;
    input [13:0] input_920;
    input [13:0] input_921;
    input [13:0] input_922;
    input [13:0] input_923;
    input [13:0] input_924;
    input [13:0] input_925;
    input [13:0] input_926;
    input [13:0] input_927;
    input [13:0] input_928;
    input [13:0] input_929;
    input [13:0] input_930;
    input [13:0] input_931;
    input [13:0] input_932;
    input [13:0] input_933;
    input [13:0] input_934;
    input [13:0] input_935;
    input [13:0] input_936;
    input [13:0] input_937;
    input [13:0] input_938;
    input [13:0] input_939;
    input [13:0] input_940;
    input [13:0] input_941;
    input [13:0] input_942;
    input [13:0] input_943;
    input [13:0] input_944;
    input [13:0] input_945;
    input [13:0] input_946;
    input [13:0] input_947;
    input [13:0] input_948;
    input [13:0] input_949;
    input [13:0] input_950;
    input [13:0] input_951;
    input [13:0] input_952;
    input [13:0] input_953;
    input [13:0] input_954;
    input [13:0] input_955;
    input [13:0] input_956;
    input [13:0] input_957;
    input [13:0] input_958;
    input [13:0] input_959;
    input [13:0] input_960;
    input [13:0] input_961;
    input [13:0] input_962;
    input [13:0] input_963;
    input [13:0] input_964;
    input [13:0] input_965;
    input [13:0] input_966;
    input [13:0] input_967;
    input [13:0] input_968;
    input [13:0] input_969;
    input [13:0] input_970;
    input [13:0] input_971;
    input [13:0] input_972;
    input [13:0] input_973;
    input [13:0] input_974;
    input [13:0] input_975;
    input [13:0] input_976;
    input [13:0] input_977;
    input [13:0] input_978;
    input [13:0] input_979;
    input [13:0] input_980;
    input [13:0] input_981;
    input [13:0] input_982;
    input [13:0] input_983;
    input [13:0] input_984;
    input [13:0] input_985;
    input [13:0] input_986;
    input [13:0] input_987;
    input [13:0] input_988;
    input [13:0] input_989;
    input [13:0] input_990;
    input [13:0] input_991;
    input [13:0] input_992;
    input [13:0] input_993;
    input [13:0] input_994;
    input [13:0] input_995;
    input [13:0] input_996;
    input [13:0] input_997;
    input [13:0] input_998;
    input [13:0] input_999;
    input [13:0] input_1000;
    input [13:0] input_1001;
    input [13:0] input_1002;
    input [13:0] input_1003;
    input [13:0] input_1004;
    input [13:0] input_1005;
    input [13:0] input_1006;
    input [13:0] input_1007;
    input [13:0] input_1008;
    input [13:0] input_1009;
    input [13:0] input_1010;
    input [13:0] input_1011;
    input [13:0] input_1012;
    input [13:0] input_1013;
    input [13:0] input_1014;
    input [13:0] input_1015;
    input [13:0] input_1016;
    input [13:0] input_1017;
    input [13:0] input_1018;
    input [13:0] input_1019;
    input [13:0] input_1020;
    input [13:0] input_1021;
    input [13:0] input_1022;
    input [13:0] input_1023;
    input [9:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      10'b0000000000 : begin
        result = input_0;
      end
      10'b0000000001 : begin
        result = input_1;
      end
      10'b0000000010 : begin
        result = input_2;
      end
      10'b0000000011 : begin
        result = input_3;
      end
      10'b0000000100 : begin
        result = input_4;
      end
      10'b0000000101 : begin
        result = input_5;
      end
      10'b0000000110 : begin
        result = input_6;
      end
      10'b0000000111 : begin
        result = input_7;
      end
      10'b0000001000 : begin
        result = input_8;
      end
      10'b0000001001 : begin
        result = input_9;
      end
      10'b0000001010 : begin
        result = input_10;
      end
      10'b0000001011 : begin
        result = input_11;
      end
      10'b0000001100 : begin
        result = input_12;
      end
      10'b0000001101 : begin
        result = input_13;
      end
      10'b0000001110 : begin
        result = input_14;
      end
      10'b0000001111 : begin
        result = input_15;
      end
      10'b0000010000 : begin
        result = input_16;
      end
      10'b0000010001 : begin
        result = input_17;
      end
      10'b0000010010 : begin
        result = input_18;
      end
      10'b0000010011 : begin
        result = input_19;
      end
      10'b0000010100 : begin
        result = input_20;
      end
      10'b0000010101 : begin
        result = input_21;
      end
      10'b0000010110 : begin
        result = input_22;
      end
      10'b0000010111 : begin
        result = input_23;
      end
      10'b0000011000 : begin
        result = input_24;
      end
      10'b0000011001 : begin
        result = input_25;
      end
      10'b0000011010 : begin
        result = input_26;
      end
      10'b0000011011 : begin
        result = input_27;
      end
      10'b0000011100 : begin
        result = input_28;
      end
      10'b0000011101 : begin
        result = input_29;
      end
      10'b0000011110 : begin
        result = input_30;
      end
      10'b0000011111 : begin
        result = input_31;
      end
      10'b0000100000 : begin
        result = input_32;
      end
      10'b0000100001 : begin
        result = input_33;
      end
      10'b0000100010 : begin
        result = input_34;
      end
      10'b0000100011 : begin
        result = input_35;
      end
      10'b0000100100 : begin
        result = input_36;
      end
      10'b0000100101 : begin
        result = input_37;
      end
      10'b0000100110 : begin
        result = input_38;
      end
      10'b0000100111 : begin
        result = input_39;
      end
      10'b0000101000 : begin
        result = input_40;
      end
      10'b0000101001 : begin
        result = input_41;
      end
      10'b0000101010 : begin
        result = input_42;
      end
      10'b0000101011 : begin
        result = input_43;
      end
      10'b0000101100 : begin
        result = input_44;
      end
      10'b0000101101 : begin
        result = input_45;
      end
      10'b0000101110 : begin
        result = input_46;
      end
      10'b0000101111 : begin
        result = input_47;
      end
      10'b0000110000 : begin
        result = input_48;
      end
      10'b0000110001 : begin
        result = input_49;
      end
      10'b0000110010 : begin
        result = input_50;
      end
      10'b0000110011 : begin
        result = input_51;
      end
      10'b0000110100 : begin
        result = input_52;
      end
      10'b0000110101 : begin
        result = input_53;
      end
      10'b0000110110 : begin
        result = input_54;
      end
      10'b0000110111 : begin
        result = input_55;
      end
      10'b0000111000 : begin
        result = input_56;
      end
      10'b0000111001 : begin
        result = input_57;
      end
      10'b0000111010 : begin
        result = input_58;
      end
      10'b0000111011 : begin
        result = input_59;
      end
      10'b0000111100 : begin
        result = input_60;
      end
      10'b0000111101 : begin
        result = input_61;
      end
      10'b0000111110 : begin
        result = input_62;
      end
      10'b0000111111 : begin
        result = input_63;
      end
      10'b0001000000 : begin
        result = input_64;
      end
      10'b0001000001 : begin
        result = input_65;
      end
      10'b0001000010 : begin
        result = input_66;
      end
      10'b0001000011 : begin
        result = input_67;
      end
      10'b0001000100 : begin
        result = input_68;
      end
      10'b0001000101 : begin
        result = input_69;
      end
      10'b0001000110 : begin
        result = input_70;
      end
      10'b0001000111 : begin
        result = input_71;
      end
      10'b0001001000 : begin
        result = input_72;
      end
      10'b0001001001 : begin
        result = input_73;
      end
      10'b0001001010 : begin
        result = input_74;
      end
      10'b0001001011 : begin
        result = input_75;
      end
      10'b0001001100 : begin
        result = input_76;
      end
      10'b0001001101 : begin
        result = input_77;
      end
      10'b0001001110 : begin
        result = input_78;
      end
      10'b0001001111 : begin
        result = input_79;
      end
      10'b0001010000 : begin
        result = input_80;
      end
      10'b0001010001 : begin
        result = input_81;
      end
      10'b0001010010 : begin
        result = input_82;
      end
      10'b0001010011 : begin
        result = input_83;
      end
      10'b0001010100 : begin
        result = input_84;
      end
      10'b0001010101 : begin
        result = input_85;
      end
      10'b0001010110 : begin
        result = input_86;
      end
      10'b0001010111 : begin
        result = input_87;
      end
      10'b0001011000 : begin
        result = input_88;
      end
      10'b0001011001 : begin
        result = input_89;
      end
      10'b0001011010 : begin
        result = input_90;
      end
      10'b0001011011 : begin
        result = input_91;
      end
      10'b0001011100 : begin
        result = input_92;
      end
      10'b0001011101 : begin
        result = input_93;
      end
      10'b0001011110 : begin
        result = input_94;
      end
      10'b0001011111 : begin
        result = input_95;
      end
      10'b0001100000 : begin
        result = input_96;
      end
      10'b0001100001 : begin
        result = input_97;
      end
      10'b0001100010 : begin
        result = input_98;
      end
      10'b0001100011 : begin
        result = input_99;
      end
      10'b0001100100 : begin
        result = input_100;
      end
      10'b0001100101 : begin
        result = input_101;
      end
      10'b0001100110 : begin
        result = input_102;
      end
      10'b0001100111 : begin
        result = input_103;
      end
      10'b0001101000 : begin
        result = input_104;
      end
      10'b0001101001 : begin
        result = input_105;
      end
      10'b0001101010 : begin
        result = input_106;
      end
      10'b0001101011 : begin
        result = input_107;
      end
      10'b0001101100 : begin
        result = input_108;
      end
      10'b0001101101 : begin
        result = input_109;
      end
      10'b0001101110 : begin
        result = input_110;
      end
      10'b0001101111 : begin
        result = input_111;
      end
      10'b0001110000 : begin
        result = input_112;
      end
      10'b0001110001 : begin
        result = input_113;
      end
      10'b0001110010 : begin
        result = input_114;
      end
      10'b0001110011 : begin
        result = input_115;
      end
      10'b0001110100 : begin
        result = input_116;
      end
      10'b0001110101 : begin
        result = input_117;
      end
      10'b0001110110 : begin
        result = input_118;
      end
      10'b0001110111 : begin
        result = input_119;
      end
      10'b0001111000 : begin
        result = input_120;
      end
      10'b0001111001 : begin
        result = input_121;
      end
      10'b0001111010 : begin
        result = input_122;
      end
      10'b0001111011 : begin
        result = input_123;
      end
      10'b0001111100 : begin
        result = input_124;
      end
      10'b0001111101 : begin
        result = input_125;
      end
      10'b0001111110 : begin
        result = input_126;
      end
      10'b0001111111 : begin
        result = input_127;
      end
      10'b0010000000 : begin
        result = input_128;
      end
      10'b0010000001 : begin
        result = input_129;
      end
      10'b0010000010 : begin
        result = input_130;
      end
      10'b0010000011 : begin
        result = input_131;
      end
      10'b0010000100 : begin
        result = input_132;
      end
      10'b0010000101 : begin
        result = input_133;
      end
      10'b0010000110 : begin
        result = input_134;
      end
      10'b0010000111 : begin
        result = input_135;
      end
      10'b0010001000 : begin
        result = input_136;
      end
      10'b0010001001 : begin
        result = input_137;
      end
      10'b0010001010 : begin
        result = input_138;
      end
      10'b0010001011 : begin
        result = input_139;
      end
      10'b0010001100 : begin
        result = input_140;
      end
      10'b0010001101 : begin
        result = input_141;
      end
      10'b0010001110 : begin
        result = input_142;
      end
      10'b0010001111 : begin
        result = input_143;
      end
      10'b0010010000 : begin
        result = input_144;
      end
      10'b0010010001 : begin
        result = input_145;
      end
      10'b0010010010 : begin
        result = input_146;
      end
      10'b0010010011 : begin
        result = input_147;
      end
      10'b0010010100 : begin
        result = input_148;
      end
      10'b0010010101 : begin
        result = input_149;
      end
      10'b0010010110 : begin
        result = input_150;
      end
      10'b0010010111 : begin
        result = input_151;
      end
      10'b0010011000 : begin
        result = input_152;
      end
      10'b0010011001 : begin
        result = input_153;
      end
      10'b0010011010 : begin
        result = input_154;
      end
      10'b0010011011 : begin
        result = input_155;
      end
      10'b0010011100 : begin
        result = input_156;
      end
      10'b0010011101 : begin
        result = input_157;
      end
      10'b0010011110 : begin
        result = input_158;
      end
      10'b0010011111 : begin
        result = input_159;
      end
      10'b0010100000 : begin
        result = input_160;
      end
      10'b0010100001 : begin
        result = input_161;
      end
      10'b0010100010 : begin
        result = input_162;
      end
      10'b0010100011 : begin
        result = input_163;
      end
      10'b0010100100 : begin
        result = input_164;
      end
      10'b0010100101 : begin
        result = input_165;
      end
      10'b0010100110 : begin
        result = input_166;
      end
      10'b0010100111 : begin
        result = input_167;
      end
      10'b0010101000 : begin
        result = input_168;
      end
      10'b0010101001 : begin
        result = input_169;
      end
      10'b0010101010 : begin
        result = input_170;
      end
      10'b0010101011 : begin
        result = input_171;
      end
      10'b0010101100 : begin
        result = input_172;
      end
      10'b0010101101 : begin
        result = input_173;
      end
      10'b0010101110 : begin
        result = input_174;
      end
      10'b0010101111 : begin
        result = input_175;
      end
      10'b0010110000 : begin
        result = input_176;
      end
      10'b0010110001 : begin
        result = input_177;
      end
      10'b0010110010 : begin
        result = input_178;
      end
      10'b0010110011 : begin
        result = input_179;
      end
      10'b0010110100 : begin
        result = input_180;
      end
      10'b0010110101 : begin
        result = input_181;
      end
      10'b0010110110 : begin
        result = input_182;
      end
      10'b0010110111 : begin
        result = input_183;
      end
      10'b0010111000 : begin
        result = input_184;
      end
      10'b0010111001 : begin
        result = input_185;
      end
      10'b0010111010 : begin
        result = input_186;
      end
      10'b0010111011 : begin
        result = input_187;
      end
      10'b0010111100 : begin
        result = input_188;
      end
      10'b0010111101 : begin
        result = input_189;
      end
      10'b0010111110 : begin
        result = input_190;
      end
      10'b0010111111 : begin
        result = input_191;
      end
      10'b0011000000 : begin
        result = input_192;
      end
      10'b0011000001 : begin
        result = input_193;
      end
      10'b0011000010 : begin
        result = input_194;
      end
      10'b0011000011 : begin
        result = input_195;
      end
      10'b0011000100 : begin
        result = input_196;
      end
      10'b0011000101 : begin
        result = input_197;
      end
      10'b0011000110 : begin
        result = input_198;
      end
      10'b0011000111 : begin
        result = input_199;
      end
      10'b0011001000 : begin
        result = input_200;
      end
      10'b0011001001 : begin
        result = input_201;
      end
      10'b0011001010 : begin
        result = input_202;
      end
      10'b0011001011 : begin
        result = input_203;
      end
      10'b0011001100 : begin
        result = input_204;
      end
      10'b0011001101 : begin
        result = input_205;
      end
      10'b0011001110 : begin
        result = input_206;
      end
      10'b0011001111 : begin
        result = input_207;
      end
      10'b0011010000 : begin
        result = input_208;
      end
      10'b0011010001 : begin
        result = input_209;
      end
      10'b0011010010 : begin
        result = input_210;
      end
      10'b0011010011 : begin
        result = input_211;
      end
      10'b0011010100 : begin
        result = input_212;
      end
      10'b0011010101 : begin
        result = input_213;
      end
      10'b0011010110 : begin
        result = input_214;
      end
      10'b0011010111 : begin
        result = input_215;
      end
      10'b0011011000 : begin
        result = input_216;
      end
      10'b0011011001 : begin
        result = input_217;
      end
      10'b0011011010 : begin
        result = input_218;
      end
      10'b0011011011 : begin
        result = input_219;
      end
      10'b0011011100 : begin
        result = input_220;
      end
      10'b0011011101 : begin
        result = input_221;
      end
      10'b0011011110 : begin
        result = input_222;
      end
      10'b0011011111 : begin
        result = input_223;
      end
      10'b0011100000 : begin
        result = input_224;
      end
      10'b0011100001 : begin
        result = input_225;
      end
      10'b0011100010 : begin
        result = input_226;
      end
      10'b0011100011 : begin
        result = input_227;
      end
      10'b0011100100 : begin
        result = input_228;
      end
      10'b0011100101 : begin
        result = input_229;
      end
      10'b0011100110 : begin
        result = input_230;
      end
      10'b0011100111 : begin
        result = input_231;
      end
      10'b0011101000 : begin
        result = input_232;
      end
      10'b0011101001 : begin
        result = input_233;
      end
      10'b0011101010 : begin
        result = input_234;
      end
      10'b0011101011 : begin
        result = input_235;
      end
      10'b0011101100 : begin
        result = input_236;
      end
      10'b0011101101 : begin
        result = input_237;
      end
      10'b0011101110 : begin
        result = input_238;
      end
      10'b0011101111 : begin
        result = input_239;
      end
      10'b0011110000 : begin
        result = input_240;
      end
      10'b0011110001 : begin
        result = input_241;
      end
      10'b0011110010 : begin
        result = input_242;
      end
      10'b0011110011 : begin
        result = input_243;
      end
      10'b0011110100 : begin
        result = input_244;
      end
      10'b0011110101 : begin
        result = input_245;
      end
      10'b0011110110 : begin
        result = input_246;
      end
      10'b0011110111 : begin
        result = input_247;
      end
      10'b0011111000 : begin
        result = input_248;
      end
      10'b0011111001 : begin
        result = input_249;
      end
      10'b0011111010 : begin
        result = input_250;
      end
      10'b0011111011 : begin
        result = input_251;
      end
      10'b0011111100 : begin
        result = input_252;
      end
      10'b0011111101 : begin
        result = input_253;
      end
      10'b0011111110 : begin
        result = input_254;
      end
      10'b0011111111 : begin
        result = input_255;
      end
      10'b0100000000 : begin
        result = input_256;
      end
      10'b0100000001 : begin
        result = input_257;
      end
      10'b0100000010 : begin
        result = input_258;
      end
      10'b0100000011 : begin
        result = input_259;
      end
      10'b0100000100 : begin
        result = input_260;
      end
      10'b0100000101 : begin
        result = input_261;
      end
      10'b0100000110 : begin
        result = input_262;
      end
      10'b0100000111 : begin
        result = input_263;
      end
      10'b0100001000 : begin
        result = input_264;
      end
      10'b0100001001 : begin
        result = input_265;
      end
      10'b0100001010 : begin
        result = input_266;
      end
      10'b0100001011 : begin
        result = input_267;
      end
      10'b0100001100 : begin
        result = input_268;
      end
      10'b0100001101 : begin
        result = input_269;
      end
      10'b0100001110 : begin
        result = input_270;
      end
      10'b0100001111 : begin
        result = input_271;
      end
      10'b0100010000 : begin
        result = input_272;
      end
      10'b0100010001 : begin
        result = input_273;
      end
      10'b0100010010 : begin
        result = input_274;
      end
      10'b0100010011 : begin
        result = input_275;
      end
      10'b0100010100 : begin
        result = input_276;
      end
      10'b0100010101 : begin
        result = input_277;
      end
      10'b0100010110 : begin
        result = input_278;
      end
      10'b0100010111 : begin
        result = input_279;
      end
      10'b0100011000 : begin
        result = input_280;
      end
      10'b0100011001 : begin
        result = input_281;
      end
      10'b0100011010 : begin
        result = input_282;
      end
      10'b0100011011 : begin
        result = input_283;
      end
      10'b0100011100 : begin
        result = input_284;
      end
      10'b0100011101 : begin
        result = input_285;
      end
      10'b0100011110 : begin
        result = input_286;
      end
      10'b0100011111 : begin
        result = input_287;
      end
      10'b0100100000 : begin
        result = input_288;
      end
      10'b0100100001 : begin
        result = input_289;
      end
      10'b0100100010 : begin
        result = input_290;
      end
      10'b0100100011 : begin
        result = input_291;
      end
      10'b0100100100 : begin
        result = input_292;
      end
      10'b0100100101 : begin
        result = input_293;
      end
      10'b0100100110 : begin
        result = input_294;
      end
      10'b0100100111 : begin
        result = input_295;
      end
      10'b0100101000 : begin
        result = input_296;
      end
      10'b0100101001 : begin
        result = input_297;
      end
      10'b0100101010 : begin
        result = input_298;
      end
      10'b0100101011 : begin
        result = input_299;
      end
      10'b0100101100 : begin
        result = input_300;
      end
      10'b0100101101 : begin
        result = input_301;
      end
      10'b0100101110 : begin
        result = input_302;
      end
      10'b0100101111 : begin
        result = input_303;
      end
      10'b0100110000 : begin
        result = input_304;
      end
      10'b0100110001 : begin
        result = input_305;
      end
      10'b0100110010 : begin
        result = input_306;
      end
      10'b0100110011 : begin
        result = input_307;
      end
      10'b0100110100 : begin
        result = input_308;
      end
      10'b0100110101 : begin
        result = input_309;
      end
      10'b0100110110 : begin
        result = input_310;
      end
      10'b0100110111 : begin
        result = input_311;
      end
      10'b0100111000 : begin
        result = input_312;
      end
      10'b0100111001 : begin
        result = input_313;
      end
      10'b0100111010 : begin
        result = input_314;
      end
      10'b0100111011 : begin
        result = input_315;
      end
      10'b0100111100 : begin
        result = input_316;
      end
      10'b0100111101 : begin
        result = input_317;
      end
      10'b0100111110 : begin
        result = input_318;
      end
      10'b0100111111 : begin
        result = input_319;
      end
      10'b0101000000 : begin
        result = input_320;
      end
      10'b0101000001 : begin
        result = input_321;
      end
      10'b0101000010 : begin
        result = input_322;
      end
      10'b0101000011 : begin
        result = input_323;
      end
      10'b0101000100 : begin
        result = input_324;
      end
      10'b0101000101 : begin
        result = input_325;
      end
      10'b0101000110 : begin
        result = input_326;
      end
      10'b0101000111 : begin
        result = input_327;
      end
      10'b0101001000 : begin
        result = input_328;
      end
      10'b0101001001 : begin
        result = input_329;
      end
      10'b0101001010 : begin
        result = input_330;
      end
      10'b0101001011 : begin
        result = input_331;
      end
      10'b0101001100 : begin
        result = input_332;
      end
      10'b0101001101 : begin
        result = input_333;
      end
      10'b0101001110 : begin
        result = input_334;
      end
      10'b0101001111 : begin
        result = input_335;
      end
      10'b0101010000 : begin
        result = input_336;
      end
      10'b0101010001 : begin
        result = input_337;
      end
      10'b0101010010 : begin
        result = input_338;
      end
      10'b0101010011 : begin
        result = input_339;
      end
      10'b0101010100 : begin
        result = input_340;
      end
      10'b0101010101 : begin
        result = input_341;
      end
      10'b0101010110 : begin
        result = input_342;
      end
      10'b0101010111 : begin
        result = input_343;
      end
      10'b0101011000 : begin
        result = input_344;
      end
      10'b0101011001 : begin
        result = input_345;
      end
      10'b0101011010 : begin
        result = input_346;
      end
      10'b0101011011 : begin
        result = input_347;
      end
      10'b0101011100 : begin
        result = input_348;
      end
      10'b0101011101 : begin
        result = input_349;
      end
      10'b0101011110 : begin
        result = input_350;
      end
      10'b0101011111 : begin
        result = input_351;
      end
      10'b0101100000 : begin
        result = input_352;
      end
      10'b0101100001 : begin
        result = input_353;
      end
      10'b0101100010 : begin
        result = input_354;
      end
      10'b0101100011 : begin
        result = input_355;
      end
      10'b0101100100 : begin
        result = input_356;
      end
      10'b0101100101 : begin
        result = input_357;
      end
      10'b0101100110 : begin
        result = input_358;
      end
      10'b0101100111 : begin
        result = input_359;
      end
      10'b0101101000 : begin
        result = input_360;
      end
      10'b0101101001 : begin
        result = input_361;
      end
      10'b0101101010 : begin
        result = input_362;
      end
      10'b0101101011 : begin
        result = input_363;
      end
      10'b0101101100 : begin
        result = input_364;
      end
      10'b0101101101 : begin
        result = input_365;
      end
      10'b0101101110 : begin
        result = input_366;
      end
      10'b0101101111 : begin
        result = input_367;
      end
      10'b0101110000 : begin
        result = input_368;
      end
      10'b0101110001 : begin
        result = input_369;
      end
      10'b0101110010 : begin
        result = input_370;
      end
      10'b0101110011 : begin
        result = input_371;
      end
      10'b0101110100 : begin
        result = input_372;
      end
      10'b0101110101 : begin
        result = input_373;
      end
      10'b0101110110 : begin
        result = input_374;
      end
      10'b0101110111 : begin
        result = input_375;
      end
      10'b0101111000 : begin
        result = input_376;
      end
      10'b0101111001 : begin
        result = input_377;
      end
      10'b0101111010 : begin
        result = input_378;
      end
      10'b0101111011 : begin
        result = input_379;
      end
      10'b0101111100 : begin
        result = input_380;
      end
      10'b0101111101 : begin
        result = input_381;
      end
      10'b0101111110 : begin
        result = input_382;
      end
      10'b0101111111 : begin
        result = input_383;
      end
      10'b0110000000 : begin
        result = input_384;
      end
      10'b0110000001 : begin
        result = input_385;
      end
      10'b0110000010 : begin
        result = input_386;
      end
      10'b0110000011 : begin
        result = input_387;
      end
      10'b0110000100 : begin
        result = input_388;
      end
      10'b0110000101 : begin
        result = input_389;
      end
      10'b0110000110 : begin
        result = input_390;
      end
      10'b0110000111 : begin
        result = input_391;
      end
      10'b0110001000 : begin
        result = input_392;
      end
      10'b0110001001 : begin
        result = input_393;
      end
      10'b0110001010 : begin
        result = input_394;
      end
      10'b0110001011 : begin
        result = input_395;
      end
      10'b0110001100 : begin
        result = input_396;
      end
      10'b0110001101 : begin
        result = input_397;
      end
      10'b0110001110 : begin
        result = input_398;
      end
      10'b0110001111 : begin
        result = input_399;
      end
      10'b0110010000 : begin
        result = input_400;
      end
      10'b0110010001 : begin
        result = input_401;
      end
      10'b0110010010 : begin
        result = input_402;
      end
      10'b0110010011 : begin
        result = input_403;
      end
      10'b0110010100 : begin
        result = input_404;
      end
      10'b0110010101 : begin
        result = input_405;
      end
      10'b0110010110 : begin
        result = input_406;
      end
      10'b0110010111 : begin
        result = input_407;
      end
      10'b0110011000 : begin
        result = input_408;
      end
      10'b0110011001 : begin
        result = input_409;
      end
      10'b0110011010 : begin
        result = input_410;
      end
      10'b0110011011 : begin
        result = input_411;
      end
      10'b0110011100 : begin
        result = input_412;
      end
      10'b0110011101 : begin
        result = input_413;
      end
      10'b0110011110 : begin
        result = input_414;
      end
      10'b0110011111 : begin
        result = input_415;
      end
      10'b0110100000 : begin
        result = input_416;
      end
      10'b0110100001 : begin
        result = input_417;
      end
      10'b0110100010 : begin
        result = input_418;
      end
      10'b0110100011 : begin
        result = input_419;
      end
      10'b0110100100 : begin
        result = input_420;
      end
      10'b0110100101 : begin
        result = input_421;
      end
      10'b0110100110 : begin
        result = input_422;
      end
      10'b0110100111 : begin
        result = input_423;
      end
      10'b0110101000 : begin
        result = input_424;
      end
      10'b0110101001 : begin
        result = input_425;
      end
      10'b0110101010 : begin
        result = input_426;
      end
      10'b0110101011 : begin
        result = input_427;
      end
      10'b0110101100 : begin
        result = input_428;
      end
      10'b0110101101 : begin
        result = input_429;
      end
      10'b0110101110 : begin
        result = input_430;
      end
      10'b0110101111 : begin
        result = input_431;
      end
      10'b0110110000 : begin
        result = input_432;
      end
      10'b0110110001 : begin
        result = input_433;
      end
      10'b0110110010 : begin
        result = input_434;
      end
      10'b0110110011 : begin
        result = input_435;
      end
      10'b0110110100 : begin
        result = input_436;
      end
      10'b0110110101 : begin
        result = input_437;
      end
      10'b0110110110 : begin
        result = input_438;
      end
      10'b0110110111 : begin
        result = input_439;
      end
      10'b0110111000 : begin
        result = input_440;
      end
      10'b0110111001 : begin
        result = input_441;
      end
      10'b0110111010 : begin
        result = input_442;
      end
      10'b0110111011 : begin
        result = input_443;
      end
      10'b0110111100 : begin
        result = input_444;
      end
      10'b0110111101 : begin
        result = input_445;
      end
      10'b0110111110 : begin
        result = input_446;
      end
      10'b0110111111 : begin
        result = input_447;
      end
      10'b0111000000 : begin
        result = input_448;
      end
      10'b0111000001 : begin
        result = input_449;
      end
      10'b0111000010 : begin
        result = input_450;
      end
      10'b0111000011 : begin
        result = input_451;
      end
      10'b0111000100 : begin
        result = input_452;
      end
      10'b0111000101 : begin
        result = input_453;
      end
      10'b0111000110 : begin
        result = input_454;
      end
      10'b0111000111 : begin
        result = input_455;
      end
      10'b0111001000 : begin
        result = input_456;
      end
      10'b0111001001 : begin
        result = input_457;
      end
      10'b0111001010 : begin
        result = input_458;
      end
      10'b0111001011 : begin
        result = input_459;
      end
      10'b0111001100 : begin
        result = input_460;
      end
      10'b0111001101 : begin
        result = input_461;
      end
      10'b0111001110 : begin
        result = input_462;
      end
      10'b0111001111 : begin
        result = input_463;
      end
      10'b0111010000 : begin
        result = input_464;
      end
      10'b0111010001 : begin
        result = input_465;
      end
      10'b0111010010 : begin
        result = input_466;
      end
      10'b0111010011 : begin
        result = input_467;
      end
      10'b0111010100 : begin
        result = input_468;
      end
      10'b0111010101 : begin
        result = input_469;
      end
      10'b0111010110 : begin
        result = input_470;
      end
      10'b0111010111 : begin
        result = input_471;
      end
      10'b0111011000 : begin
        result = input_472;
      end
      10'b0111011001 : begin
        result = input_473;
      end
      10'b0111011010 : begin
        result = input_474;
      end
      10'b0111011011 : begin
        result = input_475;
      end
      10'b0111011100 : begin
        result = input_476;
      end
      10'b0111011101 : begin
        result = input_477;
      end
      10'b0111011110 : begin
        result = input_478;
      end
      10'b0111011111 : begin
        result = input_479;
      end
      10'b0111100000 : begin
        result = input_480;
      end
      10'b0111100001 : begin
        result = input_481;
      end
      10'b0111100010 : begin
        result = input_482;
      end
      10'b0111100011 : begin
        result = input_483;
      end
      10'b0111100100 : begin
        result = input_484;
      end
      10'b0111100101 : begin
        result = input_485;
      end
      10'b0111100110 : begin
        result = input_486;
      end
      10'b0111100111 : begin
        result = input_487;
      end
      10'b0111101000 : begin
        result = input_488;
      end
      10'b0111101001 : begin
        result = input_489;
      end
      10'b0111101010 : begin
        result = input_490;
      end
      10'b0111101011 : begin
        result = input_491;
      end
      10'b0111101100 : begin
        result = input_492;
      end
      10'b0111101101 : begin
        result = input_493;
      end
      10'b0111101110 : begin
        result = input_494;
      end
      10'b0111101111 : begin
        result = input_495;
      end
      10'b0111110000 : begin
        result = input_496;
      end
      10'b0111110001 : begin
        result = input_497;
      end
      10'b0111110010 : begin
        result = input_498;
      end
      10'b0111110011 : begin
        result = input_499;
      end
      10'b0111110100 : begin
        result = input_500;
      end
      10'b0111110101 : begin
        result = input_501;
      end
      10'b0111110110 : begin
        result = input_502;
      end
      10'b0111110111 : begin
        result = input_503;
      end
      10'b0111111000 : begin
        result = input_504;
      end
      10'b0111111001 : begin
        result = input_505;
      end
      10'b0111111010 : begin
        result = input_506;
      end
      10'b0111111011 : begin
        result = input_507;
      end
      10'b0111111100 : begin
        result = input_508;
      end
      10'b0111111101 : begin
        result = input_509;
      end
      10'b0111111110 : begin
        result = input_510;
      end
      10'b0111111111 : begin
        result = input_511;
      end
      10'b1000000000 : begin
        result = input_512;
      end
      10'b1000000001 : begin
        result = input_513;
      end
      10'b1000000010 : begin
        result = input_514;
      end
      10'b1000000011 : begin
        result = input_515;
      end
      10'b1000000100 : begin
        result = input_516;
      end
      10'b1000000101 : begin
        result = input_517;
      end
      10'b1000000110 : begin
        result = input_518;
      end
      10'b1000000111 : begin
        result = input_519;
      end
      10'b1000001000 : begin
        result = input_520;
      end
      10'b1000001001 : begin
        result = input_521;
      end
      10'b1000001010 : begin
        result = input_522;
      end
      10'b1000001011 : begin
        result = input_523;
      end
      10'b1000001100 : begin
        result = input_524;
      end
      10'b1000001101 : begin
        result = input_525;
      end
      10'b1000001110 : begin
        result = input_526;
      end
      10'b1000001111 : begin
        result = input_527;
      end
      10'b1000010000 : begin
        result = input_528;
      end
      10'b1000010001 : begin
        result = input_529;
      end
      10'b1000010010 : begin
        result = input_530;
      end
      10'b1000010011 : begin
        result = input_531;
      end
      10'b1000010100 : begin
        result = input_532;
      end
      10'b1000010101 : begin
        result = input_533;
      end
      10'b1000010110 : begin
        result = input_534;
      end
      10'b1000010111 : begin
        result = input_535;
      end
      10'b1000011000 : begin
        result = input_536;
      end
      10'b1000011001 : begin
        result = input_537;
      end
      10'b1000011010 : begin
        result = input_538;
      end
      10'b1000011011 : begin
        result = input_539;
      end
      10'b1000011100 : begin
        result = input_540;
      end
      10'b1000011101 : begin
        result = input_541;
      end
      10'b1000011110 : begin
        result = input_542;
      end
      10'b1000011111 : begin
        result = input_543;
      end
      10'b1000100000 : begin
        result = input_544;
      end
      10'b1000100001 : begin
        result = input_545;
      end
      10'b1000100010 : begin
        result = input_546;
      end
      10'b1000100011 : begin
        result = input_547;
      end
      10'b1000100100 : begin
        result = input_548;
      end
      10'b1000100101 : begin
        result = input_549;
      end
      10'b1000100110 : begin
        result = input_550;
      end
      10'b1000100111 : begin
        result = input_551;
      end
      10'b1000101000 : begin
        result = input_552;
      end
      10'b1000101001 : begin
        result = input_553;
      end
      10'b1000101010 : begin
        result = input_554;
      end
      10'b1000101011 : begin
        result = input_555;
      end
      10'b1000101100 : begin
        result = input_556;
      end
      10'b1000101101 : begin
        result = input_557;
      end
      10'b1000101110 : begin
        result = input_558;
      end
      10'b1000101111 : begin
        result = input_559;
      end
      10'b1000110000 : begin
        result = input_560;
      end
      10'b1000110001 : begin
        result = input_561;
      end
      10'b1000110010 : begin
        result = input_562;
      end
      10'b1000110011 : begin
        result = input_563;
      end
      10'b1000110100 : begin
        result = input_564;
      end
      10'b1000110101 : begin
        result = input_565;
      end
      10'b1000110110 : begin
        result = input_566;
      end
      10'b1000110111 : begin
        result = input_567;
      end
      10'b1000111000 : begin
        result = input_568;
      end
      10'b1000111001 : begin
        result = input_569;
      end
      10'b1000111010 : begin
        result = input_570;
      end
      10'b1000111011 : begin
        result = input_571;
      end
      10'b1000111100 : begin
        result = input_572;
      end
      10'b1000111101 : begin
        result = input_573;
      end
      10'b1000111110 : begin
        result = input_574;
      end
      10'b1000111111 : begin
        result = input_575;
      end
      10'b1001000000 : begin
        result = input_576;
      end
      10'b1001000001 : begin
        result = input_577;
      end
      10'b1001000010 : begin
        result = input_578;
      end
      10'b1001000011 : begin
        result = input_579;
      end
      10'b1001000100 : begin
        result = input_580;
      end
      10'b1001000101 : begin
        result = input_581;
      end
      10'b1001000110 : begin
        result = input_582;
      end
      10'b1001000111 : begin
        result = input_583;
      end
      10'b1001001000 : begin
        result = input_584;
      end
      10'b1001001001 : begin
        result = input_585;
      end
      10'b1001001010 : begin
        result = input_586;
      end
      10'b1001001011 : begin
        result = input_587;
      end
      10'b1001001100 : begin
        result = input_588;
      end
      10'b1001001101 : begin
        result = input_589;
      end
      10'b1001001110 : begin
        result = input_590;
      end
      10'b1001001111 : begin
        result = input_591;
      end
      10'b1001010000 : begin
        result = input_592;
      end
      10'b1001010001 : begin
        result = input_593;
      end
      10'b1001010010 : begin
        result = input_594;
      end
      10'b1001010011 : begin
        result = input_595;
      end
      10'b1001010100 : begin
        result = input_596;
      end
      10'b1001010101 : begin
        result = input_597;
      end
      10'b1001010110 : begin
        result = input_598;
      end
      10'b1001010111 : begin
        result = input_599;
      end
      10'b1001011000 : begin
        result = input_600;
      end
      10'b1001011001 : begin
        result = input_601;
      end
      10'b1001011010 : begin
        result = input_602;
      end
      10'b1001011011 : begin
        result = input_603;
      end
      10'b1001011100 : begin
        result = input_604;
      end
      10'b1001011101 : begin
        result = input_605;
      end
      10'b1001011110 : begin
        result = input_606;
      end
      10'b1001011111 : begin
        result = input_607;
      end
      10'b1001100000 : begin
        result = input_608;
      end
      10'b1001100001 : begin
        result = input_609;
      end
      10'b1001100010 : begin
        result = input_610;
      end
      10'b1001100011 : begin
        result = input_611;
      end
      10'b1001100100 : begin
        result = input_612;
      end
      10'b1001100101 : begin
        result = input_613;
      end
      10'b1001100110 : begin
        result = input_614;
      end
      10'b1001100111 : begin
        result = input_615;
      end
      10'b1001101000 : begin
        result = input_616;
      end
      10'b1001101001 : begin
        result = input_617;
      end
      10'b1001101010 : begin
        result = input_618;
      end
      10'b1001101011 : begin
        result = input_619;
      end
      10'b1001101100 : begin
        result = input_620;
      end
      10'b1001101101 : begin
        result = input_621;
      end
      10'b1001101110 : begin
        result = input_622;
      end
      10'b1001101111 : begin
        result = input_623;
      end
      10'b1001110000 : begin
        result = input_624;
      end
      10'b1001110001 : begin
        result = input_625;
      end
      10'b1001110010 : begin
        result = input_626;
      end
      10'b1001110011 : begin
        result = input_627;
      end
      10'b1001110100 : begin
        result = input_628;
      end
      10'b1001110101 : begin
        result = input_629;
      end
      10'b1001110110 : begin
        result = input_630;
      end
      10'b1001110111 : begin
        result = input_631;
      end
      10'b1001111000 : begin
        result = input_632;
      end
      10'b1001111001 : begin
        result = input_633;
      end
      10'b1001111010 : begin
        result = input_634;
      end
      10'b1001111011 : begin
        result = input_635;
      end
      10'b1001111100 : begin
        result = input_636;
      end
      10'b1001111101 : begin
        result = input_637;
      end
      10'b1001111110 : begin
        result = input_638;
      end
      10'b1001111111 : begin
        result = input_639;
      end
      10'b1010000000 : begin
        result = input_640;
      end
      10'b1010000001 : begin
        result = input_641;
      end
      10'b1010000010 : begin
        result = input_642;
      end
      10'b1010000011 : begin
        result = input_643;
      end
      10'b1010000100 : begin
        result = input_644;
      end
      10'b1010000101 : begin
        result = input_645;
      end
      10'b1010000110 : begin
        result = input_646;
      end
      10'b1010000111 : begin
        result = input_647;
      end
      10'b1010001000 : begin
        result = input_648;
      end
      10'b1010001001 : begin
        result = input_649;
      end
      10'b1010001010 : begin
        result = input_650;
      end
      10'b1010001011 : begin
        result = input_651;
      end
      10'b1010001100 : begin
        result = input_652;
      end
      10'b1010001101 : begin
        result = input_653;
      end
      10'b1010001110 : begin
        result = input_654;
      end
      10'b1010001111 : begin
        result = input_655;
      end
      10'b1010010000 : begin
        result = input_656;
      end
      10'b1010010001 : begin
        result = input_657;
      end
      10'b1010010010 : begin
        result = input_658;
      end
      10'b1010010011 : begin
        result = input_659;
      end
      10'b1010010100 : begin
        result = input_660;
      end
      10'b1010010101 : begin
        result = input_661;
      end
      10'b1010010110 : begin
        result = input_662;
      end
      10'b1010010111 : begin
        result = input_663;
      end
      10'b1010011000 : begin
        result = input_664;
      end
      10'b1010011001 : begin
        result = input_665;
      end
      10'b1010011010 : begin
        result = input_666;
      end
      10'b1010011011 : begin
        result = input_667;
      end
      10'b1010011100 : begin
        result = input_668;
      end
      10'b1010011101 : begin
        result = input_669;
      end
      10'b1010011110 : begin
        result = input_670;
      end
      10'b1010011111 : begin
        result = input_671;
      end
      10'b1010100000 : begin
        result = input_672;
      end
      10'b1010100001 : begin
        result = input_673;
      end
      10'b1010100010 : begin
        result = input_674;
      end
      10'b1010100011 : begin
        result = input_675;
      end
      10'b1010100100 : begin
        result = input_676;
      end
      10'b1010100101 : begin
        result = input_677;
      end
      10'b1010100110 : begin
        result = input_678;
      end
      10'b1010100111 : begin
        result = input_679;
      end
      10'b1010101000 : begin
        result = input_680;
      end
      10'b1010101001 : begin
        result = input_681;
      end
      10'b1010101010 : begin
        result = input_682;
      end
      10'b1010101011 : begin
        result = input_683;
      end
      10'b1010101100 : begin
        result = input_684;
      end
      10'b1010101101 : begin
        result = input_685;
      end
      10'b1010101110 : begin
        result = input_686;
      end
      10'b1010101111 : begin
        result = input_687;
      end
      10'b1010110000 : begin
        result = input_688;
      end
      10'b1010110001 : begin
        result = input_689;
      end
      10'b1010110010 : begin
        result = input_690;
      end
      10'b1010110011 : begin
        result = input_691;
      end
      10'b1010110100 : begin
        result = input_692;
      end
      10'b1010110101 : begin
        result = input_693;
      end
      10'b1010110110 : begin
        result = input_694;
      end
      10'b1010110111 : begin
        result = input_695;
      end
      10'b1010111000 : begin
        result = input_696;
      end
      10'b1010111001 : begin
        result = input_697;
      end
      10'b1010111010 : begin
        result = input_698;
      end
      10'b1010111011 : begin
        result = input_699;
      end
      10'b1010111100 : begin
        result = input_700;
      end
      10'b1010111101 : begin
        result = input_701;
      end
      10'b1010111110 : begin
        result = input_702;
      end
      10'b1010111111 : begin
        result = input_703;
      end
      10'b1011000000 : begin
        result = input_704;
      end
      10'b1011000001 : begin
        result = input_705;
      end
      10'b1011000010 : begin
        result = input_706;
      end
      10'b1011000011 : begin
        result = input_707;
      end
      10'b1011000100 : begin
        result = input_708;
      end
      10'b1011000101 : begin
        result = input_709;
      end
      10'b1011000110 : begin
        result = input_710;
      end
      10'b1011000111 : begin
        result = input_711;
      end
      10'b1011001000 : begin
        result = input_712;
      end
      10'b1011001001 : begin
        result = input_713;
      end
      10'b1011001010 : begin
        result = input_714;
      end
      10'b1011001011 : begin
        result = input_715;
      end
      10'b1011001100 : begin
        result = input_716;
      end
      10'b1011001101 : begin
        result = input_717;
      end
      10'b1011001110 : begin
        result = input_718;
      end
      10'b1011001111 : begin
        result = input_719;
      end
      10'b1011010000 : begin
        result = input_720;
      end
      10'b1011010001 : begin
        result = input_721;
      end
      10'b1011010010 : begin
        result = input_722;
      end
      10'b1011010011 : begin
        result = input_723;
      end
      10'b1011010100 : begin
        result = input_724;
      end
      10'b1011010101 : begin
        result = input_725;
      end
      10'b1011010110 : begin
        result = input_726;
      end
      10'b1011010111 : begin
        result = input_727;
      end
      10'b1011011000 : begin
        result = input_728;
      end
      10'b1011011001 : begin
        result = input_729;
      end
      10'b1011011010 : begin
        result = input_730;
      end
      10'b1011011011 : begin
        result = input_731;
      end
      10'b1011011100 : begin
        result = input_732;
      end
      10'b1011011101 : begin
        result = input_733;
      end
      10'b1011011110 : begin
        result = input_734;
      end
      10'b1011011111 : begin
        result = input_735;
      end
      10'b1011100000 : begin
        result = input_736;
      end
      10'b1011100001 : begin
        result = input_737;
      end
      10'b1011100010 : begin
        result = input_738;
      end
      10'b1011100011 : begin
        result = input_739;
      end
      10'b1011100100 : begin
        result = input_740;
      end
      10'b1011100101 : begin
        result = input_741;
      end
      10'b1011100110 : begin
        result = input_742;
      end
      10'b1011100111 : begin
        result = input_743;
      end
      10'b1011101000 : begin
        result = input_744;
      end
      10'b1011101001 : begin
        result = input_745;
      end
      10'b1011101010 : begin
        result = input_746;
      end
      10'b1011101011 : begin
        result = input_747;
      end
      10'b1011101100 : begin
        result = input_748;
      end
      10'b1011101101 : begin
        result = input_749;
      end
      10'b1011101110 : begin
        result = input_750;
      end
      10'b1011101111 : begin
        result = input_751;
      end
      10'b1011110000 : begin
        result = input_752;
      end
      10'b1011110001 : begin
        result = input_753;
      end
      10'b1011110010 : begin
        result = input_754;
      end
      10'b1011110011 : begin
        result = input_755;
      end
      10'b1011110100 : begin
        result = input_756;
      end
      10'b1011110101 : begin
        result = input_757;
      end
      10'b1011110110 : begin
        result = input_758;
      end
      10'b1011110111 : begin
        result = input_759;
      end
      10'b1011111000 : begin
        result = input_760;
      end
      10'b1011111001 : begin
        result = input_761;
      end
      10'b1011111010 : begin
        result = input_762;
      end
      10'b1011111011 : begin
        result = input_763;
      end
      10'b1011111100 : begin
        result = input_764;
      end
      10'b1011111101 : begin
        result = input_765;
      end
      10'b1011111110 : begin
        result = input_766;
      end
      10'b1011111111 : begin
        result = input_767;
      end
      10'b1100000000 : begin
        result = input_768;
      end
      10'b1100000001 : begin
        result = input_769;
      end
      10'b1100000010 : begin
        result = input_770;
      end
      10'b1100000011 : begin
        result = input_771;
      end
      10'b1100000100 : begin
        result = input_772;
      end
      10'b1100000101 : begin
        result = input_773;
      end
      10'b1100000110 : begin
        result = input_774;
      end
      10'b1100000111 : begin
        result = input_775;
      end
      10'b1100001000 : begin
        result = input_776;
      end
      10'b1100001001 : begin
        result = input_777;
      end
      10'b1100001010 : begin
        result = input_778;
      end
      10'b1100001011 : begin
        result = input_779;
      end
      10'b1100001100 : begin
        result = input_780;
      end
      10'b1100001101 : begin
        result = input_781;
      end
      10'b1100001110 : begin
        result = input_782;
      end
      10'b1100001111 : begin
        result = input_783;
      end
      10'b1100010000 : begin
        result = input_784;
      end
      10'b1100010001 : begin
        result = input_785;
      end
      10'b1100010010 : begin
        result = input_786;
      end
      10'b1100010011 : begin
        result = input_787;
      end
      10'b1100010100 : begin
        result = input_788;
      end
      10'b1100010101 : begin
        result = input_789;
      end
      10'b1100010110 : begin
        result = input_790;
      end
      10'b1100010111 : begin
        result = input_791;
      end
      10'b1100011000 : begin
        result = input_792;
      end
      10'b1100011001 : begin
        result = input_793;
      end
      10'b1100011010 : begin
        result = input_794;
      end
      10'b1100011011 : begin
        result = input_795;
      end
      10'b1100011100 : begin
        result = input_796;
      end
      10'b1100011101 : begin
        result = input_797;
      end
      10'b1100011110 : begin
        result = input_798;
      end
      10'b1100011111 : begin
        result = input_799;
      end
      10'b1100100000 : begin
        result = input_800;
      end
      10'b1100100001 : begin
        result = input_801;
      end
      10'b1100100010 : begin
        result = input_802;
      end
      10'b1100100011 : begin
        result = input_803;
      end
      10'b1100100100 : begin
        result = input_804;
      end
      10'b1100100101 : begin
        result = input_805;
      end
      10'b1100100110 : begin
        result = input_806;
      end
      10'b1100100111 : begin
        result = input_807;
      end
      10'b1100101000 : begin
        result = input_808;
      end
      10'b1100101001 : begin
        result = input_809;
      end
      10'b1100101010 : begin
        result = input_810;
      end
      10'b1100101011 : begin
        result = input_811;
      end
      10'b1100101100 : begin
        result = input_812;
      end
      10'b1100101101 : begin
        result = input_813;
      end
      10'b1100101110 : begin
        result = input_814;
      end
      10'b1100101111 : begin
        result = input_815;
      end
      10'b1100110000 : begin
        result = input_816;
      end
      10'b1100110001 : begin
        result = input_817;
      end
      10'b1100110010 : begin
        result = input_818;
      end
      10'b1100110011 : begin
        result = input_819;
      end
      10'b1100110100 : begin
        result = input_820;
      end
      10'b1100110101 : begin
        result = input_821;
      end
      10'b1100110110 : begin
        result = input_822;
      end
      10'b1100110111 : begin
        result = input_823;
      end
      10'b1100111000 : begin
        result = input_824;
      end
      10'b1100111001 : begin
        result = input_825;
      end
      10'b1100111010 : begin
        result = input_826;
      end
      10'b1100111011 : begin
        result = input_827;
      end
      10'b1100111100 : begin
        result = input_828;
      end
      10'b1100111101 : begin
        result = input_829;
      end
      10'b1100111110 : begin
        result = input_830;
      end
      10'b1100111111 : begin
        result = input_831;
      end
      10'b1101000000 : begin
        result = input_832;
      end
      10'b1101000001 : begin
        result = input_833;
      end
      10'b1101000010 : begin
        result = input_834;
      end
      10'b1101000011 : begin
        result = input_835;
      end
      10'b1101000100 : begin
        result = input_836;
      end
      10'b1101000101 : begin
        result = input_837;
      end
      10'b1101000110 : begin
        result = input_838;
      end
      10'b1101000111 : begin
        result = input_839;
      end
      10'b1101001000 : begin
        result = input_840;
      end
      10'b1101001001 : begin
        result = input_841;
      end
      10'b1101001010 : begin
        result = input_842;
      end
      10'b1101001011 : begin
        result = input_843;
      end
      10'b1101001100 : begin
        result = input_844;
      end
      10'b1101001101 : begin
        result = input_845;
      end
      10'b1101001110 : begin
        result = input_846;
      end
      10'b1101001111 : begin
        result = input_847;
      end
      10'b1101010000 : begin
        result = input_848;
      end
      10'b1101010001 : begin
        result = input_849;
      end
      10'b1101010010 : begin
        result = input_850;
      end
      10'b1101010011 : begin
        result = input_851;
      end
      10'b1101010100 : begin
        result = input_852;
      end
      10'b1101010101 : begin
        result = input_853;
      end
      10'b1101010110 : begin
        result = input_854;
      end
      10'b1101010111 : begin
        result = input_855;
      end
      10'b1101011000 : begin
        result = input_856;
      end
      10'b1101011001 : begin
        result = input_857;
      end
      10'b1101011010 : begin
        result = input_858;
      end
      10'b1101011011 : begin
        result = input_859;
      end
      10'b1101011100 : begin
        result = input_860;
      end
      10'b1101011101 : begin
        result = input_861;
      end
      10'b1101011110 : begin
        result = input_862;
      end
      10'b1101011111 : begin
        result = input_863;
      end
      10'b1101100000 : begin
        result = input_864;
      end
      10'b1101100001 : begin
        result = input_865;
      end
      10'b1101100010 : begin
        result = input_866;
      end
      10'b1101100011 : begin
        result = input_867;
      end
      10'b1101100100 : begin
        result = input_868;
      end
      10'b1101100101 : begin
        result = input_869;
      end
      10'b1101100110 : begin
        result = input_870;
      end
      10'b1101100111 : begin
        result = input_871;
      end
      10'b1101101000 : begin
        result = input_872;
      end
      10'b1101101001 : begin
        result = input_873;
      end
      10'b1101101010 : begin
        result = input_874;
      end
      10'b1101101011 : begin
        result = input_875;
      end
      10'b1101101100 : begin
        result = input_876;
      end
      10'b1101101101 : begin
        result = input_877;
      end
      10'b1101101110 : begin
        result = input_878;
      end
      10'b1101101111 : begin
        result = input_879;
      end
      10'b1101110000 : begin
        result = input_880;
      end
      10'b1101110001 : begin
        result = input_881;
      end
      10'b1101110010 : begin
        result = input_882;
      end
      10'b1101110011 : begin
        result = input_883;
      end
      10'b1101110100 : begin
        result = input_884;
      end
      10'b1101110101 : begin
        result = input_885;
      end
      10'b1101110110 : begin
        result = input_886;
      end
      10'b1101110111 : begin
        result = input_887;
      end
      10'b1101111000 : begin
        result = input_888;
      end
      10'b1101111001 : begin
        result = input_889;
      end
      10'b1101111010 : begin
        result = input_890;
      end
      10'b1101111011 : begin
        result = input_891;
      end
      10'b1101111100 : begin
        result = input_892;
      end
      10'b1101111101 : begin
        result = input_893;
      end
      10'b1101111110 : begin
        result = input_894;
      end
      10'b1101111111 : begin
        result = input_895;
      end
      10'b1110000000 : begin
        result = input_896;
      end
      10'b1110000001 : begin
        result = input_897;
      end
      10'b1110000010 : begin
        result = input_898;
      end
      10'b1110000011 : begin
        result = input_899;
      end
      10'b1110000100 : begin
        result = input_900;
      end
      10'b1110000101 : begin
        result = input_901;
      end
      10'b1110000110 : begin
        result = input_902;
      end
      10'b1110000111 : begin
        result = input_903;
      end
      10'b1110001000 : begin
        result = input_904;
      end
      10'b1110001001 : begin
        result = input_905;
      end
      10'b1110001010 : begin
        result = input_906;
      end
      10'b1110001011 : begin
        result = input_907;
      end
      10'b1110001100 : begin
        result = input_908;
      end
      10'b1110001101 : begin
        result = input_909;
      end
      10'b1110001110 : begin
        result = input_910;
      end
      10'b1110001111 : begin
        result = input_911;
      end
      10'b1110010000 : begin
        result = input_912;
      end
      10'b1110010001 : begin
        result = input_913;
      end
      10'b1110010010 : begin
        result = input_914;
      end
      10'b1110010011 : begin
        result = input_915;
      end
      10'b1110010100 : begin
        result = input_916;
      end
      10'b1110010101 : begin
        result = input_917;
      end
      10'b1110010110 : begin
        result = input_918;
      end
      10'b1110010111 : begin
        result = input_919;
      end
      10'b1110011000 : begin
        result = input_920;
      end
      10'b1110011001 : begin
        result = input_921;
      end
      10'b1110011010 : begin
        result = input_922;
      end
      10'b1110011011 : begin
        result = input_923;
      end
      10'b1110011100 : begin
        result = input_924;
      end
      10'b1110011101 : begin
        result = input_925;
      end
      10'b1110011110 : begin
        result = input_926;
      end
      10'b1110011111 : begin
        result = input_927;
      end
      10'b1110100000 : begin
        result = input_928;
      end
      10'b1110100001 : begin
        result = input_929;
      end
      10'b1110100010 : begin
        result = input_930;
      end
      10'b1110100011 : begin
        result = input_931;
      end
      10'b1110100100 : begin
        result = input_932;
      end
      10'b1110100101 : begin
        result = input_933;
      end
      10'b1110100110 : begin
        result = input_934;
      end
      10'b1110100111 : begin
        result = input_935;
      end
      10'b1110101000 : begin
        result = input_936;
      end
      10'b1110101001 : begin
        result = input_937;
      end
      10'b1110101010 : begin
        result = input_938;
      end
      10'b1110101011 : begin
        result = input_939;
      end
      10'b1110101100 : begin
        result = input_940;
      end
      10'b1110101101 : begin
        result = input_941;
      end
      10'b1110101110 : begin
        result = input_942;
      end
      10'b1110101111 : begin
        result = input_943;
      end
      10'b1110110000 : begin
        result = input_944;
      end
      10'b1110110001 : begin
        result = input_945;
      end
      10'b1110110010 : begin
        result = input_946;
      end
      10'b1110110011 : begin
        result = input_947;
      end
      10'b1110110100 : begin
        result = input_948;
      end
      10'b1110110101 : begin
        result = input_949;
      end
      10'b1110110110 : begin
        result = input_950;
      end
      10'b1110110111 : begin
        result = input_951;
      end
      10'b1110111000 : begin
        result = input_952;
      end
      10'b1110111001 : begin
        result = input_953;
      end
      10'b1110111010 : begin
        result = input_954;
      end
      10'b1110111011 : begin
        result = input_955;
      end
      10'b1110111100 : begin
        result = input_956;
      end
      10'b1110111101 : begin
        result = input_957;
      end
      10'b1110111110 : begin
        result = input_958;
      end
      10'b1110111111 : begin
        result = input_959;
      end
      10'b1111000000 : begin
        result = input_960;
      end
      10'b1111000001 : begin
        result = input_961;
      end
      10'b1111000010 : begin
        result = input_962;
      end
      10'b1111000011 : begin
        result = input_963;
      end
      10'b1111000100 : begin
        result = input_964;
      end
      10'b1111000101 : begin
        result = input_965;
      end
      10'b1111000110 : begin
        result = input_966;
      end
      10'b1111000111 : begin
        result = input_967;
      end
      10'b1111001000 : begin
        result = input_968;
      end
      10'b1111001001 : begin
        result = input_969;
      end
      10'b1111001010 : begin
        result = input_970;
      end
      10'b1111001011 : begin
        result = input_971;
      end
      10'b1111001100 : begin
        result = input_972;
      end
      10'b1111001101 : begin
        result = input_973;
      end
      10'b1111001110 : begin
        result = input_974;
      end
      10'b1111001111 : begin
        result = input_975;
      end
      10'b1111010000 : begin
        result = input_976;
      end
      10'b1111010001 : begin
        result = input_977;
      end
      10'b1111010010 : begin
        result = input_978;
      end
      10'b1111010011 : begin
        result = input_979;
      end
      10'b1111010100 : begin
        result = input_980;
      end
      10'b1111010101 : begin
        result = input_981;
      end
      10'b1111010110 : begin
        result = input_982;
      end
      10'b1111010111 : begin
        result = input_983;
      end
      10'b1111011000 : begin
        result = input_984;
      end
      10'b1111011001 : begin
        result = input_985;
      end
      10'b1111011010 : begin
        result = input_986;
      end
      10'b1111011011 : begin
        result = input_987;
      end
      10'b1111011100 : begin
        result = input_988;
      end
      10'b1111011101 : begin
        result = input_989;
      end
      10'b1111011110 : begin
        result = input_990;
      end
      10'b1111011111 : begin
        result = input_991;
      end
      10'b1111100000 : begin
        result = input_992;
      end
      10'b1111100001 : begin
        result = input_993;
      end
      10'b1111100010 : begin
        result = input_994;
      end
      10'b1111100011 : begin
        result = input_995;
      end
      10'b1111100100 : begin
        result = input_996;
      end
      10'b1111100101 : begin
        result = input_997;
      end
      10'b1111100110 : begin
        result = input_998;
      end
      10'b1111100111 : begin
        result = input_999;
      end
      10'b1111101000 : begin
        result = input_1000;
      end
      10'b1111101001 : begin
        result = input_1001;
      end
      10'b1111101010 : begin
        result = input_1002;
      end
      10'b1111101011 : begin
        result = input_1003;
      end
      10'b1111101100 : begin
        result = input_1004;
      end
      10'b1111101101 : begin
        result = input_1005;
      end
      10'b1111101110 : begin
        result = input_1006;
      end
      10'b1111101111 : begin
        result = input_1007;
      end
      10'b1111110000 : begin
        result = input_1008;
      end
      10'b1111110001 : begin
        result = input_1009;
      end
      10'b1111110010 : begin
        result = input_1010;
      end
      10'b1111110011 : begin
        result = input_1011;
      end
      10'b1111110100 : begin
        result = input_1012;
      end
      10'b1111110101 : begin
        result = input_1013;
      end
      10'b1111110110 : begin
        result = input_1014;
      end
      10'b1111110111 : begin
        result = input_1015;
      end
      10'b1111111000 : begin
        result = input_1016;
      end
      10'b1111111001 : begin
        result = input_1017;
      end
      10'b1111111010 : begin
        result = input_1018;
      end
      10'b1111111011 : begin
        result = input_1019;
      end
      10'b1111111100 : begin
        result = input_1020;
      end
      10'b1111111101 : begin
        result = input_1021;
      end
      10'b1111111110 : begin
        result = input_1022;
      end
      default : begin
        result = input_1023;
      end
    endcase
    MUX_v_14_1024_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i10_1o64_a49ff3631daca65e62d175dd412366e6bd_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Mon May 27 10:56:36 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i10_1o64_a49ff3631daca65e62d175dd412366e6bd
// ------------------------------------------------------------------


module ROM_1i10_1o64_a49ff3631daca65e62d175dd412366e6bd (
  I_1, O_1
);
  input [9:0] I_1;
  output [63:0] O_1;


  wire[56:0] BUTTERFLY_if_BUTTERFLY_if_mux_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign BUTTERFLY_if_BUTTERFLY_if_mux_1_nl = MUX_v_57_1024_2(57'b000000000000000000000000000000000000000000000000000000000,
      57'b000000000000000000000000000000000000000000000000000000000, 57'b111100110101000001001111001100110011111110011101111001101,
      57'b111100110101000001001111001100110011111110011101111001101, 57'b111101101100100000110101111001111001100101000110101000110,
      57'b111011000011111011110001010100110101011101010100101100011, 57'b111011000011111011110001010100110101011101010100101100011,
      57'b111101101100100000110101111001111001100101000110101000110, 57'b111101111011000101001011111001111111101110101110010110000,
      57'b111001000111110001011100000111100011010011010011000001011, 57'b111100001110001110011101100111001101011100110100011001000,
      57'b111101010100110110110011000101001000011101010000110100011, 57'b111101010100110110110011000101001000011101010000110100011,
      57'b111100001110001110011101100111001101011100110100011001000, 57'b111001000111110001011100000111100011010011010011000001011,
      57'b111101111011000101001011111001111111101110101110010110000, 57'b111101111110110001000110110100011110100010010010100100110,
      57'b110111001000101111010011010111100001010011011010000101100, 57'b111100100010011001111001100100101000010010001110111010110,
      57'b111101000101111001000000001101011000101010001011101000001, 57'b111101100001110001011001011110001100000001011110110110001,
      57'b111011110001010110101110100111000000001101111011000111011, 57'b111010010100101000000011000101110110101011001111100000110,
      57'b111101110100111110100000101010110110001100010110111011010, 57'b111101110100111110100000101010110110001100010110111011010,
      57'b111010010100101000000011000101110110101011001111100000110, 57'b111011110001010110101110100111000000001101111011000111011,
      57'b111101100001110001011001011110001100000001011110110110001, 57'b111101000101111001000000001101011000101010001011101000001,
      57'b111100100010011001111001100100101000010010001110111010110, 57'b110111001000101111010011010111100001010011011010000101100,
      57'b111101111110110001000110110100011110100010010010100100110, 57'b111101111111101100010000111100011011110010110110101111110,
      57'b110101001000111110110010111110001000011011101100000010100, 57'b111100101011111010110100100110100100011001110110010100000,
      57'b111100111101101011101111100100010011010101010111110101111, 57'b111101100111011010111101011110100001111001100011101110011,
      57'b111011011010111010001000000001001111000010101110011000000, 57'b111010101100011111001101001110101101010110001111111011101,
      57'b111101110001000010010000100000100111101101000011011100101, 57'b111101111000010100111111011111011100100100011000011010111,
      57'b111001111000110011111100101111011001000010101111100011011, 57'b111100000011100111000011110011001001000101111111111101110,
      57'b111101011011100101000001101000101000110010110111000111110, 57'b111101001101100111110000001000111111100111000011101000001,
      57'b111100011000011111111011111111100111000010111000000110101, 57'b111000010110010000001000001101110100011100110000100111010,
      57'b111101111101001110101010101111111000010001010010100010111, 57'b111101111101001110101010101111111000010001010010100010111,
      57'b111000010110010000001000001101110100011100110000100111010, 57'b111100011000011111111011111111100111000010111000000110101,
      57'b111101001101100111110000001000111111100111000011101000001, 57'b111101011011100101000001101000101000110010110111000111110,
      57'b111100000011100111000011110011001001000101111111111101110, 57'b111001111000110011111100101111011001000010101111100011011,
      57'b111101111000010100111111011111011100100100011000011010111, 57'b111101110001000010010000100000100111101101000011011100101,
      57'b111010101100011111001101001110101101010110001111111011101, 57'b111011011010111010001000000001001111000010101110011000000,
      57'b111101100111011010111101011110100001111001100011101110011, 57'b111100111101101011101111100100010011010101010111110101111,
      57'b111100101011111010110100100110100100011001110110010100000, 57'b110101001000111110110010111110001000011011101100000010100,
      57'b111101111111101100010000111100011011110010110110101111110, 57'b111101111111111011000100001100000100001001100110100001101,
      57'b110011001001000010101010111110111101000110110011001111110, 57'b111100110000100001011011101010101000111010010110011011111,
      57'b111100111001011010000100000110111111011111111111110010110, 57'b111101101010000010011010011010001010011011100100100111010,
      57'b111011001111011110111100101000011101010001110110110001010, 57'b111010111000010001000010100110000111110100100010110011111,
      57'b111101101110110110001001110110110110011001100001000111100, 57'b111101111001110001111001110101100011001001110010110001001,
      57'b111001100000010111000001001101010011111100100111101100011, 57'b111100001000111101011001101010100000110110100101100100011,
      57'b111101011000010010000101001011000000101010000001000000000, 57'b111101010001010011010011110100000010001100010011110000010,
      57'b111100010011011010000010101001100110111010001001011011111, 57'b111000101111000100001010001000100100010110011111111000110,
      57'b111101111100001110110010011111010011100010100101110101001, 57'b111101111110000100110010001110000111000011001111111010011,
      57'b110111111010101100100111001010110101010010111001100001110, 57'b111100011101011111111101000101001001000000101000010111001,
      57'b111101001001110100010001001001001100100100110001111111011, 57'b111101011110101111100000010101100011011111001010100101010,
      57'b111011111100010111010010011011011111110001001101010111010, 57'b111010001000100011101001001100010101100011111011001110111,
      57'b111101110110101110100000011100111011010000100100101100011, 57'b111101110011000101000100011101100010010001110000100010010,
      57'b111010100000100110101110010010100000101110110011000000001, 57'b111011100110001100110111010011001001100011100010001011110,
      57'b111101100100101010100101100100001001101000001000111110101, 57'b111101000001110110000111000001011111111111001011101101110,
      57'b111100100111001101100101010111011111000111110010111101001, 57'b110110010110101010010000010010010110011100001100111110110,
      57'b111101111111010011100110110101101000000011000100000111010, 57'b111101111111010011100110110101101000000011000100000111010,
      57'b110110010110101010010000010010010110011100001100111110110, 57'b111100100111001101100101010111011111000111110010111101001,
      57'b111101000001110110000111000001011111111111001011101101110, 57'b111101100100101010100101100100001001101000001000111110101,
      57'b111011100110001100110111010011001001100011100010001011110, 57'b111010100000100110101110010010100000101110110011000000001,
      57'b111101110011000101000100011101100010010001110000100010010, 57'b111101110110101110100000011100111011010000100100101100011,
      57'b111010001000100011101001001100010101100011111011001110111, 57'b111011111100010111010010011011011111110001001101010111010,
      57'b111101011110101111100000010101100011011111001010100101010, 57'b111101001001110100010001001001001100100100110001111111011,
      57'b111100011101011111111101000101001001000000101000010111001, 57'b110111111010101100100111001010110101010010111001100001110,
      57'b111101111110000100110010001110000111000011001111111010011, 57'b111101111100001110110010011111010011100010100101110101001,
      57'b111000101111000100001010001000100100010110011111111000110, 57'b111100010011011010000010101001100110111010001001011011111,
      57'b111101010001010011010011110100000010001100010011110000010, 57'b111101011000010010000101001011000000101010000001000000000,
      57'b111100001000111101011001101010100000110110100101100100011, 57'b111001100000010111000001001101010011111100100111101100011,
      57'b111101111001110001111001110101100011001001110010110001001, 57'b111101101110110110001001110110110110011001100001000111100,
      57'b111010111000010001000010100110000111110100100010110011111, 57'b111011001111011110111100101000011101010001110110110001010,
      57'b111101101010000010011010011010001010011011100100100111010, 57'b111100111001011010000100000110111111011111111111110010110,
      57'b111100110000100001011011101010101000111010010110011011111, 57'b110011001001000010101010111110111101000110110011001111110,
      57'b111101111111111011000100001100000100001001100110100001101, 57'b111101111111111110110001000010110100110111001001011011011,
      57'b110001001001000011101000111111100110111101100011110000100, 57'b111100110010110010001100100100101111100000111100000111101,
      57'b111100110111001110100010001010100111010101010100010101111, 57'b111101101011010010110000101110011110010011110011010001011,
      57'b111011001001101110010101001100011101111001001001111010111, 57'b111010111110000111010100100110001000111011100110011100111,
      57'b111101101101101100101001001100010001110001010000010011011, 57'b111101111010011100110000000111011000010110010111100101101,
      57'b111001010100000101010000000100101101100000000010001010001, 57'b111100001011100110100110101100011110111101101101101001001,
      57'b111101010110100101011110010011110001000011101010100010001, 57'b111101010011000110000100100011011000000101111101011100010,
      57'b111100010000110100111100110011001001100111110101101011001, 57'b111000111011011011101100111011110010100001011111100110001,
      57'b111101111011101011001100110100011101000010010000001110111, 57'b111101111110011100001010111111101011011011010011001111011,
      57'b110111100001101111000010111000111100111101100001011010101, 57'b111100011111111101101100101010011010001010101011011010100,
      57'b111101000111110111100110010100011111011111001010000001101, 57'b111101100000010001100010000100110011100100101010101001001,
      57'b111011110110111000001100101010010111011110111100011010110, 57'b111010001110100110100010000111111010011001101101100111110,
      57'b111101110101110111101100011001000110111110000101101110100, 57'b111101110100000010111101110101011010011001101000100001101,
      57'b111010011010101000001000011000010111000011000000101010010, 57'b111011101011110010111011101011011100001101110001110001001,
      57'b111101100011001111000101100110100100010000111001110011011, 57'b111101000011111000100000000001111101110100010111010111111,
      57'b111100100100110100100010010011011100110110000100100111001, 57'b110110101111101101101000000001010100110101010010000011001,
      57'b111101111111000011100101011111100101111010101101100001001, 57'b111101111111100001001010101100101100011100111000110101101,
      57'b110101111011001010110111001111001111110000010000011100000, 57'b111100101001100101000001010010010101000110101010110010110,
      57'b111100111111110001110110011100011010101110001011101110001, 57'b111101100110000011111000011110011111111001111110001011100,
      57'b111011100000100100100100111011000000000010001111011100111, 57'b111010100110100011110001001000010011110001110011101101010,
      57'b111101110010000100110101001001011001010111100000101111110, 57'b111101110111100010111100010100011111001000111001111000010,
      57'b111010000010011111011100000001110001101111111110110101110, 57'b111100000000111001111110010000111010011000011111010110111,
      57'b111101011101001011010101001100111001101011001000011010010, 57'b111101001011101110111111011110100110001111101011101000010,
      57'b111100011011000000101100010110001000001100101100111110011, 57'b111000001001110011111000011001110110110101111010101110111,
      57'b111101111101101010111100101110001100101011101011101000001, 57'b111101111100101111111100100100100110010010000100110011011,
      57'b111000100010101010111011010110001001010010011111001011010, 57'b111100010101111101101101100100101111110101111001111101010,
      57'b111101001111011110100001111101111001010011010111110010100, 57'b111101011001111100100110100111110111101010101011100010010,
      57'b111100000110010010111000001001101010111011000100110001111, 57'b111001101100100110100111111100101010001010100001100010001,
      57'b111101111001000100101001011110111011101100011101011011010, 57'b111101101111111101010111001100010001011011011111000101011,
      57'b111010110010011000111110111011101001111110010011111000110, 57'b111011010101001101100100000101011011011010011111111001010,
      57'b111101101000101111110011101110100001111100011010111011100, 57'b111100111011100011110011101011111000000110111001001100001,
      57'b111100101110001110111101110111110011001010000000110001100, 57'b110100010110110000110010101110101100101000101010111001101,
      57'b111101111111110100111001011101111111111101111011101011101, 57'b111101111111110100111001011101111111111101111011101011101,
      57'b110100010110110000110010101110101100101000101010111001101, 57'b111100101110001110111101110111110011001010000000110001100,
      57'b111100111011100011110011101011111000000110111001001100001, 57'b111101101000101111110011101110100001111100011010111011100,
      57'b111011010101001101100100000101011011011010011111111001010, 57'b111010110010011000111110111011101001111110010011111000110,
      57'b111101101111111101010111001100010001011011011111000101011, 57'b111101111001000100101001011110111011101100011101011011010,
      57'b111001101100100110100111111100101010001010100001100010001, 57'b111100000110010010111000001001101010111011000100110001111,
      57'b111101011001111100100110100111110111101010101011100010010, 57'b111101001111011110100001111101111001010011010111110010100,
      57'b111100010101111101101101100100101111110101111001111101010, 57'b111000100010101010111011010110001001010010011111001011010,
      57'b111101111100101111111100100100100110010010000100110011011, 57'b111101111101101010111100101110001100101011101011101000001,
      57'b111000001001110011111000011001110110110101111010101110111, 57'b111100011011000000101100010110001000001100101100111110011,
      57'b111101001011101110111111011110100110001111101011101000010, 57'b111101011101001011010101001100111001101011001000011010010,
      57'b111100000000111001111110010000111010011000011111010110111, 57'b111010000010011111011100000001110001101111111110110101110,
      57'b111101110111100010111100010100011111001000111001111000010, 57'b111101110010000100110101001001011001010111100000101111110,
      57'b111010100110100011110001001000010011110001110011101101010, 57'b111011100000100100100100111011000000000010001111011100111,
      57'b111101100110000011111000011110011111111001111110001011100, 57'b111100111111110001110110011100011010101110001011101110001,
      57'b111100101001100101000001010010010101000110101010110010110, 57'b110101111011001010110111001111001111110000010000011100000,
      57'b111101111111100001001010101100101100011100111000110101101, 57'b111101111111000011100101011111100101111010101101100001001,
      57'b110110101111101101101000000001010100110101010010000011001, 57'b111100100100110100100010010011011100110110000100100111001,
      57'b111101000011111000100000000001111101110100010111010111111, 57'b111101100011001111000101100110100100010000111001110011011,
      57'b111011101011110010111011101011011100001101110001110001001, 57'b111010011010101000001000011000010111000011000000101010010,
      57'b111101110100000010111101110101011010011001101000100001101, 57'b111101110101110111101100011001000110111110000101101110100,
      57'b111010001110100110100010000111111010011001101101100111110, 57'b111011110110111000001100101010010111011110111100011010110,
      57'b111101100000010001100010000100110011100100101010101001001, 57'b111101000111110111100110010100011111011111001010000001101,
      57'b111100011111111101101100101010011010001010101011011010100, 57'b110111100001101111000010111000111100111101100001011010101,
      57'b111101111110011100001010111111101011011011010011001111011, 57'b111101111011101011001100110100011101000010010000001110111,
      57'b111000111011011011101100111011110010100001011111100110001, 57'b111100010000110100111100110011001001100111110101101011001,
      57'b111101010011000110000100100011011000000101111101011100010, 57'b111101010110100101011110010011110001000011101010100010001,
      57'b111100001011100110100110101100011110111101101101101001001, 57'b111001010100000101010000000100101101100000000010001010001,
      57'b111101111010011100110000000111011000010110010111100101101, 57'b111101101101101100101001001100010001110001010000010011011,
      57'b111010111110000111010100100110001000111011100110011100111, 57'b111011001001101110010101001100011101111001001001111010111,
      57'b111101101011010010110000101110011110010011110011010001011, 57'b111100110111001110100010001010100111010101010100010101111,
      57'b111100110010110010001100100100101111100000111100000111101, 57'b110001001001000011101000111111100110111101100011110000100,
      57'b111101111111111110110001000010110100110111001001011011011, 57'b111101111111111111101100010000101100011101000101010010010,
      57'b101111001001000011111000011111110011001110000000001110001, 57'b111100110011111001111011110000100100100011010111100010000,
      57'b111100110110001000000110101110011110000011000001001110101, 57'b111101101011111010000101100000010101110001110110011111001,
      57'b111011000110110101010010100101110110010001010010010110000, 57'b111011000001000001110001110110000010011101010101011000100,
      57'b111101101101000111000001110101001011001101000100110001000, 57'b111101111010110001010001010110001011110001001111010000100,
      57'b111001001101111011100101111110010110111000100001101100110, 57'b111100001100111010101101000001001111100101011100110111000,
      57'b111101010101101110011001001011001000101101100000011010100, 57'b111101010011111110101100001010010100111111110011010011101,
      57'b111100001111100001111000010001011101111001000011000011011, 57'b111001000001100110110011011101000100111000110010011000110,
      57'b111101111011011000011111101111101111101011011101110110111, 57'b111101111110100110111100100010100001000100000101110000100,
      57'b110111010101001111011011100100100010010010101110000000011, 57'b111100100001001011111111100010111100011100110101110110001,
      57'b111101000110111000100010100110011000101101001100011001100, 57'b111101100001000001101111000111111101010010111000110110000,
      57'b111011110100000111110000011101010111110000101000100010100, 57'b111010010001100111011101110101011110000111011101101110001,
      57'b111101110101011011011001011101000111001111010100010001110, 57'b111101110100100001000010000110110000111011111011111110010,
      57'b111010010111101000010001011011010111011000000001110000111, 57'b111011101110100101000111100010100100000011100110001011000,
      57'b111101100010100000100001000000001001010110110100100000111, 57'b111101000100111000111111010011010010011011101010010101010,
      57'b111100100011100111011010100011011100110000111001101000111, 57'b110110111100001110101100001101010010111010101101100100001,
      57'b111101111110111010101001110011111111100011111010001010110, 57'b111101111111100111000001100001111100011010101011101011100,
      57'b110101100010000101000110100010010110000001101011111100011, 57'b111100101010110000001000000111000100101110101000100110111,
      57'b111100111110101111000001101101100110000110011110110110010, 57'b111101100110101111101100110001001100010110011001011110110,
      57'b111011011101101111100111100100011000001001011110100000001, 57'b111010101001100001101100010000000101011110011110000100100,
      57'b111101110001100011110101011101000011100001100111000100101, 57'b111101110111111100010001000001100000010111001010111101100,
      57'b111001111110111001101110000011010110111111110110111111001, 57'b111100000010010000101011000100110101011100010001000011010,
      57'b111101011100011000011100011010010011101010000010011101001, 57'b111101001100101011100111100101110110110000000110100100010,
      57'b111100011001110000100000000001101000011001000111001010111, 57'b111000010000000010001011011010100111011000111101111001111,
      57'b111101111101011101000111010001110010001101100111110111011, 57'b111101111100111111100111001010101101011011011001011001000,
      57'b111000011100011101101101110110000110011011000110100010100, 57'b111100010111001111000000011100011111010001110101000010111,
      57'b111101001110100011011000111110101111010101000000011010101, 57'b111101011010110001000100111111110100100100001010000000101,
      57'b111100000100111101001000001110100000101111100010111100001, 57'b111001110010101101100101000011110000100000001101000011011,
      57'b111101111000101101000111101010011111101110010000001011101, 57'b111101110000100000000110011001010001010011000000010101100,
      57'b111010101111011100010011100110111100111101010011010010011, 57'b111011011000000100000110101101100011111110100000000001001,
      57'b111101101000000101101010011111110101100101011110110010010, 57'b111100111100101000000000001010111010011110101010111100101,
      57'b111100101101000101000110100101010010111010111001001010000, 57'b110100101111111000000000011010010100100001100110101000011,
      57'b111101111111110000111000111011010110110111000000111011111, 57'b111101111111111000010010100011101111100011101001111111000,
      57'b110011111011010010011011100110001110100011100111100000001, 57'b111100101111011000011010010010101100000110111000001110100,
      57'b111100111010011111001010010001101101010001101001010001101, 57'b111101101001011001011001000100000111000001110111110011111,
      57'b111011010010010110100000100100111110111101010000111100101, 57'b111010110101010101001110101111101110001110111111000010111,
      57'b111101101111011010000010111110111110111100100011111011010, 57'b111101111001011011100100111001001000010001001101010011101,
      57'b111001100110011111000110010110011000100101011001010000110, 57'b111100000111101000010011010111011001010101000111001111110,
      57'b111101011001000111100110101000111000000000001001110110100, 57'b111101010000011001001010111101010101110101111100100110111,
      57'b111100010100101100000011100100111011000101001110010101000, 57'b111000101000110111101111110000101100101111100010111110010,
      57'b111101111100011111101010111111111101011100100000111011011, 57'b111101111101111000001011000010111111001000100000110000110,
      57'b111000000011100101010000001000111101110101000001100011101, 57'b111100011100010000100000110000101110111111110101100100010,
      57'b111101001010110001110111111100100100011100110110111010111, 57'b111101011101111101101011111000100100100111000000011101010,
      57'b111011111111000101111011001001011111001110001001000010000, 57'b111010000101100001101100111001111110110111101101110010000,
      57'b111101110111001001000001011100010010110101001110110111100, 57'b111101110010100101001111100000100011100101001111111111100,
      57'b111010100011100101011100010100101010101110001000001010100, 57'b111011100011011000111111101001001100101110000000000001011,
      57'b111101100101010111100000101101001101000001011100100000000, 57'b111101000000110100001101100110011101101010111101011001100,
      57'b111100101000011001100000010011111010110011010000010011011, 57'b110110001010001000000000100110100110101110000100110110011,
      57'b111101111111011010101100011101100101101100111001111000100, 57'b111101111111001011111001110101111001011100011100101000000,
      57'b110110100011001100001000101111001001001110010000010010110, 57'b111100100110000001010000101000101111011000000000000000100,
      57'b111101000010110111100010100011010111010010101100011001100, 57'b111101100011111101000111001010010001000110011110011110011,
      57'b111011101001000000001011011101000111010011101101101011011, 57'b111010011101100111100111011111010000001000001010010110111,
      57'b111101110011100100010011111011011011010101001011101000100, 57'b111101110110010011011001011010011110000111011111110000100,
      57'b111010001011100101010000011010111011101100101000101110111, 57'b111011111001101000000010110010110001111111101000001100111,
      57'b111101011111100000110010011100001010100110111011111011101, 57'b111101001000110110001011001101111110101001001110110100010,
      57'b111100011110101111000001000111000110001011000001101000100, 57'b110111101110001110000111011001011101011101001111111001001,
      57'b111101111110010000110010001101100111111101011011100100001, 57'b111101111011111101010011000101001111001100011110101101110,
      57'b111000110101010000001001100000100111101100100101010110010, 57'b111100010010000111101010111111011100110001010110000011111,
      57'b111101010010001100111100011001000000100011001101011001000, 57'b111101010111011100000010010110100001111000001010001110100,
      57'b111100001010010010001010110101111001100110110110011101011, 57'b111001011010001110011001011101111001111010110011100100010,
      57'b111101111010000111101000010000101111111111001001011011101, 57'b111101101110010001101011111001011010000010000001001100000,
      57'b111010111011001100011010000001111001001000001100011110110, 57'b111011001100100110111000101100001010000011011110111111111,
      57'b111101101010101010110111101010010111010010011111010110001, 57'b111100111000010100100001010110011000101110110110101111010,
      57'b111100110001101010000001110100011000111000001101111101001, 57'b110010010110110010011011010111011111000110000111011111101,
      57'b111101111111111101001110010110100010010110101000110100001, 57'b111101111111111101001110010110100010010110101000110100001,
      57'b110010010110110010011011010111011111000110000111011111101, 57'b111100110001101010000001110100011000111000001101111101001,
      57'b111100111000010100100001010110011000101110110110101111010, 57'b111101101010101010110111101010010111010010011111010110001,
      57'b111011001100100110111000101100001010000011011110111111111, 57'b111010111011001100011010000001111001001000001100011110110,
      57'b111101101110010001101011111001011010000010000001001100000, 57'b111101111010000111101000010000101111111111001001011011101,
      57'b111001011010001110011001011101111001111010110011100100010, 57'b111100001010010010001010110101111001100110110110011101011,
      57'b111101010111011100000010010110100001111000001010001110100, 57'b111101010010001100111100011001000000100011001101011001000,
      57'b111100010010000111101010111111011100110001010110000011111, 57'b111000110101010000001001100000100111101100100101010110010,
      57'b111101111011111101010011000101001111001100011110101101110, 57'b111101111110010000110010001101100111111101011011100100001,
      57'b110111101110001110000111011001011101011101001111111001001, 57'b111100011110101111000001000111000110001011000001101000100,
      57'b111101001000110110001011001101111110101001001110110100010, 57'b111101011111100000110010011100001010100110111011111011101,
      57'b111011111001101000000010110010110001111111101000001100111, 57'b111010001011100101010000011010111011101100101000101110111,
      57'b111101110110010011011001011010011110000111011111110000100, 57'b111101110011100100010011111011011011010101001011101000100,
      57'b111010011101100111100111011111010000001000001010010110111, 57'b111011101001000000001011011101000111010011101101101011011,
      57'b111101100011111101000111001010010001000110011110011110011, 57'b111101000010110111100010100011010111010010101100011001100,
      57'b111100100110000001010000101000101111011000000000000000100, 57'b110110100011001100001000101111001001001110010000010010110,
      57'b111101111111001011111001110101111001011100011100101000000, 57'b111101111111011010101100011101100101101100111001111000100,
      57'b110110001010001000000000100110100110101110000100110110011, 57'b111100101000011001100000010011111010110011010000010011011,
      57'b111101000000110100001101100110011101101010111101011001100, 57'b111101100101010111100000101101001101000001011100100000000,
      57'b111011100011011000111111101001001100101110000000000001011, 57'b111010100011100101011100010100101010101110001000001010100,
      57'b111101110010100101001111100000100011100101001111111111100, 57'b111101110111001001000001011100010010110101001110110111100,
      57'b111010000101100001101100111001111110110111101101110010000, 57'b111011111111000101111011001001011111001110001001000010000,
      57'b111101011101111101101011111000100100100111000000011101010, 57'b111101001010110001110111111100100100011100110110111010111,
      57'b111100011100010000100000110000101110111111110101100100010, 57'b111000000011100101010000001000111101110101000001100011101,
      57'b111101111101111000001011000010111111001000100000110000110, 57'b111101111100011111101010111111111101011100100000111011011,
      57'b111000101000110111101111110000101100101111100010111110010, 57'b111100010100101100000011100100111011000101001110010101000,
      57'b111101010000011001001010111101010101110101111100100110111, 57'b111101011001000111100110101000111000000000001001110110100,
      57'b111100000111101000010011010111011001010101000111001111110, 57'b111001100110011111000110010110011000100101011001010000110,
      57'b111101111001011011100100111001001000010001001101010011101, 57'b111101101111011010000010111110111110111100100011111011010,
      57'b111010110101010101001110101111101110001110111111000010111, 57'b111011010010010110100000100100111110111101010000111100101,
      57'b111101101001011001011001000100000111000001110111110011111, 57'b111100111010011111001010010001101101010001101001010001101,
      57'b111100101111011000011010010010101100000110111000001110100, 57'b110011111011010010011011100110001110100011100111100000001,
      57'b111101111111111000010010100011101111100011101001111111000, 57'b111101111111110000111000111011010110110111000000111011111,
      57'b110100101111111000000000011010010100100001100110101000011, 57'b111100101101000101000110100101010010111010111001001010000,
      57'b111100111100101000000000001010111010011110101010111100101, 57'b111101101000000101101010011111110101100101011110110010010,
      57'b111011011000000100000110101101100011111110100000000001001, 57'b111010101111011100010011100110111100111101010011010010011,
      57'b111101110000100000000110011001010001010011000000010101100, 57'b111101111000101101000111101010011111101110010000001011101,
      57'b111001110010101101100101000011110000100000001101000011011, 57'b111100000100111101001000001110100000101111100010111100001,
      57'b111101011010110001000100111111110100100100001010000000101, 57'b111101001110100011011000111110101111010101000000011010101,
      57'b111100010111001111000000011100011111010001110101000010111, 57'b111000011100011101101101110110000110011011000110100010100,
      57'b111101111100111111100111001010101101011011011001011001000, 57'b111101111101011101000111010001110010001101100111110111011,
      57'b111000010000000010001011011010100111011000111101111001111, 57'b111100011001110000100000000001101000011001000111001010111,
      57'b111101001100101011100111100101110110110000000110100100010, 57'b111101011100011000011100011010010011101010000010011101001,
      57'b111100000010010000101011000100110101011100010001000011010, 57'b111001111110111001101110000011010110111111110110111111001,
      57'b111101110111111100010001000001100000010111001010111101100, 57'b111101110001100011110101011101000011100001100111000100101,
      57'b111010101001100001101100010000000101011110011110000100100, 57'b111011011101101111100111100100011000001001011110100000001,
      57'b111101100110101111101100110001001100010110011001011110110, 57'b111100111110101111000001101101100110000110011110110110010,
      57'b111100101010110000001000000111000100101110101000100110111, 57'b110101100010000101000110100010010110000001101011111100011,
      57'b111101111111100111000001100001111100011010101011101011100, 57'b111101111110111010101001110011111111100011111010001010110,
      57'b110110111100001110101100001101010010111010101101100100001, 57'b111100100011100111011010100011011100110000111001101000111,
      57'b111101000100111000111111010011010010011011101010010101010, 57'b111101100010100000100001000000001001010110110100100000111,
      57'b111011101110100101000111100010100100000011100110001011000, 57'b111010010111101000010001011011010111011000000001110000111,
      57'b111101110100100001000010000110110000111011111011111110010, 57'b111101110101011011011001011101000111001111010100010001110,
      57'b111010010001100111011101110101011110000111011101101110001, 57'b111011110100000111110000011101010111110000101000100010100,
      57'b111101100001000001101111000111111101010010111000110110000, 57'b111101000110111000100010100110011000101101001100011001100,
      57'b111100100001001011111111100010111100011100110101110110001, 57'b110111010101001111011011100100100010010010101110000000011,
      57'b111101111110100110111100100010100001000100000101110000100, 57'b111101111011011000011111101111101111101011011101110110111,
      57'b111001000001100110110011011101000100111000110010011000110, 57'b111100001111100001111000010001011101111001000011000011011,
      57'b111101010011111110101100001010010100111111110011010011101, 57'b111101010101101110011001001011001000101101100000011010100,
      57'b111100001100111010101101000001001111100101011100110111000, 57'b111001001101111011100101111110010110111000100001101100110,
      57'b111101111010110001010001010110001011110001001111010000100, 57'b111101101101000111000001110101001011001101000100110001000,
      57'b111011000001000001110001110110000010011101010101011000100, 57'b111011000110110101010010100101110110010001010010010110000,
      57'b111101101011111010000101100000010101110001110110011111001, 57'b111100110110001000000110101110011110000011000001001110101,
      57'b111100110011111001111011110000100100100011010111100010000, 57'b101111001001000011111000011111110011001110000000001110001,
      57'b111101111111111111101100010000101100011101000101010010010, 57'b111101111111111111111011000100001011000100001110100000010,
      57'b101101001001000011111100010111110110011001010010010111010, 57'b111100110100011101101000111101010101000011001110001110001,
      57'b111100110101100100101110011101101001011111110001010011100, 57'b111101101100001101100010010000100010001011010010001001111,
      57'b111011000101011000100101110000110110101011110110101000100, 57'b111011000010011110110101010101010111100111001000000111111,
      57'b111101101100110100000000011011101100010110011110101000110, 57'b111101111010111011010011011101101010000110110100001011101,
      57'b111001001010110110100100111101001101101100010101011111010, 57'b111100001101100100101000000010111000100110111001110111111,
      57'b111101010101010010101010001111010001011001011100110001110, 57'b111101010100011010110011101101110010101000101101011010010,
      57'b111100001110111000001101101100100110111000100100001110010, 57'b111001000100101100001011100100111110001000001100000000100,
      57'b111101111011001110111010101010110100010000011110011101110, 57'b111101111110101100000110100101101101001110101110010011110,
      57'b110111001110111111011011011101011001001001010100001011100, 57'b111100100001110010111111101011011001010100100001110000000,
      57'b111101000110011000110101001110101000110000100011001010101, 57'b111101100001011001101000101001001001100011110001111110001,
      57'b111011110010101111010100001101101001111001101100000100101, 57'b111010010011000111110011010011001010101010101010010111010,
      57'b111101110101001101000001110010011111001100101100000000000, 57'b111101110100101111110110000110110000000010110101100110000,
      57'b111010010110001000001101001001110100101010100010100100000, 57'b111011101111111101111111101100110101010010100000111011110,
      57'b111101100010001001000001100110001010000011100000000000100, 57'b111101000101011001000011100011110110111100001110110001000,
      57'b111100100011000000101101001101001001010110011001010100010, 57'b110111000010011111000011100010010110000010011000010100001,
      57'b111101111110110101111101001110101000101000101001110001100, 57'b111101111111101001101110001010100101100011011111011010011,
      57'b110101010101100010000000110111101010111111000001100010111, 57'b111100101011010101100001101010001100101110110010010011111,
      57'b111100111110001101011100010011100111000101101001100110011, 57'b111101100111000101011001100100111100110011010000001100000,
      57'b111011011100010100111100000010100111111010101011010010011, 57'b111010101011000000100000000010010111101000110011110110100,
      57'b111101110001010011000111101000100001110010001100101111010, 57'b111101111000001000101101000010100110011110111001110001100,
      57'b111001111011110110111010010000000101111010011100000000010, 57'b111100000010111011111001111101100001100011011100010110111,
      57'b111101011011111110110011010000110111001111001001011101001, 57'b111101001101001001101111110100100001010110000011010110010,
      57'b111100011001001000010000111101100010010011010011000011111, 57'b111000010011001001001100101001101111111010011010000001001,
      57'b111101111101010101111101111001011000011001111110111011100, 57'b111101111101000111001101110101100011110100001011110010001,
      57'b111000011001010110111101111111001010001010001011010100111, 57'b111100010111110111100001001001011010001000001000000010101,
      57'b111101001110000101101000100010000111100000111010111000010, 57'b111101011011001011000111100010100111111011011110001000111,
      57'b111100000100010010001000100100000001100101011000010001100, 57'b111001110101110000110101101000110001011011110001101001000,
      57'b111101111000100001001000010111100100010011000111101011111, 57'b111101110000110001010000000101111110111000110011011011001,
      57'b111010101101111101110011110001011100111011011001110110110, 57'b111011011001011111001011100011101101100110001100101110010,
      57'b111101100111110000011000011101000110011100100011001111011, 57'b111100111101001001111011100000111101111111001011111010010,
      57'b111100101100100000000000111010101111101110010001111011111, 57'b110100111100011011011101010100101100001110100011010000110,
      57'b111101111111101110101001110111011000110111001000101100100, 57'b111101111111111001110000010011100111000101010011001111001,
      57'b110011100010001010100111101001100111001010011101100011101, 57'b111100101111111100111110010111101111001010110101000010000,
      57'b111100111001111100101010110001110000001111001100101000010, 57'b111101101001101101111110001111011110010111111101111011100,
      57'b111011010000111010110010101000011101101010000101011000000, 57'b111010110110110011001100001100011100010100000110010110110,
      57'b111101101111001000001011000001111011011011000110110000001, 57'b111101111001100110110100001011010001110101010111011110000,
      57'b111001100011011011001000001010011010111010111010011011101, 57'b111100001000010010111001001001000110100001010100101010111,
      57'b111101011000101100111010000101010010011001010001011110101, 57'b111101010000110110010011011010010110000001010011101011110,
      57'b111100010100000011000101111101111010011010011110010111010, 57'b111000101011111110000000010000110010101001100101111011110,
      57'b111101111100010111010011100110111110010110100101101111000, 57'b111101111101111110100011100001111000010101000110110001000,
      57'b111000000000011101110100010101101011011111011100001011011, 57'b111100011100111000010001111100011110101100011000000101001,
      57'b111101001010010011001000011100011101011000100101001101100, 57'b111101011110010110101010011001011000011010010001100100111,
      57'b111011111101101110101011101011100001001001101001011011110, 57'b111010000111000010101101101001110000101110100100111001110,
      57'b111101110110111011110101101101010000001111000011001010001, 57'b111101110010110101001110101010101000001000110011111010011,
      57'b111010100010000110001000011011100100010010011011011110000, 57'b111011100100110010111111111000011100001100101001110001001,
      57'b111101100101000001000111100011001101110011100010001001001, 57'b111101000001010101001110000010011111101010100010111111111,
      57'b111100100111110011100110000100101110011001010010010000110, 57'b110110010000011001001011001110100111011010100010001001101,
      57'b111101111111010111001110100100101001100000100000100001111, 57'b111101111111001111110101010000101010010000010110101100000,
      57'b110110011100111011001111100010010110001011010001010011001, 57'b111100100110100111011110001101101010110001001111101111111,
      57'b111101000010010110111000100010001101011111000001111111010, 57'b111101100100010011111010110000111000000101001110000010011,
      57'b111011100111100110100101110101110111000011100110100100001, 57'b111010011111000111001101111101001011011101100001001110001,
      57'b111101110011010100110000111000101010111010101001110100111, 57'b111101110110100001000001101011110100110011001000000001001,
      57'b111010001010000100011111011101111110001101001001101111000, 57'b111011111010111111101111011100110010101101100110110100011,
      57'b111101011111001000001101101100001000100010101010011000001, 57'b111101001001010101010010000011111110001011010100000010101,
      57'b111100011110000111100010001001001100000011100010100011000, 57'b110111110100011101011011111111101111001001010101000111111,
      57'b111101111110001010110111000111011011111011001101011110110, 57'b111101111100000110000111101001010010000001100011000001100,
      57'b111000110010001010001101010000011000111011000001100001101, 57'b111100010010110000111001101001100101110110111000100010000,
      57'b111101010001110000001100001001010010110010011101111000110, 57'b111101010111110111000111111011000100111110101011110110110,
      57'b111100001001100111110100111001111111011100010010101001111, 57'b111001011101010010110001100110100111100010101110110101101,
      57'b111101111001111100110101110111100000110111011110001100101, 57'b111101101110100011111111011110011100010101001000101011010,
      57'b111010111001101110110001111001001001001100001000010010010, 57'b111011001110000010111110101000100000011011111100111110010,
      57'b111101101010010110101101100011011000110000111010100100100, 57'b111100111000110111010110010010110000011100100000110111111,
      57'b111100110001000101110010001001111111011000010001011111111, 57'b110010101111111010100110100100001111110101011001000100110,
      57'b111101111111111100001110001101000011100001100101101110111, 57'b111101111111111110000100101000011110001010011101111010001,
      57'b110001111011010100010100101101010101110011001011111001011, 57'b111100110010001110001010101000011011111110101001101011011,
      57'b111100110111110001100101010011001110010010101101101110101, 57'b111101101010111110111000101110010100010001000101001111111,
      57'b111011001011001010101010110110111101010111001010010001111, 57'b111010111100101001111010111100110000100111101111110101110,
      57'b111101101101111111001111001000011100101010111010110011010, 57'b111101111010010010010001000000110101111001010101110110100,
      57'b111001010111001001111000111010101111100111011100110101011, 57'b111100001010111100011011011100100110110111110001010111100,
      57'b111101010111000000110100011110011010001011110110011101111, 57'b111101010010101001100100100010000100100001111010100100011,
      57'b111100010001011110010110101100110001011000001001111100010, 57'b111000111000010101111110110001101000010001100010011111111,
      57'b111101111011110100010100110011100000110100011001000101010, 57'b111101111110010110100011100000011100100010100001101010100,
      57'b110111100111111110101001100111011001100000111110111000001, 57'b111100011111010110011001111101010101111100000011010000000,
      57'b111101001000010110111100101000011010101110101111011111110, 57'b111101011111111001001110100100101101000011011000101000111,
      57'b111011111000010000001100100000110101111111111011111111110, 57'b111010001101000101111011111111011111010001111001001000011,
      57'b111101110110000101100111101001011000110101111011010110010, 57'b111101110011110011101101100101001101001010001011001011010,
      57'b111010011100000111111010111100011010100111011011010101011, 57'b111011101010011001101000000101011101010000110000010011101,
      57'b111101100011100110001010110001001100111101010101011010111, 57'b111101000011011000000101000011101100110101010000110010101,
      57'b111100100101011010111100101010001011001110010001011110001, 57'b110110101001011100111011101001010010011010100110100001010,
      57'b111101111111000111110100100101011111010011101100010000110, 57'b111101111111011110000000100000010100000100110000110010001,
      57'b110110000011110110110000101001110010001100011000001100100, 57'b111100101000111111010100000011100110110011001101010100110,
      57'b111101000000010011000101101110101011011100101001011111010, 57'b111101100101101101110001000001010000000001101101010011001,
      57'b111011100001111110110110101000111001001100011000100101001, 57'b111010100101000100101001111010001000110111000001011110011,
      57'b111101110010010101000110111111111100000011100111001011110, 57'b111101110111010110000011101001100010100001010010101000100,
      57'b111010000100000000100111000000101111010110110011000011110, 57'b111100000000001110100000011001000001010111000001011100001,
      57'b111101011101100100100100110100000101101101100010000001101, 57'b111101001011010000011111101000010101111010111111111100001,
      57'b111100011011101000101001100011011100000010111111110001101, 57'b111000000110101100100110110111100101100100110011110000110,
      57'b111101111101110001101000110001101011001101010110110110111, 57'b111101111100100111111000101001111100001011010110000001000,
      57'b111000100101110001011000101111111011110011111101010001000, 57'b111100010101010100111011011101000011110101110101101011000,
      57'b111101001111111011111010011110001001100010100100111011110, 57'b111101011001100010001010110100101111100110111101111110011,
      57'b111100000110111101101000010111000010010111100010010110110, 57'b111001101001100010111011101001101001011001011110111101110,
      57'b111101111001010000001011111111100010001100000100111001110, 57'b111101101111101011110001101101010100110111010010110011100,
      57'b111010110011110111001010010011100101011010110001111001011, 57'b111011010011110010000110011010011110110111111001100011011,
      57'b111101101001000100101010111000110111001011010010011100001, 57'b111100111011000001100010100101100001100000100011101100100,
      57'b111100101110110011101111011100111001111100011010001011100, 57'b110100001010001101000010111011011010000101100000101111111,
      57'b111101111111110110101010111100100001001011111110110101110, 57'b111101111111110010111110001000010000010001100000000010100,
      57'b110100100011010100011100101101111111110000110000101111001, 57'b111100101101101010000101100100110010011110111010001001000,
      57'b111100111100000101111101100011011100100001011001101011011, 57'b111101101000011010110011100101111010110011101001010111001,
      57'b111011010110101000111001100010010010111001101110000001001, 57'b111010110000111010101100101011100100010001100001000000010,
      57'b111101110000001110110011011011001001010000000111101010100, 57'b111101111000111000111101010111110001010000100011100001000,
      57'b111001101111101010001011000111111000000010000100110011010, 57'b111100000101101000000010110000111100011111000010111101100,
      57'b111101011010010110111010000001001110111100111100100100101, 57'b111101001111000001000001011101101101101000010010001110010,
      57'b111100010110100110011001111010011010011101001101110111000, 57'b111000011111100100010111101010111110110110100100010010011,
      57'b111101111100110111110110101111100111110111101111000101001, 57'b111101111101100100000110111000110100000011101010101001101,
      57'b111000001100111011000100101000000101111100010010011100111, 57'b111100011010011000101001001010010110000010100110111100001,
      57'b111101001100001101010111011110001010001010111010110010100, 57'b111101011100110001111101000011111110110010001010101011110,
      57'b111100000001100101010111001010101111011011011110110010110, 57'b111010000000111110001100000000110101110011111110111010010,
      57'b111101110111101111101011011100101000111001010001111000000, 57'b111101110001110100011001111101100011101011100111010000101,
      57'b111010101000000010110001111011100000110010111000001001000, 57'b111011011111001010001010100010111111111111100000011011001,
      57'b111101100110011001110111000100000110000101101111010100000, 57'b111100111111010000011111110000111101100000011011010000110,
      57'b111100101010001010100111111110101000101011001110111111100, 57'b110101101110101000000011011111001100000001000111011001001,
      57'b111101111111100100001011000010100111000010011000111101101, 57'b111101111110111111001100100100010111101110011001100000111,
      57'b110110110101111110001101100111110011110011011000100101001, 57'b111100100100001110000001100110000011000001001000111111111,
      57'b111101000100011000110011011100111010010000001101110100001, 57'b111101100010110111110111101011001111111101111100001011010,
      57'b111011101101001100000110001011100111110100001000011011001, 57'b111010011001001000001111110110110001110001011101010101111,
      57'b111101110100010010000100101011011101011010110000000100101, 57'b111101110101101001100111101010001010110111000100000010001,
      57'b111010010000000111000010110000011110101110010011110111110, 57'b111011110101100000000011010010101111100100101011000100000,
      57'b111101100000101001101100111011100010001100101111001010111, 57'b111101000111011000001000010011011010010000110110001001001,
      57'b111100100000100100111001001100110001111010001000010001100, 57'b110111011011011111010011011101100001110001111011001001100,
      57'b111101111110100001101000101011000110110000110000010000111, 57'b111101111011100001111011001000011010010110111111010110111,
      57'b111000111110100001010011110111011110100101100101100011100, 57'b111100010000001011011101010100001011101010110000011010110,
      57'b111101010011100010011100011011110100111010110000011110101, 57'b111101010110001001111111110111101001111101111101011001000,
      57'b111100001100010000101100100011111001110100100011011100101, 57'b111001010001000000011111000011011000110000011000111011010,
      57'b111101111010100111000101100011111101011110010110100000111, 57'b111101101101011001111010000101100111001101000101010111001,
      57'b111010111111100100100110111010011011100110100000111100100, 57'b111011001000010001110111110000001111011110111101111010001,
      57'b111101101011100110011111101010000100011000000110111111111, 57'b111100110110101011010111111101111010010101010111111001101,
      57'b111100110011010110000111100111111010100101011001110000110, 57'b110000010110110010110101100001110010100001001011100000011,
      57'b111101111111111111010011100101100100101111000110001001111, 57'b111101111111111111010011100101100100101111000110001001111,
      57'b110000010110110010110101100001110010100001001011100000011, 57'b111100110011010110000111100111111010100101011001110000110,
      57'b111100110110101011010111111101111010010101010111111001101, 57'b111101101011100110011111101010000100011000000110111111111,
      57'b111011001000010001110111110000001111011110111101111010001, 57'b111010111111100100100110111010011011100110100000111100100,
      57'b111101101101011001111010000101100111001101000101010111001, 57'b111101111010100111000101100011111101011110010110100000111,
      57'b111001010001000000011111000011011000110000011000111011010, 57'b111100001100010000101100100011111001110100100011011100101,
      57'b111101010110001001111111110111101001111101111101011001000, 57'b111101010011100010011100011011110100111010110000011110101,
      57'b111100010000001011011101010100001011101010110000011010110, 57'b111000111110100001010011110111011110100101100101100011100,
      57'b111101111011100001111011001000011010010110111111010110111, 57'b111101111110100001101000101011000110110000110000010000111,
      57'b110111011011011111010011011101100001110001111011001001100, 57'b111100100000100100111001001100110001111010001000010001100,
      57'b111101000111011000001000010011011010010000110110001001001, 57'b111101100000101001101100111011100010001100101111001010111,
      57'b111011110101100000000011010010101111100100101011000100000, 57'b111010010000000111000010110000011110101110010011110111110,
      57'b111101110101101001100111101010001010110111000100000010001, 57'b111101110100010010000100101011011101011010110000000100101,
      57'b111010011001001000001111110110110001110001011101010101111, 57'b111011101101001100000110001011100111110100001000011011001,
      57'b111101100010110111110111101011001111111101111100001011010, 57'b111101000100011000110011011100111010010000001101110100001,
      57'b111100100100001110000001100110000011000001001000111111111, 57'b110110110101111110001101100111110011110011011000100101001,
      57'b111101111110111111001100100100010111101110011001100000111, 57'b111101111111100100001011000010100111000010011000111101101,
      57'b110101101110101000000011011111001100000001000111011001001, 57'b111100101010001010100111111110101000101011001110111111100,
      57'b111100111111010000011111110000111101100000011011010000110, 57'b111101100110011001110111000100000110000101101111010100000,
      57'b111011011111001010001010100010111111111111100000011011001, 57'b111010101000000010110001111011100000110010111000001001000,
      57'b111101110001110100011001111101100011101011100111010000101, 57'b111101110111101111101011011100101000111001010001111000000,
      57'b111010000000111110001100000000110101110011111110111010010, 57'b111100000001100101010111001010101111011011011110110010110,
      57'b111101011100110001111101000011111110110010001010101011110, 57'b111101001100001101010111011110001010001010111010110010100,
      57'b111100011010011000101001001010010110000010100110111100001, 57'b111000001100111011000100101000000101111100010010011100111,
      57'b111101111101100100000110111000110100000011101010101001101, 57'b111101111100110111110110101111100111110111101111000101001,
      57'b111000011111100100010111101010111110110110100100010010011, 57'b111100010110100110011001111010011010011101001101110111000,
      57'b111101001111000001000001011101101101101000010010001110010, 57'b111101011010010110111010000001001110111100111100100100101,
      57'b111100000101101000000010110000111100011111000010111101100, 57'b111001101111101010001011000111111000000010000100110011010,
      57'b111101111000111000111101010111110001010000100011100001000, 57'b111101110000001110110011011011001001010000000111101010100,
      57'b111010110000111010101100101011100100010001100001000000010, 57'b111011010110101000111001100010010010111001101110000001001,
      57'b111101101000011010110011100101111010110011101001010111001, 57'b111100111100000101111101100011011100100001011001101011011,
      57'b111100101101101010000101100100110010011110111010001001000, 57'b110100100011010100011100101101111111110000110000101111001,
      57'b111101111111110010111110001000010000010001100000000010100, 57'b111101111111110110101010111100100001001011111110110101110,
      57'b110100001010001101000010111011011010000101100000101111111, 57'b111100101110110011101111011100111001111100011010001011100,
      57'b111100111011000001100010100101100001100000100011101100100, 57'b111101101001000100101010111000110111001011010010011100001,
      57'b111011010011110010000110011010011110110111111001100011011, 57'b111010110011110111001010010011100101011010110001111001011,
      57'b111101101111101011110001101101010100110111010010110011100, 57'b111101111001010000001011111111100010001100000100111001110,
      57'b111001101001100010111011101001101001011001011110111101110, 57'b111100000110111101101000010111000010010111100010010110110,
      57'b111101011001100010001010110100101111100110111101111110011, 57'b111101001111111011111010011110001001100010100100111011110,
      57'b111100010101010100111011011101000011110101110101101011000, 57'b111000100101110001011000101111111011110011111101010001000,
      57'b111101111100100111111000101001111100001011010110000001000, 57'b111101111101110001101000110001101011001101010110110110111,
      57'b111000000110101100100110110111100101100100110011110000110, 57'b111100011011101000101001100011011100000010111111110001101,
      57'b111101001011010000011111101000010101111010111111111100001, 57'b111101011101100100100100110100000101101101100010000001101,
      57'b111100000000001110100000011001000001010111000001011100001, 57'b111010000100000000100111000000101111010110110011000011110,
      57'b111101110111010110000011101001100010100001010010101000100, 57'b111101110010010101000110111111111100000011100111001011110,
      57'b111010100101000100101001111010001000110111000001011110011, 57'b111011100001111110110110101000111001001100011000100101001,
      57'b111101100101101101110001000001010000000001101101010011001, 57'b111101000000010011000101101110101011011100101001011111010,
      57'b111100101000111111010100000011100110110011001101010100110, 57'b110110000011110110110000101001110010001100011000001100100,
      57'b111101111111011110000000100000010100000100110000110010001, 57'b111101111111000111110100100101011111010011101100010000110,
      57'b110110101001011100111011101001010010011010100110100001010, 57'b111100100101011010111100101010001011001110010001011110001,
      57'b111101000011011000000101000011101100110101010000110010101, 57'b111101100011100110001010110001001100111101010101011010111,
      57'b111011101010011001101000000101011101010000110000010011101, 57'b111010011100000111111010111100011010100111011011010101011,
      57'b111101110011110011101101100101001101001010001011001011010, 57'b111101110110000101100111101001011000110101111011010110010,
      57'b111010001101000101111011111111011111010001111001001000011, 57'b111011111000010000001100100000110101111111111011111111110,
      57'b111101011111111001001110100100101101000011011000101000111, 57'b111101001000010110111100101000011010101110101111011111110,
      57'b111100011111010110011001111101010101111100000011010000000, 57'b110111100111111110101001100111011001100000111110111000001,
      57'b111101111110010110100011100000011100100010100001101010100, 57'b111101111011110100010100110011100000110100011001000101010,
      57'b111000111000010101111110110001101000010001100010011111111, 57'b111100010001011110010110101100110001011000001001111100010,
      57'b111101010010101001100100100010000100100001111010100100011, 57'b111101010111000000110100011110011010001011110110011101111,
      57'b111100001010111100011011011100100110110111110001010111100, 57'b111001010111001001111000111010101111100111011100110101011,
      57'b111101111010010010010001000000110101111001010101110110100, 57'b111101101101111111001111001000011100101010111010110011010,
      57'b111010111100101001111010111100110000100111101111110101110, 57'b111011001011001010101010110110111101010111001010010001111,
      57'b111101101010111110111000101110010100010001000101001111111, 57'b111100110111110001100101010011001110010010101101101110101,
      57'b111100110010001110001010101000011011111110101001101011011, 57'b110001111011010100010100101101010101110011001011111001011,
      57'b111101111111111110000100101000011110001010011101111010001, 57'b111101111111111100001110001101000011100001100101101110111,
      57'b110010101111111010100110100100001111110101011001000100110, 57'b111100110001000101110010001001111111011000010001011111111,
      57'b111100111000110111010110010010110000011100100000110111111, 57'b111101101010010110101101100011011000110000111010100100100,
      57'b111011001110000010111110101000100000011011111100111110010, 57'b111010111001101110110001111001001001001100001000010010010,
      57'b111101101110100011111111011110011100010101001000101011010, 57'b111101111001111100110101110111100000110111011110001100101,
      57'b111001011101010010110001100110100111100010101110110101101, 57'b111100001001100111110100111001111111011100010010101001111,
      57'b111101010111110111000111111011000100111110101011110110110, 57'b111101010001110000001100001001010010110010011101111000110,
      57'b111100010010110000111001101001100101110110111000100010000, 57'b111000110010001010001101010000011000111011000001100001101,
      57'b111101111100000110000111101001010010000001100011000001100, 57'b111101111110001010110111000111011011111011001101011110110,
      57'b110111110100011101011011111111101111001001010101000111111, 57'b111100011110000111100010001001001100000011100010100011000,
      57'b111101001001010101010010000011111110001011010100000010101, 57'b111101011111001000001101101100001000100010101010011000001,
      57'b111011111010111111101111011100110010101101100110110100011, 57'b111010001010000100011111011101111110001101001001101111000,
      57'b111101110110100001000001101011110100110011001000000001001, 57'b111101110011010100110000111000101010111010101001110100111,
      57'b111010011111000111001101111101001011011101100001001110001, 57'b111011100111100110100101110101110111000011100110100100001,
      57'b111101100100010011111010110000111000000101001110000010011, 57'b111101000010010110111000100010001101011111000001111111010,
      57'b111100100110100111011110001101101010110001001111101111111, 57'b110110011100111011001111100010010110001011010001010011001,
      57'b111101111111001111110101010000101010010000010110101100000, 57'b111101111111010111001110100100101001100000100000100001111,
      57'b110110010000011001001011001110100111011010100010001001101, 57'b111100100111110011100110000100101110011001010010010000110,
      57'b111101000001010101001110000010011111101010100010111111111, 57'b111101100101000001000111100011001101110011100010001001001,
      57'b111011100100110010111111111000011100001100101001110001001, 57'b111010100010000110001000011011100100010010011011011110000,
      57'b111101110010110101001110101010101000001000110011111010011, 57'b111101110110111011110101101101010000001111000011001010001,
      57'b111010000111000010101101101001110000101110100100111001110, 57'b111011111101101110101011101011100001001001101001011011110,
      57'b111101011110010110101010011001011000011010010001100100111, 57'b111101001010010011001000011100011101011000100101001101100,
      57'b111100011100111000010001111100011110101100011000000101001, 57'b111000000000011101110100010101101011011111011100001011011,
      57'b111101111101111110100011100001111000010101000110110001000, 57'b111101111100010111010011100110111110010110100101101111000,
      57'b111000101011111110000000010000110010101001100101111011110, 57'b111100010100000011000101111101111010011010011110010111010,
      57'b111101010000110110010011011010010110000001010011101011110, 57'b111101011000101100111010000101010010011001010001011110101,
      57'b111100001000010010111001001001000110100001010100101010111, 57'b111001100011011011001000001010011010111010111010011011101,
      57'b111101111001100110110100001011010001110101010111011110000, 57'b111101101111001000001011000001111011011011000110110000001,
      57'b111010110110110011001100001100011100010100000110010110110, 57'b111011010000111010110010101000011101101010000101011000000,
      57'b111101101001101101111110001111011110010111111101111011100, 57'b111100111001111100101010110001110000001111001100101000010,
      57'b111100101111111100111110010111101111001010110101000010000, 57'b110011100010001010100111101001100111001010011101100011101,
      57'b111101111111111001110000010011100111000101010011001111001, 57'b111101111111101110101001110111011000110111001000101100100,
      57'b110100111100011011011101010100101100001110100011010000110, 57'b111100101100100000000000111010101111101110010001111011111,
      57'b111100111101001001111011100000111101111111001011111010010, 57'b111101100111110000011000011101000110011100100011001111011,
      57'b111011011001011111001011100011101101100110001100101110010, 57'b111010101101111101110011110001011100111011011001110110110,
      57'b111101110000110001010000000101111110111000110011011011001, 57'b111101111000100001001000010111100100010011000111101011111,
      57'b111001110101110000110101101000110001011011110001101001000, 57'b111100000100010010001000100100000001100101011000010001100,
      57'b111101011011001011000111100010100111111011011110001000111, 57'b111101001110000101101000100010000111100000111010111000010,
      57'b111100010111110111100001001001011010001000001000000010101, 57'b111000011001010110111101111111001010001010001011010100111,
      57'b111101111101000111001101110101100011110100001011110010001, 57'b111101111101010101111101111001011000011001111110111011100,
      57'b111000010011001001001100101001101111111010011010000001001, 57'b111100011001001000010000111101100010010011010011000011111,
      57'b111101001101001001101111110100100001010110000011010110010, 57'b111101011011111110110011010000110111001111001001011101001,
      57'b111100000010111011111001111101100001100011011100010110111, 57'b111001111011110110111010010000000101111010011100000000010,
      57'b111101111000001000101101000010100110011110111001110001100, 57'b111101110001010011000111101000100001110010001100101111010,
      57'b111010101011000000100000000010010111101000110011110110100, 57'b111011011100010100111100000010100111111010101011010010011,
      57'b111101100111000101011001100100111100110011010000001100000, 57'b111100111110001101011100010011100111000101101001100110011,
      57'b111100101011010101100001101010001100101110110010010011111, 57'b110101010101100010000000110111101010111111000001100010111,
      57'b111101111111101001101110001010100101100011011111011010011, 57'b111101111110110101111101001110101000101000101001110001100,
      57'b110111000010011111000011100010010110000010011000010100001, 57'b111100100011000000101101001101001001010110011001010100010,
      57'b111101000101011001000011100011110110111100001110110001000, 57'b111101100010001001000001100110001010000011100000000000100,
      57'b111011101111111101111111101100110101010010100000111011110, 57'b111010010110001000001101001001110100101010100010100100000,
      57'b111101110100101111110110000110110000000010110101100110000, 57'b111101110101001101000001110010011111001100101100000000000,
      57'b111010010011000111110011010011001010101010101010010111010, 57'b111011110010101111010100001101101001111001101100000100101,
      57'b111101100001011001101000101001001001100011110001111110001, 57'b111101000110011000110101001110101000110000100011001010101,
      57'b111100100001110010111111101011011001010100100001110000000, 57'b110111001110111111011011011101011001001001010100001011100,
      57'b111101111110101100000110100101101101001110101110010011110, 57'b111101111011001110111010101010110100010000011110011101110,
      57'b111001000100101100001011100100111110001000001100000000100, 57'b111100001110111000001101101100100110111000100100001110010,
      57'b111101010100011010110011101101110010101000101101011010010, 57'b111101010101010010101010001111010001011001011100110001110,
      57'b111100001101100100101000000010111000100110111001110111111, 57'b111001001010110110100100111101001101101100010101011111010,
      57'b111101111010111011010011011101101010000110110100001011101, 57'b111101101100110100000000011011101100010110011110101000110,
      57'b111011000010011110110101010101010111100111001000000111111, 57'b111011000101011000100101110000110110101011110110101000100,
      57'b111101101100001101100010010000100010001011010010001001111, 57'b111100110101100100101110011101101001011111110001010011100,
      57'b111100110100011101101000111101010101000011001110001110001, 57'b101101001001000011111100010111110110011001010010010111010,
      57'b111101111111111111111011000100001011000100001110100000010, I_1);
  assign O_1 = {(I_1[0]) , 1'b0 , (signext_62_57(BUTTERFLY_if_BUTTERFLY_if_mux_1_nl))};

  function automatic [56:0] MUX_v_57_1024_2;
    input [56:0] input_0;
    input [56:0] input_1;
    input [56:0] input_2;
    input [56:0] input_3;
    input [56:0] input_4;
    input [56:0] input_5;
    input [56:0] input_6;
    input [56:0] input_7;
    input [56:0] input_8;
    input [56:0] input_9;
    input [56:0] input_10;
    input [56:0] input_11;
    input [56:0] input_12;
    input [56:0] input_13;
    input [56:0] input_14;
    input [56:0] input_15;
    input [56:0] input_16;
    input [56:0] input_17;
    input [56:0] input_18;
    input [56:0] input_19;
    input [56:0] input_20;
    input [56:0] input_21;
    input [56:0] input_22;
    input [56:0] input_23;
    input [56:0] input_24;
    input [56:0] input_25;
    input [56:0] input_26;
    input [56:0] input_27;
    input [56:0] input_28;
    input [56:0] input_29;
    input [56:0] input_30;
    input [56:0] input_31;
    input [56:0] input_32;
    input [56:0] input_33;
    input [56:0] input_34;
    input [56:0] input_35;
    input [56:0] input_36;
    input [56:0] input_37;
    input [56:0] input_38;
    input [56:0] input_39;
    input [56:0] input_40;
    input [56:0] input_41;
    input [56:0] input_42;
    input [56:0] input_43;
    input [56:0] input_44;
    input [56:0] input_45;
    input [56:0] input_46;
    input [56:0] input_47;
    input [56:0] input_48;
    input [56:0] input_49;
    input [56:0] input_50;
    input [56:0] input_51;
    input [56:0] input_52;
    input [56:0] input_53;
    input [56:0] input_54;
    input [56:0] input_55;
    input [56:0] input_56;
    input [56:0] input_57;
    input [56:0] input_58;
    input [56:0] input_59;
    input [56:0] input_60;
    input [56:0] input_61;
    input [56:0] input_62;
    input [56:0] input_63;
    input [56:0] input_64;
    input [56:0] input_65;
    input [56:0] input_66;
    input [56:0] input_67;
    input [56:0] input_68;
    input [56:0] input_69;
    input [56:0] input_70;
    input [56:0] input_71;
    input [56:0] input_72;
    input [56:0] input_73;
    input [56:0] input_74;
    input [56:0] input_75;
    input [56:0] input_76;
    input [56:0] input_77;
    input [56:0] input_78;
    input [56:0] input_79;
    input [56:0] input_80;
    input [56:0] input_81;
    input [56:0] input_82;
    input [56:0] input_83;
    input [56:0] input_84;
    input [56:0] input_85;
    input [56:0] input_86;
    input [56:0] input_87;
    input [56:0] input_88;
    input [56:0] input_89;
    input [56:0] input_90;
    input [56:0] input_91;
    input [56:0] input_92;
    input [56:0] input_93;
    input [56:0] input_94;
    input [56:0] input_95;
    input [56:0] input_96;
    input [56:0] input_97;
    input [56:0] input_98;
    input [56:0] input_99;
    input [56:0] input_100;
    input [56:0] input_101;
    input [56:0] input_102;
    input [56:0] input_103;
    input [56:0] input_104;
    input [56:0] input_105;
    input [56:0] input_106;
    input [56:0] input_107;
    input [56:0] input_108;
    input [56:0] input_109;
    input [56:0] input_110;
    input [56:0] input_111;
    input [56:0] input_112;
    input [56:0] input_113;
    input [56:0] input_114;
    input [56:0] input_115;
    input [56:0] input_116;
    input [56:0] input_117;
    input [56:0] input_118;
    input [56:0] input_119;
    input [56:0] input_120;
    input [56:0] input_121;
    input [56:0] input_122;
    input [56:0] input_123;
    input [56:0] input_124;
    input [56:0] input_125;
    input [56:0] input_126;
    input [56:0] input_127;
    input [56:0] input_128;
    input [56:0] input_129;
    input [56:0] input_130;
    input [56:0] input_131;
    input [56:0] input_132;
    input [56:0] input_133;
    input [56:0] input_134;
    input [56:0] input_135;
    input [56:0] input_136;
    input [56:0] input_137;
    input [56:0] input_138;
    input [56:0] input_139;
    input [56:0] input_140;
    input [56:0] input_141;
    input [56:0] input_142;
    input [56:0] input_143;
    input [56:0] input_144;
    input [56:0] input_145;
    input [56:0] input_146;
    input [56:0] input_147;
    input [56:0] input_148;
    input [56:0] input_149;
    input [56:0] input_150;
    input [56:0] input_151;
    input [56:0] input_152;
    input [56:0] input_153;
    input [56:0] input_154;
    input [56:0] input_155;
    input [56:0] input_156;
    input [56:0] input_157;
    input [56:0] input_158;
    input [56:0] input_159;
    input [56:0] input_160;
    input [56:0] input_161;
    input [56:0] input_162;
    input [56:0] input_163;
    input [56:0] input_164;
    input [56:0] input_165;
    input [56:0] input_166;
    input [56:0] input_167;
    input [56:0] input_168;
    input [56:0] input_169;
    input [56:0] input_170;
    input [56:0] input_171;
    input [56:0] input_172;
    input [56:0] input_173;
    input [56:0] input_174;
    input [56:0] input_175;
    input [56:0] input_176;
    input [56:0] input_177;
    input [56:0] input_178;
    input [56:0] input_179;
    input [56:0] input_180;
    input [56:0] input_181;
    input [56:0] input_182;
    input [56:0] input_183;
    input [56:0] input_184;
    input [56:0] input_185;
    input [56:0] input_186;
    input [56:0] input_187;
    input [56:0] input_188;
    input [56:0] input_189;
    input [56:0] input_190;
    input [56:0] input_191;
    input [56:0] input_192;
    input [56:0] input_193;
    input [56:0] input_194;
    input [56:0] input_195;
    input [56:0] input_196;
    input [56:0] input_197;
    input [56:0] input_198;
    input [56:0] input_199;
    input [56:0] input_200;
    input [56:0] input_201;
    input [56:0] input_202;
    input [56:0] input_203;
    input [56:0] input_204;
    input [56:0] input_205;
    input [56:0] input_206;
    input [56:0] input_207;
    input [56:0] input_208;
    input [56:0] input_209;
    input [56:0] input_210;
    input [56:0] input_211;
    input [56:0] input_212;
    input [56:0] input_213;
    input [56:0] input_214;
    input [56:0] input_215;
    input [56:0] input_216;
    input [56:0] input_217;
    input [56:0] input_218;
    input [56:0] input_219;
    input [56:0] input_220;
    input [56:0] input_221;
    input [56:0] input_222;
    input [56:0] input_223;
    input [56:0] input_224;
    input [56:0] input_225;
    input [56:0] input_226;
    input [56:0] input_227;
    input [56:0] input_228;
    input [56:0] input_229;
    input [56:0] input_230;
    input [56:0] input_231;
    input [56:0] input_232;
    input [56:0] input_233;
    input [56:0] input_234;
    input [56:0] input_235;
    input [56:0] input_236;
    input [56:0] input_237;
    input [56:0] input_238;
    input [56:0] input_239;
    input [56:0] input_240;
    input [56:0] input_241;
    input [56:0] input_242;
    input [56:0] input_243;
    input [56:0] input_244;
    input [56:0] input_245;
    input [56:0] input_246;
    input [56:0] input_247;
    input [56:0] input_248;
    input [56:0] input_249;
    input [56:0] input_250;
    input [56:0] input_251;
    input [56:0] input_252;
    input [56:0] input_253;
    input [56:0] input_254;
    input [56:0] input_255;
    input [56:0] input_256;
    input [56:0] input_257;
    input [56:0] input_258;
    input [56:0] input_259;
    input [56:0] input_260;
    input [56:0] input_261;
    input [56:0] input_262;
    input [56:0] input_263;
    input [56:0] input_264;
    input [56:0] input_265;
    input [56:0] input_266;
    input [56:0] input_267;
    input [56:0] input_268;
    input [56:0] input_269;
    input [56:0] input_270;
    input [56:0] input_271;
    input [56:0] input_272;
    input [56:0] input_273;
    input [56:0] input_274;
    input [56:0] input_275;
    input [56:0] input_276;
    input [56:0] input_277;
    input [56:0] input_278;
    input [56:0] input_279;
    input [56:0] input_280;
    input [56:0] input_281;
    input [56:0] input_282;
    input [56:0] input_283;
    input [56:0] input_284;
    input [56:0] input_285;
    input [56:0] input_286;
    input [56:0] input_287;
    input [56:0] input_288;
    input [56:0] input_289;
    input [56:0] input_290;
    input [56:0] input_291;
    input [56:0] input_292;
    input [56:0] input_293;
    input [56:0] input_294;
    input [56:0] input_295;
    input [56:0] input_296;
    input [56:0] input_297;
    input [56:0] input_298;
    input [56:0] input_299;
    input [56:0] input_300;
    input [56:0] input_301;
    input [56:0] input_302;
    input [56:0] input_303;
    input [56:0] input_304;
    input [56:0] input_305;
    input [56:0] input_306;
    input [56:0] input_307;
    input [56:0] input_308;
    input [56:0] input_309;
    input [56:0] input_310;
    input [56:0] input_311;
    input [56:0] input_312;
    input [56:0] input_313;
    input [56:0] input_314;
    input [56:0] input_315;
    input [56:0] input_316;
    input [56:0] input_317;
    input [56:0] input_318;
    input [56:0] input_319;
    input [56:0] input_320;
    input [56:0] input_321;
    input [56:0] input_322;
    input [56:0] input_323;
    input [56:0] input_324;
    input [56:0] input_325;
    input [56:0] input_326;
    input [56:0] input_327;
    input [56:0] input_328;
    input [56:0] input_329;
    input [56:0] input_330;
    input [56:0] input_331;
    input [56:0] input_332;
    input [56:0] input_333;
    input [56:0] input_334;
    input [56:0] input_335;
    input [56:0] input_336;
    input [56:0] input_337;
    input [56:0] input_338;
    input [56:0] input_339;
    input [56:0] input_340;
    input [56:0] input_341;
    input [56:0] input_342;
    input [56:0] input_343;
    input [56:0] input_344;
    input [56:0] input_345;
    input [56:0] input_346;
    input [56:0] input_347;
    input [56:0] input_348;
    input [56:0] input_349;
    input [56:0] input_350;
    input [56:0] input_351;
    input [56:0] input_352;
    input [56:0] input_353;
    input [56:0] input_354;
    input [56:0] input_355;
    input [56:0] input_356;
    input [56:0] input_357;
    input [56:0] input_358;
    input [56:0] input_359;
    input [56:0] input_360;
    input [56:0] input_361;
    input [56:0] input_362;
    input [56:0] input_363;
    input [56:0] input_364;
    input [56:0] input_365;
    input [56:0] input_366;
    input [56:0] input_367;
    input [56:0] input_368;
    input [56:0] input_369;
    input [56:0] input_370;
    input [56:0] input_371;
    input [56:0] input_372;
    input [56:0] input_373;
    input [56:0] input_374;
    input [56:0] input_375;
    input [56:0] input_376;
    input [56:0] input_377;
    input [56:0] input_378;
    input [56:0] input_379;
    input [56:0] input_380;
    input [56:0] input_381;
    input [56:0] input_382;
    input [56:0] input_383;
    input [56:0] input_384;
    input [56:0] input_385;
    input [56:0] input_386;
    input [56:0] input_387;
    input [56:0] input_388;
    input [56:0] input_389;
    input [56:0] input_390;
    input [56:0] input_391;
    input [56:0] input_392;
    input [56:0] input_393;
    input [56:0] input_394;
    input [56:0] input_395;
    input [56:0] input_396;
    input [56:0] input_397;
    input [56:0] input_398;
    input [56:0] input_399;
    input [56:0] input_400;
    input [56:0] input_401;
    input [56:0] input_402;
    input [56:0] input_403;
    input [56:0] input_404;
    input [56:0] input_405;
    input [56:0] input_406;
    input [56:0] input_407;
    input [56:0] input_408;
    input [56:0] input_409;
    input [56:0] input_410;
    input [56:0] input_411;
    input [56:0] input_412;
    input [56:0] input_413;
    input [56:0] input_414;
    input [56:0] input_415;
    input [56:0] input_416;
    input [56:0] input_417;
    input [56:0] input_418;
    input [56:0] input_419;
    input [56:0] input_420;
    input [56:0] input_421;
    input [56:0] input_422;
    input [56:0] input_423;
    input [56:0] input_424;
    input [56:0] input_425;
    input [56:0] input_426;
    input [56:0] input_427;
    input [56:0] input_428;
    input [56:0] input_429;
    input [56:0] input_430;
    input [56:0] input_431;
    input [56:0] input_432;
    input [56:0] input_433;
    input [56:0] input_434;
    input [56:0] input_435;
    input [56:0] input_436;
    input [56:0] input_437;
    input [56:0] input_438;
    input [56:0] input_439;
    input [56:0] input_440;
    input [56:0] input_441;
    input [56:0] input_442;
    input [56:0] input_443;
    input [56:0] input_444;
    input [56:0] input_445;
    input [56:0] input_446;
    input [56:0] input_447;
    input [56:0] input_448;
    input [56:0] input_449;
    input [56:0] input_450;
    input [56:0] input_451;
    input [56:0] input_452;
    input [56:0] input_453;
    input [56:0] input_454;
    input [56:0] input_455;
    input [56:0] input_456;
    input [56:0] input_457;
    input [56:0] input_458;
    input [56:0] input_459;
    input [56:0] input_460;
    input [56:0] input_461;
    input [56:0] input_462;
    input [56:0] input_463;
    input [56:0] input_464;
    input [56:0] input_465;
    input [56:0] input_466;
    input [56:0] input_467;
    input [56:0] input_468;
    input [56:0] input_469;
    input [56:0] input_470;
    input [56:0] input_471;
    input [56:0] input_472;
    input [56:0] input_473;
    input [56:0] input_474;
    input [56:0] input_475;
    input [56:0] input_476;
    input [56:0] input_477;
    input [56:0] input_478;
    input [56:0] input_479;
    input [56:0] input_480;
    input [56:0] input_481;
    input [56:0] input_482;
    input [56:0] input_483;
    input [56:0] input_484;
    input [56:0] input_485;
    input [56:0] input_486;
    input [56:0] input_487;
    input [56:0] input_488;
    input [56:0] input_489;
    input [56:0] input_490;
    input [56:0] input_491;
    input [56:0] input_492;
    input [56:0] input_493;
    input [56:0] input_494;
    input [56:0] input_495;
    input [56:0] input_496;
    input [56:0] input_497;
    input [56:0] input_498;
    input [56:0] input_499;
    input [56:0] input_500;
    input [56:0] input_501;
    input [56:0] input_502;
    input [56:0] input_503;
    input [56:0] input_504;
    input [56:0] input_505;
    input [56:0] input_506;
    input [56:0] input_507;
    input [56:0] input_508;
    input [56:0] input_509;
    input [56:0] input_510;
    input [56:0] input_511;
    input [56:0] input_512;
    input [56:0] input_513;
    input [56:0] input_514;
    input [56:0] input_515;
    input [56:0] input_516;
    input [56:0] input_517;
    input [56:0] input_518;
    input [56:0] input_519;
    input [56:0] input_520;
    input [56:0] input_521;
    input [56:0] input_522;
    input [56:0] input_523;
    input [56:0] input_524;
    input [56:0] input_525;
    input [56:0] input_526;
    input [56:0] input_527;
    input [56:0] input_528;
    input [56:0] input_529;
    input [56:0] input_530;
    input [56:0] input_531;
    input [56:0] input_532;
    input [56:0] input_533;
    input [56:0] input_534;
    input [56:0] input_535;
    input [56:0] input_536;
    input [56:0] input_537;
    input [56:0] input_538;
    input [56:0] input_539;
    input [56:0] input_540;
    input [56:0] input_541;
    input [56:0] input_542;
    input [56:0] input_543;
    input [56:0] input_544;
    input [56:0] input_545;
    input [56:0] input_546;
    input [56:0] input_547;
    input [56:0] input_548;
    input [56:0] input_549;
    input [56:0] input_550;
    input [56:0] input_551;
    input [56:0] input_552;
    input [56:0] input_553;
    input [56:0] input_554;
    input [56:0] input_555;
    input [56:0] input_556;
    input [56:0] input_557;
    input [56:0] input_558;
    input [56:0] input_559;
    input [56:0] input_560;
    input [56:0] input_561;
    input [56:0] input_562;
    input [56:0] input_563;
    input [56:0] input_564;
    input [56:0] input_565;
    input [56:0] input_566;
    input [56:0] input_567;
    input [56:0] input_568;
    input [56:0] input_569;
    input [56:0] input_570;
    input [56:0] input_571;
    input [56:0] input_572;
    input [56:0] input_573;
    input [56:0] input_574;
    input [56:0] input_575;
    input [56:0] input_576;
    input [56:0] input_577;
    input [56:0] input_578;
    input [56:0] input_579;
    input [56:0] input_580;
    input [56:0] input_581;
    input [56:0] input_582;
    input [56:0] input_583;
    input [56:0] input_584;
    input [56:0] input_585;
    input [56:0] input_586;
    input [56:0] input_587;
    input [56:0] input_588;
    input [56:0] input_589;
    input [56:0] input_590;
    input [56:0] input_591;
    input [56:0] input_592;
    input [56:0] input_593;
    input [56:0] input_594;
    input [56:0] input_595;
    input [56:0] input_596;
    input [56:0] input_597;
    input [56:0] input_598;
    input [56:0] input_599;
    input [56:0] input_600;
    input [56:0] input_601;
    input [56:0] input_602;
    input [56:0] input_603;
    input [56:0] input_604;
    input [56:0] input_605;
    input [56:0] input_606;
    input [56:0] input_607;
    input [56:0] input_608;
    input [56:0] input_609;
    input [56:0] input_610;
    input [56:0] input_611;
    input [56:0] input_612;
    input [56:0] input_613;
    input [56:0] input_614;
    input [56:0] input_615;
    input [56:0] input_616;
    input [56:0] input_617;
    input [56:0] input_618;
    input [56:0] input_619;
    input [56:0] input_620;
    input [56:0] input_621;
    input [56:0] input_622;
    input [56:0] input_623;
    input [56:0] input_624;
    input [56:0] input_625;
    input [56:0] input_626;
    input [56:0] input_627;
    input [56:0] input_628;
    input [56:0] input_629;
    input [56:0] input_630;
    input [56:0] input_631;
    input [56:0] input_632;
    input [56:0] input_633;
    input [56:0] input_634;
    input [56:0] input_635;
    input [56:0] input_636;
    input [56:0] input_637;
    input [56:0] input_638;
    input [56:0] input_639;
    input [56:0] input_640;
    input [56:0] input_641;
    input [56:0] input_642;
    input [56:0] input_643;
    input [56:0] input_644;
    input [56:0] input_645;
    input [56:0] input_646;
    input [56:0] input_647;
    input [56:0] input_648;
    input [56:0] input_649;
    input [56:0] input_650;
    input [56:0] input_651;
    input [56:0] input_652;
    input [56:0] input_653;
    input [56:0] input_654;
    input [56:0] input_655;
    input [56:0] input_656;
    input [56:0] input_657;
    input [56:0] input_658;
    input [56:0] input_659;
    input [56:0] input_660;
    input [56:0] input_661;
    input [56:0] input_662;
    input [56:0] input_663;
    input [56:0] input_664;
    input [56:0] input_665;
    input [56:0] input_666;
    input [56:0] input_667;
    input [56:0] input_668;
    input [56:0] input_669;
    input [56:0] input_670;
    input [56:0] input_671;
    input [56:0] input_672;
    input [56:0] input_673;
    input [56:0] input_674;
    input [56:0] input_675;
    input [56:0] input_676;
    input [56:0] input_677;
    input [56:0] input_678;
    input [56:0] input_679;
    input [56:0] input_680;
    input [56:0] input_681;
    input [56:0] input_682;
    input [56:0] input_683;
    input [56:0] input_684;
    input [56:0] input_685;
    input [56:0] input_686;
    input [56:0] input_687;
    input [56:0] input_688;
    input [56:0] input_689;
    input [56:0] input_690;
    input [56:0] input_691;
    input [56:0] input_692;
    input [56:0] input_693;
    input [56:0] input_694;
    input [56:0] input_695;
    input [56:0] input_696;
    input [56:0] input_697;
    input [56:0] input_698;
    input [56:0] input_699;
    input [56:0] input_700;
    input [56:0] input_701;
    input [56:0] input_702;
    input [56:0] input_703;
    input [56:0] input_704;
    input [56:0] input_705;
    input [56:0] input_706;
    input [56:0] input_707;
    input [56:0] input_708;
    input [56:0] input_709;
    input [56:0] input_710;
    input [56:0] input_711;
    input [56:0] input_712;
    input [56:0] input_713;
    input [56:0] input_714;
    input [56:0] input_715;
    input [56:0] input_716;
    input [56:0] input_717;
    input [56:0] input_718;
    input [56:0] input_719;
    input [56:0] input_720;
    input [56:0] input_721;
    input [56:0] input_722;
    input [56:0] input_723;
    input [56:0] input_724;
    input [56:0] input_725;
    input [56:0] input_726;
    input [56:0] input_727;
    input [56:0] input_728;
    input [56:0] input_729;
    input [56:0] input_730;
    input [56:0] input_731;
    input [56:0] input_732;
    input [56:0] input_733;
    input [56:0] input_734;
    input [56:0] input_735;
    input [56:0] input_736;
    input [56:0] input_737;
    input [56:0] input_738;
    input [56:0] input_739;
    input [56:0] input_740;
    input [56:0] input_741;
    input [56:0] input_742;
    input [56:0] input_743;
    input [56:0] input_744;
    input [56:0] input_745;
    input [56:0] input_746;
    input [56:0] input_747;
    input [56:0] input_748;
    input [56:0] input_749;
    input [56:0] input_750;
    input [56:0] input_751;
    input [56:0] input_752;
    input [56:0] input_753;
    input [56:0] input_754;
    input [56:0] input_755;
    input [56:0] input_756;
    input [56:0] input_757;
    input [56:0] input_758;
    input [56:0] input_759;
    input [56:0] input_760;
    input [56:0] input_761;
    input [56:0] input_762;
    input [56:0] input_763;
    input [56:0] input_764;
    input [56:0] input_765;
    input [56:0] input_766;
    input [56:0] input_767;
    input [56:0] input_768;
    input [56:0] input_769;
    input [56:0] input_770;
    input [56:0] input_771;
    input [56:0] input_772;
    input [56:0] input_773;
    input [56:0] input_774;
    input [56:0] input_775;
    input [56:0] input_776;
    input [56:0] input_777;
    input [56:0] input_778;
    input [56:0] input_779;
    input [56:0] input_780;
    input [56:0] input_781;
    input [56:0] input_782;
    input [56:0] input_783;
    input [56:0] input_784;
    input [56:0] input_785;
    input [56:0] input_786;
    input [56:0] input_787;
    input [56:0] input_788;
    input [56:0] input_789;
    input [56:0] input_790;
    input [56:0] input_791;
    input [56:0] input_792;
    input [56:0] input_793;
    input [56:0] input_794;
    input [56:0] input_795;
    input [56:0] input_796;
    input [56:0] input_797;
    input [56:0] input_798;
    input [56:0] input_799;
    input [56:0] input_800;
    input [56:0] input_801;
    input [56:0] input_802;
    input [56:0] input_803;
    input [56:0] input_804;
    input [56:0] input_805;
    input [56:0] input_806;
    input [56:0] input_807;
    input [56:0] input_808;
    input [56:0] input_809;
    input [56:0] input_810;
    input [56:0] input_811;
    input [56:0] input_812;
    input [56:0] input_813;
    input [56:0] input_814;
    input [56:0] input_815;
    input [56:0] input_816;
    input [56:0] input_817;
    input [56:0] input_818;
    input [56:0] input_819;
    input [56:0] input_820;
    input [56:0] input_821;
    input [56:0] input_822;
    input [56:0] input_823;
    input [56:0] input_824;
    input [56:0] input_825;
    input [56:0] input_826;
    input [56:0] input_827;
    input [56:0] input_828;
    input [56:0] input_829;
    input [56:0] input_830;
    input [56:0] input_831;
    input [56:0] input_832;
    input [56:0] input_833;
    input [56:0] input_834;
    input [56:0] input_835;
    input [56:0] input_836;
    input [56:0] input_837;
    input [56:0] input_838;
    input [56:0] input_839;
    input [56:0] input_840;
    input [56:0] input_841;
    input [56:0] input_842;
    input [56:0] input_843;
    input [56:0] input_844;
    input [56:0] input_845;
    input [56:0] input_846;
    input [56:0] input_847;
    input [56:0] input_848;
    input [56:0] input_849;
    input [56:0] input_850;
    input [56:0] input_851;
    input [56:0] input_852;
    input [56:0] input_853;
    input [56:0] input_854;
    input [56:0] input_855;
    input [56:0] input_856;
    input [56:0] input_857;
    input [56:0] input_858;
    input [56:0] input_859;
    input [56:0] input_860;
    input [56:0] input_861;
    input [56:0] input_862;
    input [56:0] input_863;
    input [56:0] input_864;
    input [56:0] input_865;
    input [56:0] input_866;
    input [56:0] input_867;
    input [56:0] input_868;
    input [56:0] input_869;
    input [56:0] input_870;
    input [56:0] input_871;
    input [56:0] input_872;
    input [56:0] input_873;
    input [56:0] input_874;
    input [56:0] input_875;
    input [56:0] input_876;
    input [56:0] input_877;
    input [56:0] input_878;
    input [56:0] input_879;
    input [56:0] input_880;
    input [56:0] input_881;
    input [56:0] input_882;
    input [56:0] input_883;
    input [56:0] input_884;
    input [56:0] input_885;
    input [56:0] input_886;
    input [56:0] input_887;
    input [56:0] input_888;
    input [56:0] input_889;
    input [56:0] input_890;
    input [56:0] input_891;
    input [56:0] input_892;
    input [56:0] input_893;
    input [56:0] input_894;
    input [56:0] input_895;
    input [56:0] input_896;
    input [56:0] input_897;
    input [56:0] input_898;
    input [56:0] input_899;
    input [56:0] input_900;
    input [56:0] input_901;
    input [56:0] input_902;
    input [56:0] input_903;
    input [56:0] input_904;
    input [56:0] input_905;
    input [56:0] input_906;
    input [56:0] input_907;
    input [56:0] input_908;
    input [56:0] input_909;
    input [56:0] input_910;
    input [56:0] input_911;
    input [56:0] input_912;
    input [56:0] input_913;
    input [56:0] input_914;
    input [56:0] input_915;
    input [56:0] input_916;
    input [56:0] input_917;
    input [56:0] input_918;
    input [56:0] input_919;
    input [56:0] input_920;
    input [56:0] input_921;
    input [56:0] input_922;
    input [56:0] input_923;
    input [56:0] input_924;
    input [56:0] input_925;
    input [56:0] input_926;
    input [56:0] input_927;
    input [56:0] input_928;
    input [56:0] input_929;
    input [56:0] input_930;
    input [56:0] input_931;
    input [56:0] input_932;
    input [56:0] input_933;
    input [56:0] input_934;
    input [56:0] input_935;
    input [56:0] input_936;
    input [56:0] input_937;
    input [56:0] input_938;
    input [56:0] input_939;
    input [56:0] input_940;
    input [56:0] input_941;
    input [56:0] input_942;
    input [56:0] input_943;
    input [56:0] input_944;
    input [56:0] input_945;
    input [56:0] input_946;
    input [56:0] input_947;
    input [56:0] input_948;
    input [56:0] input_949;
    input [56:0] input_950;
    input [56:0] input_951;
    input [56:0] input_952;
    input [56:0] input_953;
    input [56:0] input_954;
    input [56:0] input_955;
    input [56:0] input_956;
    input [56:0] input_957;
    input [56:0] input_958;
    input [56:0] input_959;
    input [56:0] input_960;
    input [56:0] input_961;
    input [56:0] input_962;
    input [56:0] input_963;
    input [56:0] input_964;
    input [56:0] input_965;
    input [56:0] input_966;
    input [56:0] input_967;
    input [56:0] input_968;
    input [56:0] input_969;
    input [56:0] input_970;
    input [56:0] input_971;
    input [56:0] input_972;
    input [56:0] input_973;
    input [56:0] input_974;
    input [56:0] input_975;
    input [56:0] input_976;
    input [56:0] input_977;
    input [56:0] input_978;
    input [56:0] input_979;
    input [56:0] input_980;
    input [56:0] input_981;
    input [56:0] input_982;
    input [56:0] input_983;
    input [56:0] input_984;
    input [56:0] input_985;
    input [56:0] input_986;
    input [56:0] input_987;
    input [56:0] input_988;
    input [56:0] input_989;
    input [56:0] input_990;
    input [56:0] input_991;
    input [56:0] input_992;
    input [56:0] input_993;
    input [56:0] input_994;
    input [56:0] input_995;
    input [56:0] input_996;
    input [56:0] input_997;
    input [56:0] input_998;
    input [56:0] input_999;
    input [56:0] input_1000;
    input [56:0] input_1001;
    input [56:0] input_1002;
    input [56:0] input_1003;
    input [56:0] input_1004;
    input [56:0] input_1005;
    input [56:0] input_1006;
    input [56:0] input_1007;
    input [56:0] input_1008;
    input [56:0] input_1009;
    input [56:0] input_1010;
    input [56:0] input_1011;
    input [56:0] input_1012;
    input [56:0] input_1013;
    input [56:0] input_1014;
    input [56:0] input_1015;
    input [56:0] input_1016;
    input [56:0] input_1017;
    input [56:0] input_1018;
    input [56:0] input_1019;
    input [56:0] input_1020;
    input [56:0] input_1021;
    input [56:0] input_1022;
    input [56:0] input_1023;
    input [9:0] sel;
    reg [56:0] result;
  begin
    case (sel)
      10'b0000000000 : begin
        result = input_0;
      end
      10'b0000000001 : begin
        result = input_1;
      end
      10'b0000000010 : begin
        result = input_2;
      end
      10'b0000000011 : begin
        result = input_3;
      end
      10'b0000000100 : begin
        result = input_4;
      end
      10'b0000000101 : begin
        result = input_5;
      end
      10'b0000000110 : begin
        result = input_6;
      end
      10'b0000000111 : begin
        result = input_7;
      end
      10'b0000001000 : begin
        result = input_8;
      end
      10'b0000001001 : begin
        result = input_9;
      end
      10'b0000001010 : begin
        result = input_10;
      end
      10'b0000001011 : begin
        result = input_11;
      end
      10'b0000001100 : begin
        result = input_12;
      end
      10'b0000001101 : begin
        result = input_13;
      end
      10'b0000001110 : begin
        result = input_14;
      end
      10'b0000001111 : begin
        result = input_15;
      end
      10'b0000010000 : begin
        result = input_16;
      end
      10'b0000010001 : begin
        result = input_17;
      end
      10'b0000010010 : begin
        result = input_18;
      end
      10'b0000010011 : begin
        result = input_19;
      end
      10'b0000010100 : begin
        result = input_20;
      end
      10'b0000010101 : begin
        result = input_21;
      end
      10'b0000010110 : begin
        result = input_22;
      end
      10'b0000010111 : begin
        result = input_23;
      end
      10'b0000011000 : begin
        result = input_24;
      end
      10'b0000011001 : begin
        result = input_25;
      end
      10'b0000011010 : begin
        result = input_26;
      end
      10'b0000011011 : begin
        result = input_27;
      end
      10'b0000011100 : begin
        result = input_28;
      end
      10'b0000011101 : begin
        result = input_29;
      end
      10'b0000011110 : begin
        result = input_30;
      end
      10'b0000011111 : begin
        result = input_31;
      end
      10'b0000100000 : begin
        result = input_32;
      end
      10'b0000100001 : begin
        result = input_33;
      end
      10'b0000100010 : begin
        result = input_34;
      end
      10'b0000100011 : begin
        result = input_35;
      end
      10'b0000100100 : begin
        result = input_36;
      end
      10'b0000100101 : begin
        result = input_37;
      end
      10'b0000100110 : begin
        result = input_38;
      end
      10'b0000100111 : begin
        result = input_39;
      end
      10'b0000101000 : begin
        result = input_40;
      end
      10'b0000101001 : begin
        result = input_41;
      end
      10'b0000101010 : begin
        result = input_42;
      end
      10'b0000101011 : begin
        result = input_43;
      end
      10'b0000101100 : begin
        result = input_44;
      end
      10'b0000101101 : begin
        result = input_45;
      end
      10'b0000101110 : begin
        result = input_46;
      end
      10'b0000101111 : begin
        result = input_47;
      end
      10'b0000110000 : begin
        result = input_48;
      end
      10'b0000110001 : begin
        result = input_49;
      end
      10'b0000110010 : begin
        result = input_50;
      end
      10'b0000110011 : begin
        result = input_51;
      end
      10'b0000110100 : begin
        result = input_52;
      end
      10'b0000110101 : begin
        result = input_53;
      end
      10'b0000110110 : begin
        result = input_54;
      end
      10'b0000110111 : begin
        result = input_55;
      end
      10'b0000111000 : begin
        result = input_56;
      end
      10'b0000111001 : begin
        result = input_57;
      end
      10'b0000111010 : begin
        result = input_58;
      end
      10'b0000111011 : begin
        result = input_59;
      end
      10'b0000111100 : begin
        result = input_60;
      end
      10'b0000111101 : begin
        result = input_61;
      end
      10'b0000111110 : begin
        result = input_62;
      end
      10'b0000111111 : begin
        result = input_63;
      end
      10'b0001000000 : begin
        result = input_64;
      end
      10'b0001000001 : begin
        result = input_65;
      end
      10'b0001000010 : begin
        result = input_66;
      end
      10'b0001000011 : begin
        result = input_67;
      end
      10'b0001000100 : begin
        result = input_68;
      end
      10'b0001000101 : begin
        result = input_69;
      end
      10'b0001000110 : begin
        result = input_70;
      end
      10'b0001000111 : begin
        result = input_71;
      end
      10'b0001001000 : begin
        result = input_72;
      end
      10'b0001001001 : begin
        result = input_73;
      end
      10'b0001001010 : begin
        result = input_74;
      end
      10'b0001001011 : begin
        result = input_75;
      end
      10'b0001001100 : begin
        result = input_76;
      end
      10'b0001001101 : begin
        result = input_77;
      end
      10'b0001001110 : begin
        result = input_78;
      end
      10'b0001001111 : begin
        result = input_79;
      end
      10'b0001010000 : begin
        result = input_80;
      end
      10'b0001010001 : begin
        result = input_81;
      end
      10'b0001010010 : begin
        result = input_82;
      end
      10'b0001010011 : begin
        result = input_83;
      end
      10'b0001010100 : begin
        result = input_84;
      end
      10'b0001010101 : begin
        result = input_85;
      end
      10'b0001010110 : begin
        result = input_86;
      end
      10'b0001010111 : begin
        result = input_87;
      end
      10'b0001011000 : begin
        result = input_88;
      end
      10'b0001011001 : begin
        result = input_89;
      end
      10'b0001011010 : begin
        result = input_90;
      end
      10'b0001011011 : begin
        result = input_91;
      end
      10'b0001011100 : begin
        result = input_92;
      end
      10'b0001011101 : begin
        result = input_93;
      end
      10'b0001011110 : begin
        result = input_94;
      end
      10'b0001011111 : begin
        result = input_95;
      end
      10'b0001100000 : begin
        result = input_96;
      end
      10'b0001100001 : begin
        result = input_97;
      end
      10'b0001100010 : begin
        result = input_98;
      end
      10'b0001100011 : begin
        result = input_99;
      end
      10'b0001100100 : begin
        result = input_100;
      end
      10'b0001100101 : begin
        result = input_101;
      end
      10'b0001100110 : begin
        result = input_102;
      end
      10'b0001100111 : begin
        result = input_103;
      end
      10'b0001101000 : begin
        result = input_104;
      end
      10'b0001101001 : begin
        result = input_105;
      end
      10'b0001101010 : begin
        result = input_106;
      end
      10'b0001101011 : begin
        result = input_107;
      end
      10'b0001101100 : begin
        result = input_108;
      end
      10'b0001101101 : begin
        result = input_109;
      end
      10'b0001101110 : begin
        result = input_110;
      end
      10'b0001101111 : begin
        result = input_111;
      end
      10'b0001110000 : begin
        result = input_112;
      end
      10'b0001110001 : begin
        result = input_113;
      end
      10'b0001110010 : begin
        result = input_114;
      end
      10'b0001110011 : begin
        result = input_115;
      end
      10'b0001110100 : begin
        result = input_116;
      end
      10'b0001110101 : begin
        result = input_117;
      end
      10'b0001110110 : begin
        result = input_118;
      end
      10'b0001110111 : begin
        result = input_119;
      end
      10'b0001111000 : begin
        result = input_120;
      end
      10'b0001111001 : begin
        result = input_121;
      end
      10'b0001111010 : begin
        result = input_122;
      end
      10'b0001111011 : begin
        result = input_123;
      end
      10'b0001111100 : begin
        result = input_124;
      end
      10'b0001111101 : begin
        result = input_125;
      end
      10'b0001111110 : begin
        result = input_126;
      end
      10'b0001111111 : begin
        result = input_127;
      end
      10'b0010000000 : begin
        result = input_128;
      end
      10'b0010000001 : begin
        result = input_129;
      end
      10'b0010000010 : begin
        result = input_130;
      end
      10'b0010000011 : begin
        result = input_131;
      end
      10'b0010000100 : begin
        result = input_132;
      end
      10'b0010000101 : begin
        result = input_133;
      end
      10'b0010000110 : begin
        result = input_134;
      end
      10'b0010000111 : begin
        result = input_135;
      end
      10'b0010001000 : begin
        result = input_136;
      end
      10'b0010001001 : begin
        result = input_137;
      end
      10'b0010001010 : begin
        result = input_138;
      end
      10'b0010001011 : begin
        result = input_139;
      end
      10'b0010001100 : begin
        result = input_140;
      end
      10'b0010001101 : begin
        result = input_141;
      end
      10'b0010001110 : begin
        result = input_142;
      end
      10'b0010001111 : begin
        result = input_143;
      end
      10'b0010010000 : begin
        result = input_144;
      end
      10'b0010010001 : begin
        result = input_145;
      end
      10'b0010010010 : begin
        result = input_146;
      end
      10'b0010010011 : begin
        result = input_147;
      end
      10'b0010010100 : begin
        result = input_148;
      end
      10'b0010010101 : begin
        result = input_149;
      end
      10'b0010010110 : begin
        result = input_150;
      end
      10'b0010010111 : begin
        result = input_151;
      end
      10'b0010011000 : begin
        result = input_152;
      end
      10'b0010011001 : begin
        result = input_153;
      end
      10'b0010011010 : begin
        result = input_154;
      end
      10'b0010011011 : begin
        result = input_155;
      end
      10'b0010011100 : begin
        result = input_156;
      end
      10'b0010011101 : begin
        result = input_157;
      end
      10'b0010011110 : begin
        result = input_158;
      end
      10'b0010011111 : begin
        result = input_159;
      end
      10'b0010100000 : begin
        result = input_160;
      end
      10'b0010100001 : begin
        result = input_161;
      end
      10'b0010100010 : begin
        result = input_162;
      end
      10'b0010100011 : begin
        result = input_163;
      end
      10'b0010100100 : begin
        result = input_164;
      end
      10'b0010100101 : begin
        result = input_165;
      end
      10'b0010100110 : begin
        result = input_166;
      end
      10'b0010100111 : begin
        result = input_167;
      end
      10'b0010101000 : begin
        result = input_168;
      end
      10'b0010101001 : begin
        result = input_169;
      end
      10'b0010101010 : begin
        result = input_170;
      end
      10'b0010101011 : begin
        result = input_171;
      end
      10'b0010101100 : begin
        result = input_172;
      end
      10'b0010101101 : begin
        result = input_173;
      end
      10'b0010101110 : begin
        result = input_174;
      end
      10'b0010101111 : begin
        result = input_175;
      end
      10'b0010110000 : begin
        result = input_176;
      end
      10'b0010110001 : begin
        result = input_177;
      end
      10'b0010110010 : begin
        result = input_178;
      end
      10'b0010110011 : begin
        result = input_179;
      end
      10'b0010110100 : begin
        result = input_180;
      end
      10'b0010110101 : begin
        result = input_181;
      end
      10'b0010110110 : begin
        result = input_182;
      end
      10'b0010110111 : begin
        result = input_183;
      end
      10'b0010111000 : begin
        result = input_184;
      end
      10'b0010111001 : begin
        result = input_185;
      end
      10'b0010111010 : begin
        result = input_186;
      end
      10'b0010111011 : begin
        result = input_187;
      end
      10'b0010111100 : begin
        result = input_188;
      end
      10'b0010111101 : begin
        result = input_189;
      end
      10'b0010111110 : begin
        result = input_190;
      end
      10'b0010111111 : begin
        result = input_191;
      end
      10'b0011000000 : begin
        result = input_192;
      end
      10'b0011000001 : begin
        result = input_193;
      end
      10'b0011000010 : begin
        result = input_194;
      end
      10'b0011000011 : begin
        result = input_195;
      end
      10'b0011000100 : begin
        result = input_196;
      end
      10'b0011000101 : begin
        result = input_197;
      end
      10'b0011000110 : begin
        result = input_198;
      end
      10'b0011000111 : begin
        result = input_199;
      end
      10'b0011001000 : begin
        result = input_200;
      end
      10'b0011001001 : begin
        result = input_201;
      end
      10'b0011001010 : begin
        result = input_202;
      end
      10'b0011001011 : begin
        result = input_203;
      end
      10'b0011001100 : begin
        result = input_204;
      end
      10'b0011001101 : begin
        result = input_205;
      end
      10'b0011001110 : begin
        result = input_206;
      end
      10'b0011001111 : begin
        result = input_207;
      end
      10'b0011010000 : begin
        result = input_208;
      end
      10'b0011010001 : begin
        result = input_209;
      end
      10'b0011010010 : begin
        result = input_210;
      end
      10'b0011010011 : begin
        result = input_211;
      end
      10'b0011010100 : begin
        result = input_212;
      end
      10'b0011010101 : begin
        result = input_213;
      end
      10'b0011010110 : begin
        result = input_214;
      end
      10'b0011010111 : begin
        result = input_215;
      end
      10'b0011011000 : begin
        result = input_216;
      end
      10'b0011011001 : begin
        result = input_217;
      end
      10'b0011011010 : begin
        result = input_218;
      end
      10'b0011011011 : begin
        result = input_219;
      end
      10'b0011011100 : begin
        result = input_220;
      end
      10'b0011011101 : begin
        result = input_221;
      end
      10'b0011011110 : begin
        result = input_222;
      end
      10'b0011011111 : begin
        result = input_223;
      end
      10'b0011100000 : begin
        result = input_224;
      end
      10'b0011100001 : begin
        result = input_225;
      end
      10'b0011100010 : begin
        result = input_226;
      end
      10'b0011100011 : begin
        result = input_227;
      end
      10'b0011100100 : begin
        result = input_228;
      end
      10'b0011100101 : begin
        result = input_229;
      end
      10'b0011100110 : begin
        result = input_230;
      end
      10'b0011100111 : begin
        result = input_231;
      end
      10'b0011101000 : begin
        result = input_232;
      end
      10'b0011101001 : begin
        result = input_233;
      end
      10'b0011101010 : begin
        result = input_234;
      end
      10'b0011101011 : begin
        result = input_235;
      end
      10'b0011101100 : begin
        result = input_236;
      end
      10'b0011101101 : begin
        result = input_237;
      end
      10'b0011101110 : begin
        result = input_238;
      end
      10'b0011101111 : begin
        result = input_239;
      end
      10'b0011110000 : begin
        result = input_240;
      end
      10'b0011110001 : begin
        result = input_241;
      end
      10'b0011110010 : begin
        result = input_242;
      end
      10'b0011110011 : begin
        result = input_243;
      end
      10'b0011110100 : begin
        result = input_244;
      end
      10'b0011110101 : begin
        result = input_245;
      end
      10'b0011110110 : begin
        result = input_246;
      end
      10'b0011110111 : begin
        result = input_247;
      end
      10'b0011111000 : begin
        result = input_248;
      end
      10'b0011111001 : begin
        result = input_249;
      end
      10'b0011111010 : begin
        result = input_250;
      end
      10'b0011111011 : begin
        result = input_251;
      end
      10'b0011111100 : begin
        result = input_252;
      end
      10'b0011111101 : begin
        result = input_253;
      end
      10'b0011111110 : begin
        result = input_254;
      end
      10'b0011111111 : begin
        result = input_255;
      end
      10'b0100000000 : begin
        result = input_256;
      end
      10'b0100000001 : begin
        result = input_257;
      end
      10'b0100000010 : begin
        result = input_258;
      end
      10'b0100000011 : begin
        result = input_259;
      end
      10'b0100000100 : begin
        result = input_260;
      end
      10'b0100000101 : begin
        result = input_261;
      end
      10'b0100000110 : begin
        result = input_262;
      end
      10'b0100000111 : begin
        result = input_263;
      end
      10'b0100001000 : begin
        result = input_264;
      end
      10'b0100001001 : begin
        result = input_265;
      end
      10'b0100001010 : begin
        result = input_266;
      end
      10'b0100001011 : begin
        result = input_267;
      end
      10'b0100001100 : begin
        result = input_268;
      end
      10'b0100001101 : begin
        result = input_269;
      end
      10'b0100001110 : begin
        result = input_270;
      end
      10'b0100001111 : begin
        result = input_271;
      end
      10'b0100010000 : begin
        result = input_272;
      end
      10'b0100010001 : begin
        result = input_273;
      end
      10'b0100010010 : begin
        result = input_274;
      end
      10'b0100010011 : begin
        result = input_275;
      end
      10'b0100010100 : begin
        result = input_276;
      end
      10'b0100010101 : begin
        result = input_277;
      end
      10'b0100010110 : begin
        result = input_278;
      end
      10'b0100010111 : begin
        result = input_279;
      end
      10'b0100011000 : begin
        result = input_280;
      end
      10'b0100011001 : begin
        result = input_281;
      end
      10'b0100011010 : begin
        result = input_282;
      end
      10'b0100011011 : begin
        result = input_283;
      end
      10'b0100011100 : begin
        result = input_284;
      end
      10'b0100011101 : begin
        result = input_285;
      end
      10'b0100011110 : begin
        result = input_286;
      end
      10'b0100011111 : begin
        result = input_287;
      end
      10'b0100100000 : begin
        result = input_288;
      end
      10'b0100100001 : begin
        result = input_289;
      end
      10'b0100100010 : begin
        result = input_290;
      end
      10'b0100100011 : begin
        result = input_291;
      end
      10'b0100100100 : begin
        result = input_292;
      end
      10'b0100100101 : begin
        result = input_293;
      end
      10'b0100100110 : begin
        result = input_294;
      end
      10'b0100100111 : begin
        result = input_295;
      end
      10'b0100101000 : begin
        result = input_296;
      end
      10'b0100101001 : begin
        result = input_297;
      end
      10'b0100101010 : begin
        result = input_298;
      end
      10'b0100101011 : begin
        result = input_299;
      end
      10'b0100101100 : begin
        result = input_300;
      end
      10'b0100101101 : begin
        result = input_301;
      end
      10'b0100101110 : begin
        result = input_302;
      end
      10'b0100101111 : begin
        result = input_303;
      end
      10'b0100110000 : begin
        result = input_304;
      end
      10'b0100110001 : begin
        result = input_305;
      end
      10'b0100110010 : begin
        result = input_306;
      end
      10'b0100110011 : begin
        result = input_307;
      end
      10'b0100110100 : begin
        result = input_308;
      end
      10'b0100110101 : begin
        result = input_309;
      end
      10'b0100110110 : begin
        result = input_310;
      end
      10'b0100110111 : begin
        result = input_311;
      end
      10'b0100111000 : begin
        result = input_312;
      end
      10'b0100111001 : begin
        result = input_313;
      end
      10'b0100111010 : begin
        result = input_314;
      end
      10'b0100111011 : begin
        result = input_315;
      end
      10'b0100111100 : begin
        result = input_316;
      end
      10'b0100111101 : begin
        result = input_317;
      end
      10'b0100111110 : begin
        result = input_318;
      end
      10'b0100111111 : begin
        result = input_319;
      end
      10'b0101000000 : begin
        result = input_320;
      end
      10'b0101000001 : begin
        result = input_321;
      end
      10'b0101000010 : begin
        result = input_322;
      end
      10'b0101000011 : begin
        result = input_323;
      end
      10'b0101000100 : begin
        result = input_324;
      end
      10'b0101000101 : begin
        result = input_325;
      end
      10'b0101000110 : begin
        result = input_326;
      end
      10'b0101000111 : begin
        result = input_327;
      end
      10'b0101001000 : begin
        result = input_328;
      end
      10'b0101001001 : begin
        result = input_329;
      end
      10'b0101001010 : begin
        result = input_330;
      end
      10'b0101001011 : begin
        result = input_331;
      end
      10'b0101001100 : begin
        result = input_332;
      end
      10'b0101001101 : begin
        result = input_333;
      end
      10'b0101001110 : begin
        result = input_334;
      end
      10'b0101001111 : begin
        result = input_335;
      end
      10'b0101010000 : begin
        result = input_336;
      end
      10'b0101010001 : begin
        result = input_337;
      end
      10'b0101010010 : begin
        result = input_338;
      end
      10'b0101010011 : begin
        result = input_339;
      end
      10'b0101010100 : begin
        result = input_340;
      end
      10'b0101010101 : begin
        result = input_341;
      end
      10'b0101010110 : begin
        result = input_342;
      end
      10'b0101010111 : begin
        result = input_343;
      end
      10'b0101011000 : begin
        result = input_344;
      end
      10'b0101011001 : begin
        result = input_345;
      end
      10'b0101011010 : begin
        result = input_346;
      end
      10'b0101011011 : begin
        result = input_347;
      end
      10'b0101011100 : begin
        result = input_348;
      end
      10'b0101011101 : begin
        result = input_349;
      end
      10'b0101011110 : begin
        result = input_350;
      end
      10'b0101011111 : begin
        result = input_351;
      end
      10'b0101100000 : begin
        result = input_352;
      end
      10'b0101100001 : begin
        result = input_353;
      end
      10'b0101100010 : begin
        result = input_354;
      end
      10'b0101100011 : begin
        result = input_355;
      end
      10'b0101100100 : begin
        result = input_356;
      end
      10'b0101100101 : begin
        result = input_357;
      end
      10'b0101100110 : begin
        result = input_358;
      end
      10'b0101100111 : begin
        result = input_359;
      end
      10'b0101101000 : begin
        result = input_360;
      end
      10'b0101101001 : begin
        result = input_361;
      end
      10'b0101101010 : begin
        result = input_362;
      end
      10'b0101101011 : begin
        result = input_363;
      end
      10'b0101101100 : begin
        result = input_364;
      end
      10'b0101101101 : begin
        result = input_365;
      end
      10'b0101101110 : begin
        result = input_366;
      end
      10'b0101101111 : begin
        result = input_367;
      end
      10'b0101110000 : begin
        result = input_368;
      end
      10'b0101110001 : begin
        result = input_369;
      end
      10'b0101110010 : begin
        result = input_370;
      end
      10'b0101110011 : begin
        result = input_371;
      end
      10'b0101110100 : begin
        result = input_372;
      end
      10'b0101110101 : begin
        result = input_373;
      end
      10'b0101110110 : begin
        result = input_374;
      end
      10'b0101110111 : begin
        result = input_375;
      end
      10'b0101111000 : begin
        result = input_376;
      end
      10'b0101111001 : begin
        result = input_377;
      end
      10'b0101111010 : begin
        result = input_378;
      end
      10'b0101111011 : begin
        result = input_379;
      end
      10'b0101111100 : begin
        result = input_380;
      end
      10'b0101111101 : begin
        result = input_381;
      end
      10'b0101111110 : begin
        result = input_382;
      end
      10'b0101111111 : begin
        result = input_383;
      end
      10'b0110000000 : begin
        result = input_384;
      end
      10'b0110000001 : begin
        result = input_385;
      end
      10'b0110000010 : begin
        result = input_386;
      end
      10'b0110000011 : begin
        result = input_387;
      end
      10'b0110000100 : begin
        result = input_388;
      end
      10'b0110000101 : begin
        result = input_389;
      end
      10'b0110000110 : begin
        result = input_390;
      end
      10'b0110000111 : begin
        result = input_391;
      end
      10'b0110001000 : begin
        result = input_392;
      end
      10'b0110001001 : begin
        result = input_393;
      end
      10'b0110001010 : begin
        result = input_394;
      end
      10'b0110001011 : begin
        result = input_395;
      end
      10'b0110001100 : begin
        result = input_396;
      end
      10'b0110001101 : begin
        result = input_397;
      end
      10'b0110001110 : begin
        result = input_398;
      end
      10'b0110001111 : begin
        result = input_399;
      end
      10'b0110010000 : begin
        result = input_400;
      end
      10'b0110010001 : begin
        result = input_401;
      end
      10'b0110010010 : begin
        result = input_402;
      end
      10'b0110010011 : begin
        result = input_403;
      end
      10'b0110010100 : begin
        result = input_404;
      end
      10'b0110010101 : begin
        result = input_405;
      end
      10'b0110010110 : begin
        result = input_406;
      end
      10'b0110010111 : begin
        result = input_407;
      end
      10'b0110011000 : begin
        result = input_408;
      end
      10'b0110011001 : begin
        result = input_409;
      end
      10'b0110011010 : begin
        result = input_410;
      end
      10'b0110011011 : begin
        result = input_411;
      end
      10'b0110011100 : begin
        result = input_412;
      end
      10'b0110011101 : begin
        result = input_413;
      end
      10'b0110011110 : begin
        result = input_414;
      end
      10'b0110011111 : begin
        result = input_415;
      end
      10'b0110100000 : begin
        result = input_416;
      end
      10'b0110100001 : begin
        result = input_417;
      end
      10'b0110100010 : begin
        result = input_418;
      end
      10'b0110100011 : begin
        result = input_419;
      end
      10'b0110100100 : begin
        result = input_420;
      end
      10'b0110100101 : begin
        result = input_421;
      end
      10'b0110100110 : begin
        result = input_422;
      end
      10'b0110100111 : begin
        result = input_423;
      end
      10'b0110101000 : begin
        result = input_424;
      end
      10'b0110101001 : begin
        result = input_425;
      end
      10'b0110101010 : begin
        result = input_426;
      end
      10'b0110101011 : begin
        result = input_427;
      end
      10'b0110101100 : begin
        result = input_428;
      end
      10'b0110101101 : begin
        result = input_429;
      end
      10'b0110101110 : begin
        result = input_430;
      end
      10'b0110101111 : begin
        result = input_431;
      end
      10'b0110110000 : begin
        result = input_432;
      end
      10'b0110110001 : begin
        result = input_433;
      end
      10'b0110110010 : begin
        result = input_434;
      end
      10'b0110110011 : begin
        result = input_435;
      end
      10'b0110110100 : begin
        result = input_436;
      end
      10'b0110110101 : begin
        result = input_437;
      end
      10'b0110110110 : begin
        result = input_438;
      end
      10'b0110110111 : begin
        result = input_439;
      end
      10'b0110111000 : begin
        result = input_440;
      end
      10'b0110111001 : begin
        result = input_441;
      end
      10'b0110111010 : begin
        result = input_442;
      end
      10'b0110111011 : begin
        result = input_443;
      end
      10'b0110111100 : begin
        result = input_444;
      end
      10'b0110111101 : begin
        result = input_445;
      end
      10'b0110111110 : begin
        result = input_446;
      end
      10'b0110111111 : begin
        result = input_447;
      end
      10'b0111000000 : begin
        result = input_448;
      end
      10'b0111000001 : begin
        result = input_449;
      end
      10'b0111000010 : begin
        result = input_450;
      end
      10'b0111000011 : begin
        result = input_451;
      end
      10'b0111000100 : begin
        result = input_452;
      end
      10'b0111000101 : begin
        result = input_453;
      end
      10'b0111000110 : begin
        result = input_454;
      end
      10'b0111000111 : begin
        result = input_455;
      end
      10'b0111001000 : begin
        result = input_456;
      end
      10'b0111001001 : begin
        result = input_457;
      end
      10'b0111001010 : begin
        result = input_458;
      end
      10'b0111001011 : begin
        result = input_459;
      end
      10'b0111001100 : begin
        result = input_460;
      end
      10'b0111001101 : begin
        result = input_461;
      end
      10'b0111001110 : begin
        result = input_462;
      end
      10'b0111001111 : begin
        result = input_463;
      end
      10'b0111010000 : begin
        result = input_464;
      end
      10'b0111010001 : begin
        result = input_465;
      end
      10'b0111010010 : begin
        result = input_466;
      end
      10'b0111010011 : begin
        result = input_467;
      end
      10'b0111010100 : begin
        result = input_468;
      end
      10'b0111010101 : begin
        result = input_469;
      end
      10'b0111010110 : begin
        result = input_470;
      end
      10'b0111010111 : begin
        result = input_471;
      end
      10'b0111011000 : begin
        result = input_472;
      end
      10'b0111011001 : begin
        result = input_473;
      end
      10'b0111011010 : begin
        result = input_474;
      end
      10'b0111011011 : begin
        result = input_475;
      end
      10'b0111011100 : begin
        result = input_476;
      end
      10'b0111011101 : begin
        result = input_477;
      end
      10'b0111011110 : begin
        result = input_478;
      end
      10'b0111011111 : begin
        result = input_479;
      end
      10'b0111100000 : begin
        result = input_480;
      end
      10'b0111100001 : begin
        result = input_481;
      end
      10'b0111100010 : begin
        result = input_482;
      end
      10'b0111100011 : begin
        result = input_483;
      end
      10'b0111100100 : begin
        result = input_484;
      end
      10'b0111100101 : begin
        result = input_485;
      end
      10'b0111100110 : begin
        result = input_486;
      end
      10'b0111100111 : begin
        result = input_487;
      end
      10'b0111101000 : begin
        result = input_488;
      end
      10'b0111101001 : begin
        result = input_489;
      end
      10'b0111101010 : begin
        result = input_490;
      end
      10'b0111101011 : begin
        result = input_491;
      end
      10'b0111101100 : begin
        result = input_492;
      end
      10'b0111101101 : begin
        result = input_493;
      end
      10'b0111101110 : begin
        result = input_494;
      end
      10'b0111101111 : begin
        result = input_495;
      end
      10'b0111110000 : begin
        result = input_496;
      end
      10'b0111110001 : begin
        result = input_497;
      end
      10'b0111110010 : begin
        result = input_498;
      end
      10'b0111110011 : begin
        result = input_499;
      end
      10'b0111110100 : begin
        result = input_500;
      end
      10'b0111110101 : begin
        result = input_501;
      end
      10'b0111110110 : begin
        result = input_502;
      end
      10'b0111110111 : begin
        result = input_503;
      end
      10'b0111111000 : begin
        result = input_504;
      end
      10'b0111111001 : begin
        result = input_505;
      end
      10'b0111111010 : begin
        result = input_506;
      end
      10'b0111111011 : begin
        result = input_507;
      end
      10'b0111111100 : begin
        result = input_508;
      end
      10'b0111111101 : begin
        result = input_509;
      end
      10'b0111111110 : begin
        result = input_510;
      end
      10'b0111111111 : begin
        result = input_511;
      end
      10'b1000000000 : begin
        result = input_512;
      end
      10'b1000000001 : begin
        result = input_513;
      end
      10'b1000000010 : begin
        result = input_514;
      end
      10'b1000000011 : begin
        result = input_515;
      end
      10'b1000000100 : begin
        result = input_516;
      end
      10'b1000000101 : begin
        result = input_517;
      end
      10'b1000000110 : begin
        result = input_518;
      end
      10'b1000000111 : begin
        result = input_519;
      end
      10'b1000001000 : begin
        result = input_520;
      end
      10'b1000001001 : begin
        result = input_521;
      end
      10'b1000001010 : begin
        result = input_522;
      end
      10'b1000001011 : begin
        result = input_523;
      end
      10'b1000001100 : begin
        result = input_524;
      end
      10'b1000001101 : begin
        result = input_525;
      end
      10'b1000001110 : begin
        result = input_526;
      end
      10'b1000001111 : begin
        result = input_527;
      end
      10'b1000010000 : begin
        result = input_528;
      end
      10'b1000010001 : begin
        result = input_529;
      end
      10'b1000010010 : begin
        result = input_530;
      end
      10'b1000010011 : begin
        result = input_531;
      end
      10'b1000010100 : begin
        result = input_532;
      end
      10'b1000010101 : begin
        result = input_533;
      end
      10'b1000010110 : begin
        result = input_534;
      end
      10'b1000010111 : begin
        result = input_535;
      end
      10'b1000011000 : begin
        result = input_536;
      end
      10'b1000011001 : begin
        result = input_537;
      end
      10'b1000011010 : begin
        result = input_538;
      end
      10'b1000011011 : begin
        result = input_539;
      end
      10'b1000011100 : begin
        result = input_540;
      end
      10'b1000011101 : begin
        result = input_541;
      end
      10'b1000011110 : begin
        result = input_542;
      end
      10'b1000011111 : begin
        result = input_543;
      end
      10'b1000100000 : begin
        result = input_544;
      end
      10'b1000100001 : begin
        result = input_545;
      end
      10'b1000100010 : begin
        result = input_546;
      end
      10'b1000100011 : begin
        result = input_547;
      end
      10'b1000100100 : begin
        result = input_548;
      end
      10'b1000100101 : begin
        result = input_549;
      end
      10'b1000100110 : begin
        result = input_550;
      end
      10'b1000100111 : begin
        result = input_551;
      end
      10'b1000101000 : begin
        result = input_552;
      end
      10'b1000101001 : begin
        result = input_553;
      end
      10'b1000101010 : begin
        result = input_554;
      end
      10'b1000101011 : begin
        result = input_555;
      end
      10'b1000101100 : begin
        result = input_556;
      end
      10'b1000101101 : begin
        result = input_557;
      end
      10'b1000101110 : begin
        result = input_558;
      end
      10'b1000101111 : begin
        result = input_559;
      end
      10'b1000110000 : begin
        result = input_560;
      end
      10'b1000110001 : begin
        result = input_561;
      end
      10'b1000110010 : begin
        result = input_562;
      end
      10'b1000110011 : begin
        result = input_563;
      end
      10'b1000110100 : begin
        result = input_564;
      end
      10'b1000110101 : begin
        result = input_565;
      end
      10'b1000110110 : begin
        result = input_566;
      end
      10'b1000110111 : begin
        result = input_567;
      end
      10'b1000111000 : begin
        result = input_568;
      end
      10'b1000111001 : begin
        result = input_569;
      end
      10'b1000111010 : begin
        result = input_570;
      end
      10'b1000111011 : begin
        result = input_571;
      end
      10'b1000111100 : begin
        result = input_572;
      end
      10'b1000111101 : begin
        result = input_573;
      end
      10'b1000111110 : begin
        result = input_574;
      end
      10'b1000111111 : begin
        result = input_575;
      end
      10'b1001000000 : begin
        result = input_576;
      end
      10'b1001000001 : begin
        result = input_577;
      end
      10'b1001000010 : begin
        result = input_578;
      end
      10'b1001000011 : begin
        result = input_579;
      end
      10'b1001000100 : begin
        result = input_580;
      end
      10'b1001000101 : begin
        result = input_581;
      end
      10'b1001000110 : begin
        result = input_582;
      end
      10'b1001000111 : begin
        result = input_583;
      end
      10'b1001001000 : begin
        result = input_584;
      end
      10'b1001001001 : begin
        result = input_585;
      end
      10'b1001001010 : begin
        result = input_586;
      end
      10'b1001001011 : begin
        result = input_587;
      end
      10'b1001001100 : begin
        result = input_588;
      end
      10'b1001001101 : begin
        result = input_589;
      end
      10'b1001001110 : begin
        result = input_590;
      end
      10'b1001001111 : begin
        result = input_591;
      end
      10'b1001010000 : begin
        result = input_592;
      end
      10'b1001010001 : begin
        result = input_593;
      end
      10'b1001010010 : begin
        result = input_594;
      end
      10'b1001010011 : begin
        result = input_595;
      end
      10'b1001010100 : begin
        result = input_596;
      end
      10'b1001010101 : begin
        result = input_597;
      end
      10'b1001010110 : begin
        result = input_598;
      end
      10'b1001010111 : begin
        result = input_599;
      end
      10'b1001011000 : begin
        result = input_600;
      end
      10'b1001011001 : begin
        result = input_601;
      end
      10'b1001011010 : begin
        result = input_602;
      end
      10'b1001011011 : begin
        result = input_603;
      end
      10'b1001011100 : begin
        result = input_604;
      end
      10'b1001011101 : begin
        result = input_605;
      end
      10'b1001011110 : begin
        result = input_606;
      end
      10'b1001011111 : begin
        result = input_607;
      end
      10'b1001100000 : begin
        result = input_608;
      end
      10'b1001100001 : begin
        result = input_609;
      end
      10'b1001100010 : begin
        result = input_610;
      end
      10'b1001100011 : begin
        result = input_611;
      end
      10'b1001100100 : begin
        result = input_612;
      end
      10'b1001100101 : begin
        result = input_613;
      end
      10'b1001100110 : begin
        result = input_614;
      end
      10'b1001100111 : begin
        result = input_615;
      end
      10'b1001101000 : begin
        result = input_616;
      end
      10'b1001101001 : begin
        result = input_617;
      end
      10'b1001101010 : begin
        result = input_618;
      end
      10'b1001101011 : begin
        result = input_619;
      end
      10'b1001101100 : begin
        result = input_620;
      end
      10'b1001101101 : begin
        result = input_621;
      end
      10'b1001101110 : begin
        result = input_622;
      end
      10'b1001101111 : begin
        result = input_623;
      end
      10'b1001110000 : begin
        result = input_624;
      end
      10'b1001110001 : begin
        result = input_625;
      end
      10'b1001110010 : begin
        result = input_626;
      end
      10'b1001110011 : begin
        result = input_627;
      end
      10'b1001110100 : begin
        result = input_628;
      end
      10'b1001110101 : begin
        result = input_629;
      end
      10'b1001110110 : begin
        result = input_630;
      end
      10'b1001110111 : begin
        result = input_631;
      end
      10'b1001111000 : begin
        result = input_632;
      end
      10'b1001111001 : begin
        result = input_633;
      end
      10'b1001111010 : begin
        result = input_634;
      end
      10'b1001111011 : begin
        result = input_635;
      end
      10'b1001111100 : begin
        result = input_636;
      end
      10'b1001111101 : begin
        result = input_637;
      end
      10'b1001111110 : begin
        result = input_638;
      end
      10'b1001111111 : begin
        result = input_639;
      end
      10'b1010000000 : begin
        result = input_640;
      end
      10'b1010000001 : begin
        result = input_641;
      end
      10'b1010000010 : begin
        result = input_642;
      end
      10'b1010000011 : begin
        result = input_643;
      end
      10'b1010000100 : begin
        result = input_644;
      end
      10'b1010000101 : begin
        result = input_645;
      end
      10'b1010000110 : begin
        result = input_646;
      end
      10'b1010000111 : begin
        result = input_647;
      end
      10'b1010001000 : begin
        result = input_648;
      end
      10'b1010001001 : begin
        result = input_649;
      end
      10'b1010001010 : begin
        result = input_650;
      end
      10'b1010001011 : begin
        result = input_651;
      end
      10'b1010001100 : begin
        result = input_652;
      end
      10'b1010001101 : begin
        result = input_653;
      end
      10'b1010001110 : begin
        result = input_654;
      end
      10'b1010001111 : begin
        result = input_655;
      end
      10'b1010010000 : begin
        result = input_656;
      end
      10'b1010010001 : begin
        result = input_657;
      end
      10'b1010010010 : begin
        result = input_658;
      end
      10'b1010010011 : begin
        result = input_659;
      end
      10'b1010010100 : begin
        result = input_660;
      end
      10'b1010010101 : begin
        result = input_661;
      end
      10'b1010010110 : begin
        result = input_662;
      end
      10'b1010010111 : begin
        result = input_663;
      end
      10'b1010011000 : begin
        result = input_664;
      end
      10'b1010011001 : begin
        result = input_665;
      end
      10'b1010011010 : begin
        result = input_666;
      end
      10'b1010011011 : begin
        result = input_667;
      end
      10'b1010011100 : begin
        result = input_668;
      end
      10'b1010011101 : begin
        result = input_669;
      end
      10'b1010011110 : begin
        result = input_670;
      end
      10'b1010011111 : begin
        result = input_671;
      end
      10'b1010100000 : begin
        result = input_672;
      end
      10'b1010100001 : begin
        result = input_673;
      end
      10'b1010100010 : begin
        result = input_674;
      end
      10'b1010100011 : begin
        result = input_675;
      end
      10'b1010100100 : begin
        result = input_676;
      end
      10'b1010100101 : begin
        result = input_677;
      end
      10'b1010100110 : begin
        result = input_678;
      end
      10'b1010100111 : begin
        result = input_679;
      end
      10'b1010101000 : begin
        result = input_680;
      end
      10'b1010101001 : begin
        result = input_681;
      end
      10'b1010101010 : begin
        result = input_682;
      end
      10'b1010101011 : begin
        result = input_683;
      end
      10'b1010101100 : begin
        result = input_684;
      end
      10'b1010101101 : begin
        result = input_685;
      end
      10'b1010101110 : begin
        result = input_686;
      end
      10'b1010101111 : begin
        result = input_687;
      end
      10'b1010110000 : begin
        result = input_688;
      end
      10'b1010110001 : begin
        result = input_689;
      end
      10'b1010110010 : begin
        result = input_690;
      end
      10'b1010110011 : begin
        result = input_691;
      end
      10'b1010110100 : begin
        result = input_692;
      end
      10'b1010110101 : begin
        result = input_693;
      end
      10'b1010110110 : begin
        result = input_694;
      end
      10'b1010110111 : begin
        result = input_695;
      end
      10'b1010111000 : begin
        result = input_696;
      end
      10'b1010111001 : begin
        result = input_697;
      end
      10'b1010111010 : begin
        result = input_698;
      end
      10'b1010111011 : begin
        result = input_699;
      end
      10'b1010111100 : begin
        result = input_700;
      end
      10'b1010111101 : begin
        result = input_701;
      end
      10'b1010111110 : begin
        result = input_702;
      end
      10'b1010111111 : begin
        result = input_703;
      end
      10'b1011000000 : begin
        result = input_704;
      end
      10'b1011000001 : begin
        result = input_705;
      end
      10'b1011000010 : begin
        result = input_706;
      end
      10'b1011000011 : begin
        result = input_707;
      end
      10'b1011000100 : begin
        result = input_708;
      end
      10'b1011000101 : begin
        result = input_709;
      end
      10'b1011000110 : begin
        result = input_710;
      end
      10'b1011000111 : begin
        result = input_711;
      end
      10'b1011001000 : begin
        result = input_712;
      end
      10'b1011001001 : begin
        result = input_713;
      end
      10'b1011001010 : begin
        result = input_714;
      end
      10'b1011001011 : begin
        result = input_715;
      end
      10'b1011001100 : begin
        result = input_716;
      end
      10'b1011001101 : begin
        result = input_717;
      end
      10'b1011001110 : begin
        result = input_718;
      end
      10'b1011001111 : begin
        result = input_719;
      end
      10'b1011010000 : begin
        result = input_720;
      end
      10'b1011010001 : begin
        result = input_721;
      end
      10'b1011010010 : begin
        result = input_722;
      end
      10'b1011010011 : begin
        result = input_723;
      end
      10'b1011010100 : begin
        result = input_724;
      end
      10'b1011010101 : begin
        result = input_725;
      end
      10'b1011010110 : begin
        result = input_726;
      end
      10'b1011010111 : begin
        result = input_727;
      end
      10'b1011011000 : begin
        result = input_728;
      end
      10'b1011011001 : begin
        result = input_729;
      end
      10'b1011011010 : begin
        result = input_730;
      end
      10'b1011011011 : begin
        result = input_731;
      end
      10'b1011011100 : begin
        result = input_732;
      end
      10'b1011011101 : begin
        result = input_733;
      end
      10'b1011011110 : begin
        result = input_734;
      end
      10'b1011011111 : begin
        result = input_735;
      end
      10'b1011100000 : begin
        result = input_736;
      end
      10'b1011100001 : begin
        result = input_737;
      end
      10'b1011100010 : begin
        result = input_738;
      end
      10'b1011100011 : begin
        result = input_739;
      end
      10'b1011100100 : begin
        result = input_740;
      end
      10'b1011100101 : begin
        result = input_741;
      end
      10'b1011100110 : begin
        result = input_742;
      end
      10'b1011100111 : begin
        result = input_743;
      end
      10'b1011101000 : begin
        result = input_744;
      end
      10'b1011101001 : begin
        result = input_745;
      end
      10'b1011101010 : begin
        result = input_746;
      end
      10'b1011101011 : begin
        result = input_747;
      end
      10'b1011101100 : begin
        result = input_748;
      end
      10'b1011101101 : begin
        result = input_749;
      end
      10'b1011101110 : begin
        result = input_750;
      end
      10'b1011101111 : begin
        result = input_751;
      end
      10'b1011110000 : begin
        result = input_752;
      end
      10'b1011110001 : begin
        result = input_753;
      end
      10'b1011110010 : begin
        result = input_754;
      end
      10'b1011110011 : begin
        result = input_755;
      end
      10'b1011110100 : begin
        result = input_756;
      end
      10'b1011110101 : begin
        result = input_757;
      end
      10'b1011110110 : begin
        result = input_758;
      end
      10'b1011110111 : begin
        result = input_759;
      end
      10'b1011111000 : begin
        result = input_760;
      end
      10'b1011111001 : begin
        result = input_761;
      end
      10'b1011111010 : begin
        result = input_762;
      end
      10'b1011111011 : begin
        result = input_763;
      end
      10'b1011111100 : begin
        result = input_764;
      end
      10'b1011111101 : begin
        result = input_765;
      end
      10'b1011111110 : begin
        result = input_766;
      end
      10'b1011111111 : begin
        result = input_767;
      end
      10'b1100000000 : begin
        result = input_768;
      end
      10'b1100000001 : begin
        result = input_769;
      end
      10'b1100000010 : begin
        result = input_770;
      end
      10'b1100000011 : begin
        result = input_771;
      end
      10'b1100000100 : begin
        result = input_772;
      end
      10'b1100000101 : begin
        result = input_773;
      end
      10'b1100000110 : begin
        result = input_774;
      end
      10'b1100000111 : begin
        result = input_775;
      end
      10'b1100001000 : begin
        result = input_776;
      end
      10'b1100001001 : begin
        result = input_777;
      end
      10'b1100001010 : begin
        result = input_778;
      end
      10'b1100001011 : begin
        result = input_779;
      end
      10'b1100001100 : begin
        result = input_780;
      end
      10'b1100001101 : begin
        result = input_781;
      end
      10'b1100001110 : begin
        result = input_782;
      end
      10'b1100001111 : begin
        result = input_783;
      end
      10'b1100010000 : begin
        result = input_784;
      end
      10'b1100010001 : begin
        result = input_785;
      end
      10'b1100010010 : begin
        result = input_786;
      end
      10'b1100010011 : begin
        result = input_787;
      end
      10'b1100010100 : begin
        result = input_788;
      end
      10'b1100010101 : begin
        result = input_789;
      end
      10'b1100010110 : begin
        result = input_790;
      end
      10'b1100010111 : begin
        result = input_791;
      end
      10'b1100011000 : begin
        result = input_792;
      end
      10'b1100011001 : begin
        result = input_793;
      end
      10'b1100011010 : begin
        result = input_794;
      end
      10'b1100011011 : begin
        result = input_795;
      end
      10'b1100011100 : begin
        result = input_796;
      end
      10'b1100011101 : begin
        result = input_797;
      end
      10'b1100011110 : begin
        result = input_798;
      end
      10'b1100011111 : begin
        result = input_799;
      end
      10'b1100100000 : begin
        result = input_800;
      end
      10'b1100100001 : begin
        result = input_801;
      end
      10'b1100100010 : begin
        result = input_802;
      end
      10'b1100100011 : begin
        result = input_803;
      end
      10'b1100100100 : begin
        result = input_804;
      end
      10'b1100100101 : begin
        result = input_805;
      end
      10'b1100100110 : begin
        result = input_806;
      end
      10'b1100100111 : begin
        result = input_807;
      end
      10'b1100101000 : begin
        result = input_808;
      end
      10'b1100101001 : begin
        result = input_809;
      end
      10'b1100101010 : begin
        result = input_810;
      end
      10'b1100101011 : begin
        result = input_811;
      end
      10'b1100101100 : begin
        result = input_812;
      end
      10'b1100101101 : begin
        result = input_813;
      end
      10'b1100101110 : begin
        result = input_814;
      end
      10'b1100101111 : begin
        result = input_815;
      end
      10'b1100110000 : begin
        result = input_816;
      end
      10'b1100110001 : begin
        result = input_817;
      end
      10'b1100110010 : begin
        result = input_818;
      end
      10'b1100110011 : begin
        result = input_819;
      end
      10'b1100110100 : begin
        result = input_820;
      end
      10'b1100110101 : begin
        result = input_821;
      end
      10'b1100110110 : begin
        result = input_822;
      end
      10'b1100110111 : begin
        result = input_823;
      end
      10'b1100111000 : begin
        result = input_824;
      end
      10'b1100111001 : begin
        result = input_825;
      end
      10'b1100111010 : begin
        result = input_826;
      end
      10'b1100111011 : begin
        result = input_827;
      end
      10'b1100111100 : begin
        result = input_828;
      end
      10'b1100111101 : begin
        result = input_829;
      end
      10'b1100111110 : begin
        result = input_830;
      end
      10'b1100111111 : begin
        result = input_831;
      end
      10'b1101000000 : begin
        result = input_832;
      end
      10'b1101000001 : begin
        result = input_833;
      end
      10'b1101000010 : begin
        result = input_834;
      end
      10'b1101000011 : begin
        result = input_835;
      end
      10'b1101000100 : begin
        result = input_836;
      end
      10'b1101000101 : begin
        result = input_837;
      end
      10'b1101000110 : begin
        result = input_838;
      end
      10'b1101000111 : begin
        result = input_839;
      end
      10'b1101001000 : begin
        result = input_840;
      end
      10'b1101001001 : begin
        result = input_841;
      end
      10'b1101001010 : begin
        result = input_842;
      end
      10'b1101001011 : begin
        result = input_843;
      end
      10'b1101001100 : begin
        result = input_844;
      end
      10'b1101001101 : begin
        result = input_845;
      end
      10'b1101001110 : begin
        result = input_846;
      end
      10'b1101001111 : begin
        result = input_847;
      end
      10'b1101010000 : begin
        result = input_848;
      end
      10'b1101010001 : begin
        result = input_849;
      end
      10'b1101010010 : begin
        result = input_850;
      end
      10'b1101010011 : begin
        result = input_851;
      end
      10'b1101010100 : begin
        result = input_852;
      end
      10'b1101010101 : begin
        result = input_853;
      end
      10'b1101010110 : begin
        result = input_854;
      end
      10'b1101010111 : begin
        result = input_855;
      end
      10'b1101011000 : begin
        result = input_856;
      end
      10'b1101011001 : begin
        result = input_857;
      end
      10'b1101011010 : begin
        result = input_858;
      end
      10'b1101011011 : begin
        result = input_859;
      end
      10'b1101011100 : begin
        result = input_860;
      end
      10'b1101011101 : begin
        result = input_861;
      end
      10'b1101011110 : begin
        result = input_862;
      end
      10'b1101011111 : begin
        result = input_863;
      end
      10'b1101100000 : begin
        result = input_864;
      end
      10'b1101100001 : begin
        result = input_865;
      end
      10'b1101100010 : begin
        result = input_866;
      end
      10'b1101100011 : begin
        result = input_867;
      end
      10'b1101100100 : begin
        result = input_868;
      end
      10'b1101100101 : begin
        result = input_869;
      end
      10'b1101100110 : begin
        result = input_870;
      end
      10'b1101100111 : begin
        result = input_871;
      end
      10'b1101101000 : begin
        result = input_872;
      end
      10'b1101101001 : begin
        result = input_873;
      end
      10'b1101101010 : begin
        result = input_874;
      end
      10'b1101101011 : begin
        result = input_875;
      end
      10'b1101101100 : begin
        result = input_876;
      end
      10'b1101101101 : begin
        result = input_877;
      end
      10'b1101101110 : begin
        result = input_878;
      end
      10'b1101101111 : begin
        result = input_879;
      end
      10'b1101110000 : begin
        result = input_880;
      end
      10'b1101110001 : begin
        result = input_881;
      end
      10'b1101110010 : begin
        result = input_882;
      end
      10'b1101110011 : begin
        result = input_883;
      end
      10'b1101110100 : begin
        result = input_884;
      end
      10'b1101110101 : begin
        result = input_885;
      end
      10'b1101110110 : begin
        result = input_886;
      end
      10'b1101110111 : begin
        result = input_887;
      end
      10'b1101111000 : begin
        result = input_888;
      end
      10'b1101111001 : begin
        result = input_889;
      end
      10'b1101111010 : begin
        result = input_890;
      end
      10'b1101111011 : begin
        result = input_891;
      end
      10'b1101111100 : begin
        result = input_892;
      end
      10'b1101111101 : begin
        result = input_893;
      end
      10'b1101111110 : begin
        result = input_894;
      end
      10'b1101111111 : begin
        result = input_895;
      end
      10'b1110000000 : begin
        result = input_896;
      end
      10'b1110000001 : begin
        result = input_897;
      end
      10'b1110000010 : begin
        result = input_898;
      end
      10'b1110000011 : begin
        result = input_899;
      end
      10'b1110000100 : begin
        result = input_900;
      end
      10'b1110000101 : begin
        result = input_901;
      end
      10'b1110000110 : begin
        result = input_902;
      end
      10'b1110000111 : begin
        result = input_903;
      end
      10'b1110001000 : begin
        result = input_904;
      end
      10'b1110001001 : begin
        result = input_905;
      end
      10'b1110001010 : begin
        result = input_906;
      end
      10'b1110001011 : begin
        result = input_907;
      end
      10'b1110001100 : begin
        result = input_908;
      end
      10'b1110001101 : begin
        result = input_909;
      end
      10'b1110001110 : begin
        result = input_910;
      end
      10'b1110001111 : begin
        result = input_911;
      end
      10'b1110010000 : begin
        result = input_912;
      end
      10'b1110010001 : begin
        result = input_913;
      end
      10'b1110010010 : begin
        result = input_914;
      end
      10'b1110010011 : begin
        result = input_915;
      end
      10'b1110010100 : begin
        result = input_916;
      end
      10'b1110010101 : begin
        result = input_917;
      end
      10'b1110010110 : begin
        result = input_918;
      end
      10'b1110010111 : begin
        result = input_919;
      end
      10'b1110011000 : begin
        result = input_920;
      end
      10'b1110011001 : begin
        result = input_921;
      end
      10'b1110011010 : begin
        result = input_922;
      end
      10'b1110011011 : begin
        result = input_923;
      end
      10'b1110011100 : begin
        result = input_924;
      end
      10'b1110011101 : begin
        result = input_925;
      end
      10'b1110011110 : begin
        result = input_926;
      end
      10'b1110011111 : begin
        result = input_927;
      end
      10'b1110100000 : begin
        result = input_928;
      end
      10'b1110100001 : begin
        result = input_929;
      end
      10'b1110100010 : begin
        result = input_930;
      end
      10'b1110100011 : begin
        result = input_931;
      end
      10'b1110100100 : begin
        result = input_932;
      end
      10'b1110100101 : begin
        result = input_933;
      end
      10'b1110100110 : begin
        result = input_934;
      end
      10'b1110100111 : begin
        result = input_935;
      end
      10'b1110101000 : begin
        result = input_936;
      end
      10'b1110101001 : begin
        result = input_937;
      end
      10'b1110101010 : begin
        result = input_938;
      end
      10'b1110101011 : begin
        result = input_939;
      end
      10'b1110101100 : begin
        result = input_940;
      end
      10'b1110101101 : begin
        result = input_941;
      end
      10'b1110101110 : begin
        result = input_942;
      end
      10'b1110101111 : begin
        result = input_943;
      end
      10'b1110110000 : begin
        result = input_944;
      end
      10'b1110110001 : begin
        result = input_945;
      end
      10'b1110110010 : begin
        result = input_946;
      end
      10'b1110110011 : begin
        result = input_947;
      end
      10'b1110110100 : begin
        result = input_948;
      end
      10'b1110110101 : begin
        result = input_949;
      end
      10'b1110110110 : begin
        result = input_950;
      end
      10'b1110110111 : begin
        result = input_951;
      end
      10'b1110111000 : begin
        result = input_952;
      end
      10'b1110111001 : begin
        result = input_953;
      end
      10'b1110111010 : begin
        result = input_954;
      end
      10'b1110111011 : begin
        result = input_955;
      end
      10'b1110111100 : begin
        result = input_956;
      end
      10'b1110111101 : begin
        result = input_957;
      end
      10'b1110111110 : begin
        result = input_958;
      end
      10'b1110111111 : begin
        result = input_959;
      end
      10'b1111000000 : begin
        result = input_960;
      end
      10'b1111000001 : begin
        result = input_961;
      end
      10'b1111000010 : begin
        result = input_962;
      end
      10'b1111000011 : begin
        result = input_963;
      end
      10'b1111000100 : begin
        result = input_964;
      end
      10'b1111000101 : begin
        result = input_965;
      end
      10'b1111000110 : begin
        result = input_966;
      end
      10'b1111000111 : begin
        result = input_967;
      end
      10'b1111001000 : begin
        result = input_968;
      end
      10'b1111001001 : begin
        result = input_969;
      end
      10'b1111001010 : begin
        result = input_970;
      end
      10'b1111001011 : begin
        result = input_971;
      end
      10'b1111001100 : begin
        result = input_972;
      end
      10'b1111001101 : begin
        result = input_973;
      end
      10'b1111001110 : begin
        result = input_974;
      end
      10'b1111001111 : begin
        result = input_975;
      end
      10'b1111010000 : begin
        result = input_976;
      end
      10'b1111010001 : begin
        result = input_977;
      end
      10'b1111010010 : begin
        result = input_978;
      end
      10'b1111010011 : begin
        result = input_979;
      end
      10'b1111010100 : begin
        result = input_980;
      end
      10'b1111010101 : begin
        result = input_981;
      end
      10'b1111010110 : begin
        result = input_982;
      end
      10'b1111010111 : begin
        result = input_983;
      end
      10'b1111011000 : begin
        result = input_984;
      end
      10'b1111011001 : begin
        result = input_985;
      end
      10'b1111011010 : begin
        result = input_986;
      end
      10'b1111011011 : begin
        result = input_987;
      end
      10'b1111011100 : begin
        result = input_988;
      end
      10'b1111011101 : begin
        result = input_989;
      end
      10'b1111011110 : begin
        result = input_990;
      end
      10'b1111011111 : begin
        result = input_991;
      end
      10'b1111100000 : begin
        result = input_992;
      end
      10'b1111100001 : begin
        result = input_993;
      end
      10'b1111100010 : begin
        result = input_994;
      end
      10'b1111100011 : begin
        result = input_995;
      end
      10'b1111100100 : begin
        result = input_996;
      end
      10'b1111100101 : begin
        result = input_997;
      end
      10'b1111100110 : begin
        result = input_998;
      end
      10'b1111100111 : begin
        result = input_999;
      end
      10'b1111101000 : begin
        result = input_1000;
      end
      10'b1111101001 : begin
        result = input_1001;
      end
      10'b1111101010 : begin
        result = input_1002;
      end
      10'b1111101011 : begin
        result = input_1003;
      end
      10'b1111101100 : begin
        result = input_1004;
      end
      10'b1111101101 : begin
        result = input_1005;
      end
      10'b1111101110 : begin
        result = input_1006;
      end
      10'b1111101111 : begin
        result = input_1007;
      end
      10'b1111110000 : begin
        result = input_1008;
      end
      10'b1111110001 : begin
        result = input_1009;
      end
      10'b1111110010 : begin
        result = input_1010;
      end
      10'b1111110011 : begin
        result = input_1011;
      end
      10'b1111110100 : begin
        result = input_1012;
      end
      10'b1111110101 : begin
        result = input_1013;
      end
      10'b1111110110 : begin
        result = input_1014;
      end
      10'b1111110111 : begin
        result = input_1015;
      end
      10'b1111111000 : begin
        result = input_1016;
      end
      10'b1111111001 : begin
        result = input_1017;
      end
      10'b1111111010 : begin
        result = input_1018;
      end
      10'b1111111011 : begin
        result = input_1019;
      end
      10'b1111111100 : begin
        result = input_1020;
      end
      10'b1111111101 : begin
        result = input_1021;
      end
      10'b1111111110 : begin
        result = input_1022;
      end
      default : begin
        result = input_1023;
      end
    endcase
    MUX_v_57_1024_2 = result;
  end
  endfunction


  function automatic [61:0] signext_62_57;
    input [56:0] vector;
  begin
    signext_62_57= {{5{vector[56]}}, vector};
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i10_1o62_e041a31844d9eff753e17f0437c907cdbd_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Mon May 27 10:57:40 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i10_1o62_e041a31844d9eff753e17f0437c907cdbd
// ------------------------------------------------------------------


module ROM_1i10_1o62_e041a31844d9eff753e17f0437c907cdbd (
  I_1, O_1
);
  input [9:0] I_1;
  output [61:0] O_1;


  wire[56:0] r_ac_ieee_float_base_slc_gm_im_tab_d_rom_1_BUTTERFLY_if_r_ac_ieee_float_base_mux_nl;

  // Interconnect Declarations for Component Instantiations 
  assign r_ac_ieee_float_base_slc_gm_im_tab_d_rom_1_BUTTERFLY_if_r_ac_ieee_float_base_mux_nl
      = MUX_v_57_1024_2(57'b000000000000000000000000000000000000000000000000000000000,
      57'b111110000000000000000000000000000000000000000000000000000, 57'b111100110101000001001111001100110011111110011101111001101,
      57'b111100110101000001001111001100110011111110011101111001101, 57'b111011000011111011110001010100110101011101010100101100011,
      57'b111101101100100000110101111001111001100101000110101000110, 57'b111101101100100000110101111001111001100101000110101000110,
      57'b111011000011111011110001010100110101011101010100101100011, 57'b111001000111110001011100000111100011010011010011000001011,
      57'b111101111011000101001011111001111111101110101110010110000, 57'b111101010100110110110011000101001000011101010000110100011,
      57'b111100001110001110011101100111001101011100110100011001000, 57'b111100001110001110011101100111001101011100110100011001000,
      57'b111101010100110110110011000101001000011101010000110100011, 57'b111101111011000101001011111001111111101110101110010110000,
      57'b111001000111110001011100000111100011010011010011000001011, 57'b110111001000101111010011010111100001010011011010000101100,
      57'b111101111110110001000110110100011110100010010010100100110, 57'b111101000101111001000000001101011000101010001011101000001,
      57'b111100100010011001111001100100101000010010001110111010110, 57'b111011110001010110101110100111000000001101111011000111011,
      57'b111101100001110001011001011110001100000001011110110110001, 57'b111101110100111110100000101010110110001100010110111011010,
      57'b111010010100101000000011000101110110101011001111100000110, 57'b111010010100101000000011000101110110101011001111100000110,
      57'b111101110100111110100000101010110110001100010110111011010, 57'b111101100001110001011001011110001100000001011110110110001,
      57'b111011110001010110101110100111000000001101111011000111011, 57'b111100100010011001111001100100101000010010001110111010110,
      57'b111101000101111001000000001101011000101010001011101000001, 57'b111101111110110001000110110100011110100010010010100100110,
      57'b110111001000101111010011010111100001010011011010000101100, 57'b110101001000111110110010111110001000011011101100000010100,
      57'b111101111111101100010000111100011011110010110110101111110, 57'b111100111101101011101111100100010011010101010111110101111,
      57'b111100101011111010110100100110100100011001110110010100000, 57'b111011011010111010001000000001001111000010101110011000000,
      57'b111101100111011010111101011110100001111001100011101110011, 57'b111101110001000010010000100000100111101101000011011100101,
      57'b111010101100011111001101001110101101010110001111111011101, 57'b111001111000110011111100101111011001000010101111100011011,
      57'b111101111000010100111111011111011100100100011000011010111, 57'b111101011011100101000001101000101000110010110111000111110,
      57'b111100000011100111000011110011001001000101111111111101110, 57'b111100011000011111111011111111100111000010111000000110101,
      57'b111101001101100111110000001000111111100111000011101000001, 57'b111101111101001110101010101111111000010001010010100010111,
      57'b111000010110010000001000001101110100011100110000100111010, 57'b111000010110010000001000001101110100011100110000100111010,
      57'b111101111101001110101010101111111000010001010010100010111, 57'b111101001101100111110000001000111111100111000011101000001,
      57'b111100011000011111111011111111100111000010111000000110101, 57'b111100000011100111000011110011001001000101111111111101110,
      57'b111101011011100101000001101000101000110010110111000111110, 57'b111101111000010100111111011111011100100100011000011010111,
      57'b111001111000110011111100101111011001000010101111100011011, 57'b111010101100011111001101001110101101010110001111111011101,
      57'b111101110001000010010000100000100111101101000011011100101, 57'b111101100111011010111101011110100001111001100011101110011,
      57'b111011011010111010001000000001001111000010101110011000000, 57'b111100101011111010110100100110100100011001110110010100000,
      57'b111100111101101011101111100100010011010101010111110101111, 57'b111101111111101100010000111100011011110010110110101111110,
      57'b110101001000111110110010111110001000011011101100000010100, 57'b110011001001000010101010111110111101000110110011001111110,
      57'b111101111111111011000100001100000100001001100110100001101, 57'b111100111001011010000100000110111111011111111111110010110,
      57'b111100110000100001011011101010101000111010010110011011111, 57'b111011001111011110111100101000011101010001110110110001010,
      57'b111101101010000010011010011010001010011011100100100111010, 57'b111101101110110110001001110110110110011001100001000111100,
      57'b111010111000010001000010100110000111110100100010110011111, 57'b111001100000010111000001001101010011111100100111101100011,
      57'b111101111001110001111001110101100011001001110010110001001, 57'b111101011000010010000101001011000000101010000001000000000,
      57'b111100001000111101011001101010100000110110100101100100011, 57'b111100010011011010000010101001100110111010001001011011111,
      57'b111101010001010011010011110100000010001100010011110000010, 57'b111101111100001110110010011111010011100010100101110101001,
      57'b111000101111000100001010001000100100010110011111111000110, 57'b110111111010101100100111001010110101010010111001100001110,
      57'b111101111110000100110010001110000111000011001111111010011, 57'b111101001001110100010001001001001100100100110001111111011,
      57'b111100011101011111111101000101001001000000101000010111001, 57'b111011111100010111010010011011011111110001001101010111010,
      57'b111101011110101111100000010101100011011111001010100101010, 57'b111101110110101110100000011100111011010000100100101100011,
      57'b111010001000100011101001001100010101100011111011001110111, 57'b111010100000100110101110010010100000101110110011000000001,
      57'b111101110011000101000100011101100010010001110000100010010, 57'b111101100100101010100101100100001001101000001000111110101,
      57'b111011100110001100110111010011001001100011100010001011110, 57'b111100100111001101100101010111011111000111110010111101001,
      57'b111101000001110110000111000001011111111111001011101101110, 57'b111101111111010011100110110101101000000011000100000111010,
      57'b110110010110101010010000010010010110011100001100111110110, 57'b110110010110101010010000010010010110011100001100111110110,
      57'b111101111111010011100110110101101000000011000100000111010, 57'b111101000001110110000111000001011111111111001011101101110,
      57'b111100100111001101100101010111011111000111110010111101001, 57'b111011100110001100110111010011001001100011100010001011110,
      57'b111101100100101010100101100100001001101000001000111110101, 57'b111101110011000101000100011101100010010001110000100010010,
      57'b111010100000100110101110010010100000101110110011000000001, 57'b111010001000100011101001001100010101100011111011001110111,
      57'b111101110110101110100000011100111011010000100100101100011, 57'b111101011110101111100000010101100011011111001010100101010,
      57'b111011111100010111010010011011011111110001001101010111010, 57'b111100011101011111111101000101001001000000101000010111001,
      57'b111101001001110100010001001001001100100100110001111111011, 57'b111101111110000100110010001110000111000011001111111010011,
      57'b110111111010101100100111001010110101010010111001100001110, 57'b111000101111000100001010001000100100010110011111111000110,
      57'b111101111100001110110010011111010011100010100101110101001, 57'b111101010001010011010011110100000010001100010011110000010,
      57'b111100010011011010000010101001100110111010001001011011111, 57'b111100001000111101011001101010100000110110100101100100011,
      57'b111101011000010010000101001011000000101010000001000000000, 57'b111101111001110001111001110101100011001001110010110001001,
      57'b111001100000010111000001001101010011111100100111101100011, 57'b111010111000010001000010100110000111110100100010110011111,
      57'b111101101110110110001001110110110110011001100001000111100, 57'b111101101010000010011010011010001010011011100100100111010,
      57'b111011001111011110111100101000011101010001110110110001010, 57'b111100110000100001011011101010101000111010010110011011111,
      57'b111100111001011010000100000110111111011111111111110010110, 57'b111101111111111011000100001100000100001001100110100001101,
      57'b110011001001000010101010111110111101000110110011001111110, 57'b110001001001000011101000111111100110111101100011110000100,
      57'b111101111111111110110001000010110100110111001001011011011, 57'b111100110111001110100010001010100111010101010100010101111,
      57'b111100110010110010001100100100101111100000111100000111101, 57'b111011001001101110010101001100011101111001001001111010111,
      57'b111101101011010010110000101110011110010011110011010001011, 57'b111101101101101100101001001100010001110001010000010011011,
      57'b111010111110000111010100100110001000111011100110011100111, 57'b111001010100000101010000000100101101100000000010001010001,
      57'b111101111010011100110000000111011000010110010111100101101, 57'b111101010110100101011110010011110001000011101010100010001,
      57'b111100001011100110100110101100011110111101101101101001001, 57'b111100010000110100111100110011001001100111110101101011001,
      57'b111101010011000110000100100011011000000101111101011100010, 57'b111101111011101011001100110100011101000010010000001110111,
      57'b111000111011011011101100111011110010100001011111100110001, 57'b110111100001101111000010111000111100111101100001011010101,
      57'b111101111110011100001010111111101011011011010011001111011, 57'b111101000111110111100110010100011111011111001010000001101,
      57'b111100011111111101101100101010011010001010101011011010100, 57'b111011110110111000001100101010010111011110111100011010110,
      57'b111101100000010001100010000100110011100100101010101001001, 57'b111101110101110111101100011001000110111110000101101110100,
      57'b111010001110100110100010000111111010011001101101100111110, 57'b111010011010101000001000011000010111000011000000101010010,
      57'b111101110100000010111101110101011010011001101000100001101, 57'b111101100011001111000101100110100100010000111001110011011,
      57'b111011101011110010111011101011011100001101110001110001001, 57'b111100100100110100100010010011011100110110000100100111001,
      57'b111101000011111000100000000001111101110100010111010111111, 57'b111101111111000011100101011111100101111010101101100001001,
      57'b110110101111101101101000000001010100110101010010000011001, 57'b110101111011001010110111001111001111110000010000011100000,
      57'b111101111111100001001010101100101100011100111000110101101, 57'b111100111111110001110110011100011010101110001011101110001,
      57'b111100101001100101000001010010010101000110101010110010110, 57'b111011100000100100100100111011000000000010001111011100111,
      57'b111101100110000011111000011110011111111001111110001011100, 57'b111101110010000100110101001001011001010111100000101111110,
      57'b111010100110100011110001001000010011110001110011101101010, 57'b111010000010011111011100000001110001101111111110110101110,
      57'b111101110111100010111100010100011111001000111001111000010, 57'b111101011101001011010101001100111001101011001000011010010,
      57'b111100000000111001111110010000111010011000011111010110111, 57'b111100011011000000101100010110001000001100101100111110011,
      57'b111101001011101110111111011110100110001111101011101000010, 57'b111101111101101010111100101110001100101011101011101000001,
      57'b111000001001110011111000011001110110110101111010101110111, 57'b111000100010101010111011010110001001010010011111001011010,
      57'b111101111100101111111100100100100110010010000100110011011, 57'b111101001111011110100001111101111001010011010111110010100,
      57'b111100010101111101101101100100101111110101111001111101010, 57'b111100000110010010111000001001101010111011000100110001111,
      57'b111101011001111100100110100111110111101010101011100010010, 57'b111101111001000100101001011110111011101100011101011011010,
      57'b111001101100100110100111111100101010001010100001100010001, 57'b111010110010011000111110111011101001111110010011111000110,
      57'b111101101111111101010111001100010001011011011111000101011, 57'b111101101000101111110011101110100001111100011010111011100,
      57'b111011010101001101100100000101011011011010011111111001010, 57'b111100101110001110111101110111110011001010000000110001100,
      57'b111100111011100011110011101011111000000110111001001100001, 57'b111101111111110100111001011101111111111101111011101011101,
      57'b110100010110110000110010101110101100101000101010111001101, 57'b110100010110110000110010101110101100101000101010111001101,
      57'b111101111111110100111001011101111111111101111011101011101, 57'b111100111011100011110011101011111000000110111001001100001,
      57'b111100101110001110111101110111110011001010000000110001100, 57'b111011010101001101100100000101011011011010011111111001010,
      57'b111101101000101111110011101110100001111100011010111011100, 57'b111101101111111101010111001100010001011011011111000101011,
      57'b111010110010011000111110111011101001111110010011111000110, 57'b111001101100100110100111111100101010001010100001100010001,
      57'b111101111001000100101001011110111011101100011101011011010, 57'b111101011001111100100110100111110111101010101011100010010,
      57'b111100000110010010111000001001101010111011000100110001111, 57'b111100010101111101101101100100101111110101111001111101010,
      57'b111101001111011110100001111101111001010011010111110010100, 57'b111101111100101111111100100100100110010010000100110011011,
      57'b111000100010101010111011010110001001010010011111001011010, 57'b111000001001110011111000011001110110110101111010101110111,
      57'b111101111101101010111100101110001100101011101011101000001, 57'b111101001011101110111111011110100110001111101011101000010,
      57'b111100011011000000101100010110001000001100101100111110011, 57'b111100000000111001111110010000111010011000011111010110111,
      57'b111101011101001011010101001100111001101011001000011010010, 57'b111101110111100010111100010100011111001000111001111000010,
      57'b111010000010011111011100000001110001101111111110110101110, 57'b111010100110100011110001001000010011110001110011101101010,
      57'b111101110010000100110101001001011001010111100000101111110, 57'b111101100110000011111000011110011111111001111110001011100,
      57'b111011100000100100100100111011000000000010001111011100111, 57'b111100101001100101000001010010010101000110101010110010110,
      57'b111100111111110001110110011100011010101110001011101110001, 57'b111101111111100001001010101100101100011100111000110101101,
      57'b110101111011001010110111001111001111110000010000011100000, 57'b110110101111101101101000000001010100110101010010000011001,
      57'b111101111111000011100101011111100101111010101101100001001, 57'b111101000011111000100000000001111101110100010111010111111,
      57'b111100100100110100100010010011011100110110000100100111001, 57'b111011101011110010111011101011011100001101110001110001001,
      57'b111101100011001111000101100110100100010000111001110011011, 57'b111101110100000010111101110101011010011001101000100001101,
      57'b111010011010101000001000011000010111000011000000101010010, 57'b111010001110100110100010000111111010011001101101100111110,
      57'b111101110101110111101100011001000110111110000101101110100, 57'b111101100000010001100010000100110011100100101010101001001,
      57'b111011110110111000001100101010010111011110111100011010110, 57'b111100011111111101101100101010011010001010101011011010100,
      57'b111101000111110111100110010100011111011111001010000001101, 57'b111101111110011100001010111111101011011011010011001111011,
      57'b110111100001101111000010111000111100111101100001011010101, 57'b111000111011011011101100111011110010100001011111100110001,
      57'b111101111011101011001100110100011101000010010000001110111, 57'b111101010011000110000100100011011000000101111101011100010,
      57'b111100010000110100111100110011001001100111110101101011001, 57'b111100001011100110100110101100011110111101101101101001001,
      57'b111101010110100101011110010011110001000011101010100010001, 57'b111101111010011100110000000111011000010110010111100101101,
      57'b111001010100000101010000000100101101100000000010001010001, 57'b111010111110000111010100100110001000111011100110011100111,
      57'b111101101101101100101001001100010001110001010000010011011, 57'b111101101011010010110000101110011110010011110011010001011,
      57'b111011001001101110010101001100011101111001001001111010111, 57'b111100110010110010001100100100101111100000111100000111101,
      57'b111100110111001110100010001010100111010101010100010101111, 57'b111101111111111110110001000010110100110111001001011011011,
      57'b110001001001000011101000111111100110111101100011110000100, 57'b101111001001000011111000011111110011001110000000001110001,
      57'b111101111111111111101100010000101100011101000101010010010, 57'b111100110110001000000110101110011110000011000001001110101,
      57'b111100110011111001111011110000100100100011010111100010000, 57'b111011000110110101010010100101110110010001010010010110000,
      57'b111101101011111010000101100000010101110001110110011111001, 57'b111101101101000111000001110101001011001101000100110001000,
      57'b111011000001000001110001110110000010011101010101011000100, 57'b111001001101111011100101111110010110111000100001101100110,
      57'b111101111010110001010001010110001011110001001111010000100, 57'b111101010101101110011001001011001000101101100000011010100,
      57'b111100001100111010101101000001001111100101011100110111000, 57'b111100001111100001111000010001011101111001000011000011011,
      57'b111101010011111110101100001010010100111111110011010011101, 57'b111101111011011000011111101111101111101011011101110110111,
      57'b111001000001100110110011011101000100111000110010011000110, 57'b110111010101001111011011100100100010010010101110000000011,
      57'b111101111110100110111100100010100001000100000101110000100, 57'b111101000110111000100010100110011000101101001100011001100,
      57'b111100100001001011111111100010111100011100110101110110001, 57'b111011110100000111110000011101010111110000101000100010100,
      57'b111101100001000001101111000111111101010010111000110110000, 57'b111101110101011011011001011101000111001111010100010001110,
      57'b111010010001100111011101110101011110000111011101101110001, 57'b111010010111101000010001011011010111011000000001110000111,
      57'b111101110100100001000010000110110000111011111011111110010, 57'b111101100010100000100001000000001001010110110100100000111,
      57'b111011101110100101000111100010100100000011100110001011000, 57'b111100100011100111011010100011011100110000111001101000111,
      57'b111101000100111000111111010011010010011011101010010101010, 57'b111101111110111010101001110011111111100011111010001010110,
      57'b110110111100001110101100001101010010111010101101100100001, 57'b110101100010000101000110100010010110000001101011111100011,
      57'b111101111111100111000001100001111100011010101011101011100, 57'b111100111110101111000001101101100110000110011110110110010,
      57'b111100101010110000001000000111000100101110101000100110111, 57'b111011011101101111100111100100011000001001011110100000001,
      57'b111101100110101111101100110001001100010110011001011110110, 57'b111101110001100011110101011101000011100001100111000100101,
      57'b111010101001100001101100010000000101011110011110000100100, 57'b111001111110111001101110000011010110111111110110111111001,
      57'b111101110111111100010001000001100000010111001010111101100, 57'b111101011100011000011100011010010011101010000010011101001,
      57'b111100000010010000101011000100110101011100010001000011010, 57'b111100011001110000100000000001101000011001000111001010111,
      57'b111101001100101011100111100101110110110000000110100100010, 57'b111101111101011101000111010001110010001101100111110111011,
      57'b111000010000000010001011011010100111011000111101111001111, 57'b111000011100011101101101110110000110011011000110100010100,
      57'b111101111100111111100111001010101101011011011001011001000, 57'b111101001110100011011000111110101111010101000000011010101,
      57'b111100010111001111000000011100011111010001110101000010111, 57'b111100000100111101001000001110100000101111100010111100001,
      57'b111101011010110001000100111111110100100100001010000000101, 57'b111101111000101101000111101010011111101110010000001011101,
      57'b111001110010101101100101000011110000100000001101000011011, 57'b111010101111011100010011100110111100111101010011010010011,
      57'b111101110000100000000110011001010001010011000000010101100, 57'b111101101000000101101010011111110101100101011110110010010,
      57'b111011011000000100000110101101100011111110100000000001001, 57'b111100101101000101000110100101010010111010111001001010000,
      57'b111100111100101000000000001010111010011110101010111100101, 57'b111101111111110000111000111011010110110111000000111011111,
      57'b110100101111111000000000011010010100100001100110101000011, 57'b110011111011010010011011100110001110100011100111100000001,
      57'b111101111111111000010010100011101111100011101001111111000, 57'b111100111010011111001010010001101101010001101001010001101,
      57'b111100101111011000011010010010101100000110111000001110100, 57'b111011010010010110100000100100111110111101010000111100101,
      57'b111101101001011001011001000100000111000001110111110011111, 57'b111101101111011010000010111110111110111100100011111011010,
      57'b111010110101010101001110101111101110001110111111000010111, 57'b111001100110011111000110010110011000100101011001010000110,
      57'b111101111001011011100100111001001000010001001101010011101, 57'b111101011001000111100110101000111000000000001001110110100,
      57'b111100000111101000010011010111011001010101000111001111110, 57'b111100010100101100000011100100111011000101001110010101000,
      57'b111101010000011001001010111101010101110101111100100110111, 57'b111101111100011111101010111111111101011100100000111011011,
      57'b111000101000110111101111110000101100101111100010111110010, 57'b111000000011100101010000001000111101110101000001100011101,
      57'b111101111101111000001011000010111111001000100000110000110, 57'b111101001010110001110111111100100100011100110110111010111,
      57'b111100011100010000100000110000101110111111110101100100010, 57'b111011111111000101111011001001011111001110001001000010000,
      57'b111101011101111101101011111000100100100111000000011101010, 57'b111101110111001001000001011100010010110101001110110111100,
      57'b111010000101100001101100111001111110110111101101110010000, 57'b111010100011100101011100010100101010101110001000001010100,
      57'b111101110010100101001111100000100011100101001111111111100, 57'b111101100101010111100000101101001101000001011100100000000,
      57'b111011100011011000111111101001001100101110000000000001011, 57'b111100101000011001100000010011111010110011010000010011011,
      57'b111101000000110100001101100110011101101010111101011001100, 57'b111101111111011010101100011101100101101100111001111000100,
      57'b110110001010001000000000100110100110101110000100110110011, 57'b110110100011001100001000101111001001001110010000010010110,
      57'b111101111111001011111001110101111001011100011100101000000, 57'b111101000010110111100010100011010111010010101100011001100,
      57'b111100100110000001010000101000101111011000000000000000100, 57'b111011101001000000001011011101000111010011101101101011011,
      57'b111101100011111101000111001010010001000110011110011110011, 57'b111101110011100100010011111011011011010101001011101000100,
      57'b111010011101100111100111011111010000001000001010010110111, 57'b111010001011100101010000011010111011101100101000101110111,
      57'b111101110110010011011001011010011110000111011111110000100, 57'b111101011111100000110010011100001010100110111011111011101,
      57'b111011111001101000000010110010110001111111101000001100111, 57'b111100011110101111000001000111000110001011000001101000100,
      57'b111101001000110110001011001101111110101001001110110100010, 57'b111101111110010000110010001101100111111101011011100100001,
      57'b110111101110001110000111011001011101011101001111111001001, 57'b111000110101010000001001100000100111101100100101010110010,
      57'b111101111011111101010011000101001111001100011110101101110, 57'b111101010010001100111100011001000000100011001101011001000,
      57'b111100010010000111101010111111011100110001010110000011111, 57'b111100001010010010001010110101111001100110110110011101011,
      57'b111101010111011100000010010110100001111000001010001110100, 57'b111101111010000111101000010000101111111111001001011011101,
      57'b111001011010001110011001011101111001111010110011100100010, 57'b111010111011001100011010000001111001001000001100011110110,
      57'b111101101110010001101011111001011010000010000001001100000, 57'b111101101010101010110111101010010111010010011111010110001,
      57'b111011001100100110111000101100001010000011011110111111111, 57'b111100110001101010000001110100011000111000001101111101001,
      57'b111100111000010100100001010110011000101110110110101111010, 57'b111101111111111101001110010110100010010110101000110100001,
      57'b110010010110110010011011010111011111000110000111011111101, 57'b110010010110110010011011010111011111000110000111011111101,
      57'b111101111111111101001110010110100010010110101000110100001, 57'b111100111000010100100001010110011000101110110110101111010,
      57'b111100110001101010000001110100011000111000001101111101001, 57'b111011001100100110111000101100001010000011011110111111111,
      57'b111101101010101010110111101010010111010010011111010110001, 57'b111101101110010001101011111001011010000010000001001100000,
      57'b111010111011001100011010000001111001001000001100011110110, 57'b111001011010001110011001011101111001111010110011100100010,
      57'b111101111010000111101000010000101111111111001001011011101, 57'b111101010111011100000010010110100001111000001010001110100,
      57'b111100001010010010001010110101111001100110110110011101011, 57'b111100010010000111101010111111011100110001010110000011111,
      57'b111101010010001100111100011001000000100011001101011001000, 57'b111101111011111101010011000101001111001100011110101101110,
      57'b111000110101010000001001100000100111101100100101010110010, 57'b110111101110001110000111011001011101011101001111111001001,
      57'b111101111110010000110010001101100111111101011011100100001, 57'b111101001000110110001011001101111110101001001110110100010,
      57'b111100011110101111000001000111000110001011000001101000100, 57'b111011111001101000000010110010110001111111101000001100111,
      57'b111101011111100000110010011100001010100110111011111011101, 57'b111101110110010011011001011010011110000111011111110000100,
      57'b111010001011100101010000011010111011101100101000101110111, 57'b111010011101100111100111011111010000001000001010010110111,
      57'b111101110011100100010011111011011011010101001011101000100, 57'b111101100011111101000111001010010001000110011110011110011,
      57'b111011101001000000001011011101000111010011101101101011011, 57'b111100100110000001010000101000101111011000000000000000100,
      57'b111101000010110111100010100011010111010010101100011001100, 57'b111101111111001011111001110101111001011100011100101000000,
      57'b110110100011001100001000101111001001001110010000010010110, 57'b110110001010001000000000100110100110101110000100110110011,
      57'b111101111111011010101100011101100101101100111001111000100, 57'b111101000000110100001101100110011101101010111101011001100,
      57'b111100101000011001100000010011111010110011010000010011011, 57'b111011100011011000111111101001001100101110000000000001011,
      57'b111101100101010111100000101101001101000001011100100000000, 57'b111101110010100101001111100000100011100101001111111111100,
      57'b111010100011100101011100010100101010101110001000001010100, 57'b111010000101100001101100111001111110110111101101110010000,
      57'b111101110111001001000001011100010010110101001110110111100, 57'b111101011101111101101011111000100100100111000000011101010,
      57'b111011111111000101111011001001011111001110001001000010000, 57'b111100011100010000100000110000101110111111110101100100010,
      57'b111101001010110001110111111100100100011100110110111010111, 57'b111101111101111000001011000010111111001000100000110000110,
      57'b111000000011100101010000001000111101110101000001100011101, 57'b111000101000110111101111110000101100101111100010111110010,
      57'b111101111100011111101010111111111101011100100000111011011, 57'b111101010000011001001010111101010101110101111100100110111,
      57'b111100010100101100000011100100111011000101001110010101000, 57'b111100000111101000010011010111011001010101000111001111110,
      57'b111101011001000111100110101000111000000000001001110110100, 57'b111101111001011011100100111001001000010001001101010011101,
      57'b111001100110011111000110010110011000100101011001010000110, 57'b111010110101010101001110101111101110001110111111000010111,
      57'b111101101111011010000010111110111110111100100011111011010, 57'b111101101001011001011001000100000111000001110111110011111,
      57'b111011010010010110100000100100111110111101010000111100101, 57'b111100101111011000011010010010101100000110111000001110100,
      57'b111100111010011111001010010001101101010001101001010001101, 57'b111101111111111000010010100011101111100011101001111111000,
      57'b110011111011010010011011100110001110100011100111100000001, 57'b110100101111111000000000011010010100100001100110101000011,
      57'b111101111111110000111000111011010110110111000000111011111, 57'b111100111100101000000000001010111010011110101010111100101,
      57'b111100101101000101000110100101010010111010111001001010000, 57'b111011011000000100000110101101100011111110100000000001001,
      57'b111101101000000101101010011111110101100101011110110010010, 57'b111101110000100000000110011001010001010011000000010101100,
      57'b111010101111011100010011100110111100111101010011010010011, 57'b111001110010101101100101000011110000100000001101000011011,
      57'b111101111000101101000111101010011111101110010000001011101, 57'b111101011010110001000100111111110100100100001010000000101,
      57'b111100000100111101001000001110100000101111100010111100001, 57'b111100010111001111000000011100011111010001110101000010111,
      57'b111101001110100011011000111110101111010101000000011010101, 57'b111101111100111111100111001010101101011011011001011001000,
      57'b111000011100011101101101110110000110011011000110100010100, 57'b111000010000000010001011011010100111011000111101111001111,
      57'b111101111101011101000111010001110010001101100111110111011, 57'b111101001100101011100111100101110110110000000110100100010,
      57'b111100011001110000100000000001101000011001000111001010111, 57'b111100000010010000101011000100110101011100010001000011010,
      57'b111101011100011000011100011010010011101010000010011101001, 57'b111101110111111100010001000001100000010111001010111101100,
      57'b111001111110111001101110000011010110111111110110111111001, 57'b111010101001100001101100010000000101011110011110000100100,
      57'b111101110001100011110101011101000011100001100111000100101, 57'b111101100110101111101100110001001100010110011001011110110,
      57'b111011011101101111100111100100011000001001011110100000001, 57'b111100101010110000001000000111000100101110101000100110111,
      57'b111100111110101111000001101101100110000110011110110110010, 57'b111101111111100111000001100001111100011010101011101011100,
      57'b110101100010000101000110100010010110000001101011111100011, 57'b110110111100001110101100001101010010111010101101100100001,
      57'b111101111110111010101001110011111111100011111010001010110, 57'b111101000100111000111111010011010010011011101010010101010,
      57'b111100100011100111011010100011011100110000111001101000111, 57'b111011101110100101000111100010100100000011100110001011000,
      57'b111101100010100000100001000000001001010110110100100000111, 57'b111101110100100001000010000110110000111011111011111110010,
      57'b111010010111101000010001011011010111011000000001110000111, 57'b111010010001100111011101110101011110000111011101101110001,
      57'b111101110101011011011001011101000111001111010100010001110, 57'b111101100001000001101111000111111101010010111000110110000,
      57'b111011110100000111110000011101010111110000101000100010100, 57'b111100100001001011111111100010111100011100110101110110001,
      57'b111101000110111000100010100110011000101101001100011001100, 57'b111101111110100110111100100010100001000100000101110000100,
      57'b110111010101001111011011100100100010010010101110000000011, 57'b111001000001100110110011011101000100111000110010011000110,
      57'b111101111011011000011111101111101111101011011101110110111, 57'b111101010011111110101100001010010100111111110011010011101,
      57'b111100001111100001111000010001011101111001000011000011011, 57'b111100001100111010101101000001001111100101011100110111000,
      57'b111101010101101110011001001011001000101101100000011010100, 57'b111101111010110001010001010110001011110001001111010000100,
      57'b111001001101111011100101111110010110111000100001101100110, 57'b111011000001000001110001110110000010011101010101011000100,
      57'b111101101101000111000001110101001011001101000100110001000, 57'b111101101011111010000101100000010101110001110110011111001,
      57'b111011000110110101010010100101110110010001010010010110000, 57'b111100110011111001111011110000100100100011010111100010000,
      57'b111100110110001000000110101110011110000011000001001110101, 57'b111101111111111111101100010000101100011101000101010010010,
      57'b101111001001000011111000011111110011001110000000001110001, 57'b101101001001000011111100010111110110011001010010010111010,
      57'b111101111111111111111011000100001011000100001110100000010, 57'b111100110101100100101110011101101001011111110001010011100,
      57'b111100110100011101101000111101010101000011001110001110001, 57'b111011000101011000100101110000110110101011110110101000100,
      57'b111101101100001101100010010000100010001011010010001001111, 57'b111101101100110100000000011011101100010110011110101000110,
      57'b111011000010011110110101010101010111100111001000000111111, 57'b111001001010110110100100111101001101101100010101011111010,
      57'b111101111010111011010011011101101010000110110100001011101, 57'b111101010101010010101010001111010001011001011100110001110,
      57'b111100001101100100101000000010111000100110111001110111111, 57'b111100001110111000001101101100100110111000100100001110010,
      57'b111101010100011010110011101101110010101000101101011010010, 57'b111101111011001110111010101010110100010000011110011101110,
      57'b111001000100101100001011100100111110001000001100000000100, 57'b110111001110111111011011011101011001001001010100001011100,
      57'b111101111110101100000110100101101101001110101110010011110, 57'b111101000110011000110101001110101000110000100011001010101,
      57'b111100100001110010111111101011011001010100100001110000000, 57'b111011110010101111010100001101101001111001101100000100101,
      57'b111101100001011001101000101001001001100011110001111110001, 57'b111101110101001101000001110010011111001100101100000000000,
      57'b111010010011000111110011010011001010101010101010010111010, 57'b111010010110001000001101001001110100101010100010100100000,
      57'b111101110100101111110110000110110000000010110101100110000, 57'b111101100010001001000001100110001010000011100000000000100,
      57'b111011101111111101111111101100110101010010100000111011110, 57'b111100100011000000101101001101001001010110011001010100010,
      57'b111101000101011001000011100011110110111100001110110001000, 57'b111101111110110101111101001110101000101000101001110001100,
      57'b110111000010011111000011100010010110000010011000010100001, 57'b110101010101100010000000110111101010111111000001100010111,
      57'b111101111111101001101110001010100101100011011111011010011, 57'b111100111110001101011100010011100111000101101001100110011,
      57'b111100101011010101100001101010001100101110110010010011111, 57'b111011011100010100111100000010100111111010101011010010011,
      57'b111101100111000101011001100100111100110011010000001100000, 57'b111101110001010011000111101000100001110010001100101111010,
      57'b111010101011000000100000000010010111101000110011110110100, 57'b111001111011110110111010010000000101111010011100000000010,
      57'b111101111000001000101101000010100110011110111001110001100, 57'b111101011011111110110011010000110111001111001001011101001,
      57'b111100000010111011111001111101100001100011011100010110111, 57'b111100011001001000010000111101100010010011010011000011111,
      57'b111101001101001001101111110100100001010110000011010110010, 57'b111101111101010101111101111001011000011001111110111011100,
      57'b111000010011001001001100101001101111111010011010000001001, 57'b111000011001010110111101111111001010001010001011010100111,
      57'b111101111101000111001101110101100011110100001011110010001, 57'b111101001110000101101000100010000111100000111010111000010,
      57'b111100010111110111100001001001011010001000001000000010101, 57'b111100000100010010001000100100000001100101011000010001100,
      57'b111101011011001011000111100010100111111011011110001000111, 57'b111101111000100001001000010111100100010011000111101011111,
      57'b111001110101110000110101101000110001011011110001101001000, 57'b111010101101111101110011110001011100111011011001110110110,
      57'b111101110000110001010000000101111110111000110011011011001, 57'b111101100111110000011000011101000110011100100011001111011,
      57'b111011011001011111001011100011101101100110001100101110010, 57'b111100101100100000000000111010101111101110010001111011111,
      57'b111100111101001001111011100000111101111111001011111010010, 57'b111101111111101110101001110111011000110111001000101100100,
      57'b110100111100011011011101010100101100001110100011010000110, 57'b110011100010001010100111101001100111001010011101100011101,
      57'b111101111111111001110000010011100111000101010011001111001, 57'b111100111001111100101010110001110000001111001100101000010,
      57'b111100101111111100111110010111101111001010110101000010000, 57'b111011010000111010110010101000011101101010000101011000000,
      57'b111101101001101101111110001111011110010111111101111011100, 57'b111101101111001000001011000001111011011011000110110000001,
      57'b111010110110110011001100001100011100010100000110010110110, 57'b111001100011011011001000001010011010111010111010011011101,
      57'b111101111001100110110100001011010001110101010111011110000, 57'b111101011000101100111010000101010010011001010001011110101,
      57'b111100001000010010111001001001000110100001010100101010111, 57'b111100010100000011000101111101111010011010011110010111010,
      57'b111101010000110110010011011010010110000001010011101011110, 57'b111101111100010111010011100110111110010110100101101111000,
      57'b111000101011111110000000010000110010101001100101111011110, 57'b111000000000011101110100010101101011011111011100001011011,
      57'b111101111101111110100011100001111000010101000110110001000, 57'b111101001010010011001000011100011101011000100101001101100,
      57'b111100011100111000010001111100011110101100011000000101001, 57'b111011111101101110101011101011100001001001101001011011110,
      57'b111101011110010110101010011001011000011010010001100100111, 57'b111101110110111011110101101101010000001111000011001010001,
      57'b111010000111000010101101101001110000101110100100111001110, 57'b111010100010000110001000011011100100010010011011011110000,
      57'b111101110010110101001110101010101000001000110011111010011, 57'b111101100101000001000111100011001101110011100010001001001,
      57'b111011100100110010111111111000011100001100101001110001001, 57'b111100100111110011100110000100101110011001010010010000110,
      57'b111101000001010101001110000010011111101010100010111111111, 57'b111101111111010111001110100100101001100000100000100001111,
      57'b110110010000011001001011001110100111011010100010001001101, 57'b110110011100111011001111100010010110001011010001010011001,
      57'b111101111111001111110101010000101010010000010110101100000, 57'b111101000010010110111000100010001101011111000001111111010,
      57'b111100100110100111011110001101101010110001001111101111111, 57'b111011100111100110100101110101110111000011100110100100001,
      57'b111101100100010011111010110000111000000101001110000010011, 57'b111101110011010100110000111000101010111010101001110100111,
      57'b111010011111000111001101111101001011011101100001001110001, 57'b111010001010000100011111011101111110001101001001101111000,
      57'b111101110110100001000001101011110100110011001000000001001, 57'b111101011111001000001101101100001000100010101010011000001,
      57'b111011111010111111101111011100110010101101100110110100011, 57'b111100011110000111100010001001001100000011100010100011000,
      57'b111101001001010101010010000011111110001011010100000010101, 57'b111101111110001010110111000111011011111011001101011110110,
      57'b110111110100011101011011111111101111001001010101000111111, 57'b111000110010001010001101010000011000111011000001100001101,
      57'b111101111100000110000111101001010010000001100011000001100, 57'b111101010001110000001100001001010010110010011101111000110,
      57'b111100010010110000111001101001100101110110111000100010000, 57'b111100001001100111110100111001111111011100010010101001111,
      57'b111101010111110111000111111011000100111110101011110110110, 57'b111101111001111100110101110111100000110111011110001100101,
      57'b111001011101010010110001100110100111100010101110110101101, 57'b111010111001101110110001111001001001001100001000010010010,
      57'b111101101110100011111111011110011100010101001000101011010, 57'b111101101010010110101101100011011000110000111010100100100,
      57'b111011001110000010111110101000100000011011111100111110010, 57'b111100110001000101110010001001111111011000010001011111111,
      57'b111100111000110111010110010010110000011100100000110111111, 57'b111101111111111100001110001101000011100001100101101110111,
      57'b110010101111111010100110100100001111110101011001000100110, 57'b110001111011010100010100101101010101110011001011111001011,
      57'b111101111111111110000100101000011110001010011101111010001, 57'b111100110111110001100101010011001110010010101101101110101,
      57'b111100110010001110001010101000011011111110101001101011011, 57'b111011001011001010101010110110111101010111001010010001111,
      57'b111101101010111110111000101110010100010001000101001111111, 57'b111101101101111111001111001000011100101010111010110011010,
      57'b111010111100101001111010111100110000100111101111110101110, 57'b111001010111001001111000111010101111100111011100110101011,
      57'b111101111010010010010001000000110101111001010101110110100, 57'b111101010111000000110100011110011010001011110110011101111,
      57'b111100001010111100011011011100100110110111110001010111100, 57'b111100010001011110010110101100110001011000001001111100010,
      57'b111101010010101001100100100010000100100001111010100100011, 57'b111101111011110100010100110011100000110100011001000101010,
      57'b111000111000010101111110110001101000010001100010011111111, 57'b110111100111111110101001100111011001100000111110111000001,
      57'b111101111110010110100011100000011100100010100001101010100, 57'b111101001000010110111100101000011010101110101111011111110,
      57'b111100011111010110011001111101010101111100000011010000000, 57'b111011111000010000001100100000110101111111111011111111110,
      57'b111101011111111001001110100100101101000011011000101000111, 57'b111101110110000101100111101001011000110101111011010110010,
      57'b111010001101000101111011111111011111010001111001001000011, 57'b111010011100000111111010111100011010100111011011010101011,
      57'b111101110011110011101101100101001101001010001011001011010, 57'b111101100011100110001010110001001100111101010101011010111,
      57'b111011101010011001101000000101011101010000110000010011101, 57'b111100100101011010111100101010001011001110010001011110001,
      57'b111101000011011000000101000011101100110101010000110010101, 57'b111101111111000111110100100101011111010011101100010000110,
      57'b110110101001011100111011101001010010011010100110100001010, 57'b110110000011110110110000101001110010001100011000001100100,
      57'b111101111111011110000000100000010100000100110000110010001, 57'b111101000000010011000101101110101011011100101001011111010,
      57'b111100101000111111010100000011100110110011001101010100110, 57'b111011100001111110110110101000111001001100011000100101001,
      57'b111101100101101101110001000001010000000001101101010011001, 57'b111101110010010101000110111111111100000011100111001011110,
      57'b111010100101000100101001111010001000110111000001011110011, 57'b111010000100000000100111000000101111010110110011000011110,
      57'b111101110111010110000011101001100010100001010010101000100, 57'b111101011101100100100100110100000101101101100010000001101,
      57'b111100000000001110100000011001000001010111000001011100001, 57'b111100011011101000101001100011011100000010111111110001101,
      57'b111101001011010000011111101000010101111010111111111100001, 57'b111101111101110001101000110001101011001101010110110110111,
      57'b111000000110101100100110110111100101100100110011110000110, 57'b111000100101110001011000101111111011110011111101010001000,
      57'b111101111100100111111000101001111100001011010110000001000, 57'b111101001111111011111010011110001001100010100100111011110,
      57'b111100010101010100111011011101000011110101110101101011000, 57'b111100000110111101101000010111000010010111100010010110110,
      57'b111101011001100010001010110100101111100110111101111110011, 57'b111101111001010000001011111111100010001100000100111001110,
      57'b111001101001100010111011101001101001011001011110111101110, 57'b111010110011110111001010010011100101011010110001111001011,
      57'b111101101111101011110001101101010100110111010010110011100, 57'b111101101001000100101010111000110111001011010010011100001,
      57'b111011010011110010000110011010011110110111111001100011011, 57'b111100101110110011101111011100111001111100011010001011100,
      57'b111100111011000001100010100101100001100000100011101100100, 57'b111101111111110110101010111100100001001011111110110101110,
      57'b110100001010001101000010111011011010000101100000101111111, 57'b110100100011010100011100101101111111110000110000101111001,
      57'b111101111111110010111110001000010000010001100000000010100, 57'b111100111100000101111101100011011100100001011001101011011,
      57'b111100101101101010000101100100110010011110111010001001000, 57'b111011010110101000111001100010010010111001101110000001001,
      57'b111101101000011010110011100101111010110011101001010111001, 57'b111101110000001110110011011011001001010000000111101010100,
      57'b111010110000111010101100101011100100010001100001000000010, 57'b111001101111101010001011000111111000000010000100110011010,
      57'b111101111000111000111101010111110001010000100011100001000, 57'b111101011010010110111010000001001110111100111100100100101,
      57'b111100000101101000000010110000111100011111000010111101100, 57'b111100010110100110011001111010011010011101001101110111000,
      57'b111101001111000001000001011101101101101000010010001110010, 57'b111101111100110111110110101111100111110111101111000101001,
      57'b111000011111100100010111101010111110110110100100010010011, 57'b111000001100111011000100101000000101111100010010011100111,
      57'b111101111101100100000110111000110100000011101010101001101, 57'b111101001100001101010111011110001010001010111010110010100,
      57'b111100011010011000101001001010010110000010100110111100001, 57'b111100000001100101010111001010101111011011011110110010110,
      57'b111101011100110001111101000011111110110010001010101011110, 57'b111101110111101111101011011100101000111001010001111000000,
      57'b111010000000111110001100000000110101110011111110111010010, 57'b111010101000000010110001111011100000110010111000001001000,
      57'b111101110001110100011001111101100011101011100111010000101, 57'b111101100110011001110111000100000110000101101111010100000,
      57'b111011011111001010001010100010111111111111100000011011001, 57'b111100101010001010100111111110101000101011001110111111100,
      57'b111100111111010000011111110000111101100000011011010000110, 57'b111101111111100100001011000010100111000010011000111101101,
      57'b110101101110101000000011011111001100000001000111011001001, 57'b110110110101111110001101100111110011110011011000100101001,
      57'b111101111110111111001100100100010111101110011001100000111, 57'b111101000100011000110011011100111010010000001101110100001,
      57'b111100100100001110000001100110000011000001001000111111111, 57'b111011101101001100000110001011100111110100001000011011001,
      57'b111101100010110111110111101011001111111101111100001011010, 57'b111101110100010010000100101011011101011010110000000100101,
      57'b111010011001001000001111110110110001110001011101010101111, 57'b111010010000000111000010110000011110101110010011110111110,
      57'b111101110101101001100111101010001010110111000100000010001, 57'b111101100000101001101100111011100010001100101111001010111,
      57'b111011110101100000000011010010101111100100101011000100000, 57'b111100100000100100111001001100110001111010001000010001100,
      57'b111101000111011000001000010011011010010000110110001001001, 57'b111101111110100001101000101011000110110000110000010000111,
      57'b110111011011011111010011011101100001110001111011001001100, 57'b111000111110100001010011110111011110100101100101100011100,
      57'b111101111011100001111011001000011010010110111111010110111, 57'b111101010011100010011100011011110100111010110000011110101,
      57'b111100010000001011011101010100001011101010110000011010110, 57'b111100001100010000101100100011111001110100100011011100101,
      57'b111101010110001001111111110111101001111101111101011001000, 57'b111101111010100111000101100011111101011110010110100000111,
      57'b111001010001000000011111000011011000110000011000111011010, 57'b111010111111100100100110111010011011100110100000111100100,
      57'b111101101101011001111010000101100111001101000101010111001, 57'b111101101011100110011111101010000100011000000110111111111,
      57'b111011001000010001110111110000001111011110111101111010001, 57'b111100110011010110000111100111111010100101011001110000110,
      57'b111100110110101011010111111101111010010101010111111001101, 57'b111101111111111111010011100101100100101111000110001001111,
      57'b110000010110110010110101100001110010100001001011100000011, 57'b110000010110110010110101100001110010100001001011100000011,
      57'b111101111111111111010011100101100100101111000110001001111, 57'b111100110110101011010111111101111010010101010111111001101,
      57'b111100110011010110000111100111111010100101011001110000110, 57'b111011001000010001110111110000001111011110111101111010001,
      57'b111101101011100110011111101010000100011000000110111111111, 57'b111101101101011001111010000101100111001101000101010111001,
      57'b111010111111100100100110111010011011100110100000111100100, 57'b111001010001000000011111000011011000110000011000111011010,
      57'b111101111010100111000101100011111101011110010110100000111, 57'b111101010110001001111111110111101001111101111101011001000,
      57'b111100001100010000101100100011111001110100100011011100101, 57'b111100010000001011011101010100001011101010110000011010110,
      57'b111101010011100010011100011011110100111010110000011110101, 57'b111101111011100001111011001000011010010110111111010110111,
      57'b111000111110100001010011110111011110100101100101100011100, 57'b110111011011011111010011011101100001110001111011001001100,
      57'b111101111110100001101000101011000110110000110000010000111, 57'b111101000111011000001000010011011010010000110110001001001,
      57'b111100100000100100111001001100110001111010001000010001100, 57'b111011110101100000000011010010101111100100101011000100000,
      57'b111101100000101001101100111011100010001100101111001010111, 57'b111101110101101001100111101010001010110111000100000010001,
      57'b111010010000000111000010110000011110101110010011110111110, 57'b111010011001001000001111110110110001110001011101010101111,
      57'b111101110100010010000100101011011101011010110000000100101, 57'b111101100010110111110111101011001111111101111100001011010,
      57'b111011101101001100000110001011100111110100001000011011001, 57'b111100100100001110000001100110000011000001001000111111111,
      57'b111101000100011000110011011100111010010000001101110100001, 57'b111101111110111111001100100100010111101110011001100000111,
      57'b110110110101111110001101100111110011110011011000100101001, 57'b110101101110101000000011011111001100000001000111011001001,
      57'b111101111111100100001011000010100111000010011000111101101, 57'b111100111111010000011111110000111101100000011011010000110,
      57'b111100101010001010100111111110101000101011001110111111100, 57'b111011011111001010001010100010111111111111100000011011001,
      57'b111101100110011001110111000100000110000101101111010100000, 57'b111101110001110100011001111101100011101011100111010000101,
      57'b111010101000000010110001111011100000110010111000001001000, 57'b111010000000111110001100000000110101110011111110111010010,
      57'b111101110111101111101011011100101000111001010001111000000, 57'b111101011100110001111101000011111110110010001010101011110,
      57'b111100000001100101010111001010101111011011011110110010110, 57'b111100011010011000101001001010010110000010100110111100001,
      57'b111101001100001101010111011110001010001010111010110010100, 57'b111101111101100100000110111000110100000011101010101001101,
      57'b111000001100111011000100101000000101111100010010011100111, 57'b111000011111100100010111101010111110110110100100010010011,
      57'b111101111100110111110110101111100111110111101111000101001, 57'b111101001111000001000001011101101101101000010010001110010,
      57'b111100010110100110011001111010011010011101001101110111000, 57'b111100000101101000000010110000111100011111000010111101100,
      57'b111101011010010110111010000001001110111100111100100100101, 57'b111101111000111000111101010111110001010000100011100001000,
      57'b111001101111101010001011000111111000000010000100110011010, 57'b111010110000111010101100101011100100010001100001000000010,
      57'b111101110000001110110011011011001001010000000111101010100, 57'b111101101000011010110011100101111010110011101001010111001,
      57'b111011010110101000111001100010010010111001101110000001001, 57'b111100101101101010000101100100110010011110111010001001000,
      57'b111100111100000101111101100011011100100001011001101011011, 57'b111101111111110010111110001000010000010001100000000010100,
      57'b110100100011010100011100101101111111110000110000101111001, 57'b110100001010001101000010111011011010000101100000101111111,
      57'b111101111111110110101010111100100001001011111110110101110, 57'b111100111011000001100010100101100001100000100011101100100,
      57'b111100101110110011101111011100111001111100011010001011100, 57'b111011010011110010000110011010011110110111111001100011011,
      57'b111101101001000100101010111000110111001011010010011100001, 57'b111101101111101011110001101101010100110111010010110011100,
      57'b111010110011110111001010010011100101011010110001111001011, 57'b111001101001100010111011101001101001011001011110111101110,
      57'b111101111001010000001011111111100010001100000100111001110, 57'b111101011001100010001010110100101111100110111101111110011,
      57'b111100000110111101101000010111000010010111100010010110110, 57'b111100010101010100111011011101000011110101110101101011000,
      57'b111101001111111011111010011110001001100010100100111011110, 57'b111101111100100111111000101001111100001011010110000001000,
      57'b111000100101110001011000101111111011110011111101010001000, 57'b111000000110101100100110110111100101100100110011110000110,
      57'b111101111101110001101000110001101011001101010110110110111, 57'b111101001011010000011111101000010101111010111111111100001,
      57'b111100011011101000101001100011011100000010111111110001101, 57'b111100000000001110100000011001000001010111000001011100001,
      57'b111101011101100100100100110100000101101101100010000001101, 57'b111101110111010110000011101001100010100001010010101000100,
      57'b111010000100000000100111000000101111010110110011000011110, 57'b111010100101000100101001111010001000110111000001011110011,
      57'b111101110010010101000110111111111100000011100111001011110, 57'b111101100101101101110001000001010000000001101101010011001,
      57'b111011100001111110110110101000111001001100011000100101001, 57'b111100101000111111010100000011100110110011001101010100110,
      57'b111101000000010011000101101110101011011100101001011111010, 57'b111101111111011110000000100000010100000100110000110010001,
      57'b110110000011110110110000101001110010001100011000001100100, 57'b110110101001011100111011101001010010011010100110100001010,
      57'b111101111111000111110100100101011111010011101100010000110, 57'b111101000011011000000101000011101100110101010000110010101,
      57'b111100100101011010111100101010001011001110010001011110001, 57'b111011101010011001101000000101011101010000110000010011101,
      57'b111101100011100110001010110001001100111101010101011010111, 57'b111101110011110011101101100101001101001010001011001011010,
      57'b111010011100000111111010111100011010100111011011010101011, 57'b111010001101000101111011111111011111010001111001001000011,
      57'b111101110110000101100111101001011000110101111011010110010, 57'b111101011111111001001110100100101101000011011000101000111,
      57'b111011111000010000001100100000110101111111111011111111110, 57'b111100011111010110011001111101010101111100000011010000000,
      57'b111101001000010110111100101000011010101110101111011111110, 57'b111101111110010110100011100000011100100010100001101010100,
      57'b110111100111111110101001100111011001100000111110111000001, 57'b111000111000010101111110110001101000010001100010011111111,
      57'b111101111011110100010100110011100000110100011001000101010, 57'b111101010010101001100100100010000100100001111010100100011,
      57'b111100010001011110010110101100110001011000001001111100010, 57'b111100001010111100011011011100100110110111110001010111100,
      57'b111101010111000000110100011110011010001011110110011101111, 57'b111101111010010010010001000000110101111001010101110110100,
      57'b111001010111001001111000111010101111100111011100110101011, 57'b111010111100101001111010111100110000100111101111110101110,
      57'b111101101101111111001111001000011100101010111010110011010, 57'b111101101010111110111000101110010100010001000101001111111,
      57'b111011001011001010101010110110111101010111001010010001111, 57'b111100110010001110001010101000011011111110101001101011011,
      57'b111100110111110001100101010011001110010010101101101110101, 57'b111101111111111110000100101000011110001010011101111010001,
      57'b110001111011010100010100101101010101110011001011111001011, 57'b110010101111111010100110100100001111110101011001000100110,
      57'b111101111111111100001110001101000011100001100101101110111, 57'b111100111000110111010110010010110000011100100000110111111,
      57'b111100110001000101110010001001111111011000010001011111111, 57'b111011001110000010111110101000100000011011111100111110010,
      57'b111101101010010110101101100011011000110000111010100100100, 57'b111101101110100011111111011110011100010101001000101011010,
      57'b111010111001101110110001111001001001001100001000010010010, 57'b111001011101010010110001100110100111100010101110110101101,
      57'b111101111001111100110101110111100000110111011110001100101, 57'b111101010111110111000111111011000100111110101011110110110,
      57'b111100001001100111110100111001111111011100010010101001111, 57'b111100010010110000111001101001100101110110111000100010000,
      57'b111101010001110000001100001001010010110010011101111000110, 57'b111101111100000110000111101001010010000001100011000001100,
      57'b111000110010001010001101010000011000111011000001100001101, 57'b110111110100011101011011111111101111001001010101000111111,
      57'b111101111110001010110111000111011011111011001101011110110, 57'b111101001001010101010010000011111110001011010100000010101,
      57'b111100011110000111100010001001001100000011100010100011000, 57'b111011111010111111101111011100110010101101100110110100011,
      57'b111101011111001000001101101100001000100010101010011000001, 57'b111101110110100001000001101011110100110011001000000001001,
      57'b111010001010000100011111011101111110001101001001101111000, 57'b111010011111000111001101111101001011011101100001001110001,
      57'b111101110011010100110000111000101010111010101001110100111, 57'b111101100100010011111010110000111000000101001110000010011,
      57'b111011100111100110100101110101110111000011100110100100001, 57'b111100100110100111011110001101101010110001001111101111111,
      57'b111101000010010110111000100010001101011111000001111111010, 57'b111101111111001111110101010000101010010000010110101100000,
      57'b110110011100111011001111100010010110001011010001010011001, 57'b110110010000011001001011001110100111011010100010001001101,
      57'b111101111111010111001110100100101001100000100000100001111, 57'b111101000001010101001110000010011111101010100010111111111,
      57'b111100100111110011100110000100101110011001010010010000110, 57'b111011100100110010111111111000011100001100101001110001001,
      57'b111101100101000001000111100011001101110011100010001001001, 57'b111101110010110101001110101010101000001000110011111010011,
      57'b111010100010000110001000011011100100010010011011011110000, 57'b111010000111000010101101101001110000101110100100111001110,
      57'b111101110110111011110101101101010000001111000011001010001, 57'b111101011110010110101010011001011000011010010001100100111,
      57'b111011111101101110101011101011100001001001101001011011110, 57'b111100011100111000010001111100011110101100011000000101001,
      57'b111101001010010011001000011100011101011000100101001101100, 57'b111101111101111110100011100001111000010101000110110001000,
      57'b111000000000011101110100010101101011011111011100001011011, 57'b111000101011111110000000010000110010101001100101111011110,
      57'b111101111100010111010011100110111110010110100101101111000, 57'b111101010000110110010011011010010110000001010011101011110,
      57'b111100010100000011000101111101111010011010011110010111010, 57'b111100001000010010111001001001000110100001010100101010111,
      57'b111101011000101100111010000101010010011001010001011110101, 57'b111101111001100110110100001011010001110101010111011110000,
      57'b111001100011011011001000001010011010111010111010011011101, 57'b111010110110110011001100001100011100010100000110010110110,
      57'b111101101111001000001011000001111011011011000110110000001, 57'b111101101001101101111110001111011110010111111101111011100,
      57'b111011010000111010110010101000011101101010000101011000000, 57'b111100101111111100111110010111101111001010110101000010000,
      57'b111100111001111100101010110001110000001111001100101000010, 57'b111101111111111001110000010011100111000101010011001111001,
      57'b110011100010001010100111101001100111001010011101100011101, 57'b110100111100011011011101010100101100001110100011010000110,
      57'b111101111111101110101001110111011000110111001000101100100, 57'b111100111101001001111011100000111101111111001011111010010,
      57'b111100101100100000000000111010101111101110010001111011111, 57'b111011011001011111001011100011101101100110001100101110010,
      57'b111101100111110000011000011101000110011100100011001111011, 57'b111101110000110001010000000101111110111000110011011011001,
      57'b111010101101111101110011110001011100111011011001110110110, 57'b111001110101110000110101101000110001011011110001101001000,
      57'b111101111000100001001000010111100100010011000111101011111, 57'b111101011011001011000111100010100111111011011110001000111,
      57'b111100000100010010001000100100000001100101011000010001100, 57'b111100010111110111100001001001011010001000001000000010101,
      57'b111101001110000101101000100010000111100000111010111000010, 57'b111101111101000111001101110101100011110100001011110010001,
      57'b111000011001010110111101111111001010001010001011010100111, 57'b111000010011001001001100101001101111111010011010000001001,
      57'b111101111101010101111101111001011000011001111110111011100, 57'b111101001101001001101111110100100001010110000011010110010,
      57'b111100011001001000010000111101100010010011010011000011111, 57'b111100000010111011111001111101100001100011011100010110111,
      57'b111101011011111110110011010000110111001111001001011101001, 57'b111101111000001000101101000010100110011110111001110001100,
      57'b111001111011110110111010010000000101111010011100000000010, 57'b111010101011000000100000000010010111101000110011110110100,
      57'b111101110001010011000111101000100001110010001100101111010, 57'b111101100111000101011001100100111100110011010000001100000,
      57'b111011011100010100111100000010100111111010101011010010011, 57'b111100101011010101100001101010001100101110110010010011111,
      57'b111100111110001101011100010011100111000101101001100110011, 57'b111101111111101001101110001010100101100011011111011010011,
      57'b110101010101100010000000110111101010111111000001100010111, 57'b110111000010011111000011100010010110000010011000010100001,
      57'b111101111110110101111101001110101000101000101001110001100, 57'b111101000101011001000011100011110110111100001110110001000,
      57'b111100100011000000101101001101001001010110011001010100010, 57'b111011101111111101111111101100110101010010100000111011110,
      57'b111101100010001001000001100110001010000011100000000000100, 57'b111101110100101111110110000110110000000010110101100110000,
      57'b111010010110001000001101001001110100101010100010100100000, 57'b111010010011000111110011010011001010101010101010010111010,
      57'b111101110101001101000001110010011111001100101100000000000, 57'b111101100001011001101000101001001001100011110001111110001,
      57'b111011110010101111010100001101101001111001101100000100101, 57'b111100100001110010111111101011011001010100100001110000000,
      57'b111101000110011000110101001110101000110000100011001010101, 57'b111101111110101100000110100101101101001110101110010011110,
      57'b110111001110111111011011011101011001001001010100001011100, 57'b111001000100101100001011100100111110001000001100000000100,
      57'b111101111011001110111010101010110100010000011110011101110, 57'b111101010100011010110011101101110010101000101101011010010,
      57'b111100001110111000001101101100100110111000100100001110010, 57'b111100001101100100101000000010111000100110111001110111111,
      57'b111101010101010010101010001111010001011001011100110001110, 57'b111101111010111011010011011101101010000110110100001011101,
      57'b111001001010110110100100111101001101101100010101011111010, 57'b111011000010011110110101010101010111100111001000000111111,
      57'b111101101100110100000000011011101100010110011110101000110, 57'b111101101100001101100010010000100010001011010010001001111,
      57'b111011000101011000100101110000110110101011110110101000100, 57'b111100110100011101101000111101010101000011001110001110001,
      57'b111100110101100100101110011101101001011111110001010011100, 57'b111101111111111111111011000100001011000100001110100000010,
      57'b101101001001000011111100010111110110011001010010010111010, I_1);
  assign O_1 = signext_62_57(r_ac_ieee_float_base_slc_gm_im_tab_d_rom_1_BUTTERFLY_if_r_ac_ieee_float_base_mux_nl);

  function automatic [56:0] MUX_v_57_1024_2;
    input [56:0] input_0;
    input [56:0] input_1;
    input [56:0] input_2;
    input [56:0] input_3;
    input [56:0] input_4;
    input [56:0] input_5;
    input [56:0] input_6;
    input [56:0] input_7;
    input [56:0] input_8;
    input [56:0] input_9;
    input [56:0] input_10;
    input [56:0] input_11;
    input [56:0] input_12;
    input [56:0] input_13;
    input [56:0] input_14;
    input [56:0] input_15;
    input [56:0] input_16;
    input [56:0] input_17;
    input [56:0] input_18;
    input [56:0] input_19;
    input [56:0] input_20;
    input [56:0] input_21;
    input [56:0] input_22;
    input [56:0] input_23;
    input [56:0] input_24;
    input [56:0] input_25;
    input [56:0] input_26;
    input [56:0] input_27;
    input [56:0] input_28;
    input [56:0] input_29;
    input [56:0] input_30;
    input [56:0] input_31;
    input [56:0] input_32;
    input [56:0] input_33;
    input [56:0] input_34;
    input [56:0] input_35;
    input [56:0] input_36;
    input [56:0] input_37;
    input [56:0] input_38;
    input [56:0] input_39;
    input [56:0] input_40;
    input [56:0] input_41;
    input [56:0] input_42;
    input [56:0] input_43;
    input [56:0] input_44;
    input [56:0] input_45;
    input [56:0] input_46;
    input [56:0] input_47;
    input [56:0] input_48;
    input [56:0] input_49;
    input [56:0] input_50;
    input [56:0] input_51;
    input [56:0] input_52;
    input [56:0] input_53;
    input [56:0] input_54;
    input [56:0] input_55;
    input [56:0] input_56;
    input [56:0] input_57;
    input [56:0] input_58;
    input [56:0] input_59;
    input [56:0] input_60;
    input [56:0] input_61;
    input [56:0] input_62;
    input [56:0] input_63;
    input [56:0] input_64;
    input [56:0] input_65;
    input [56:0] input_66;
    input [56:0] input_67;
    input [56:0] input_68;
    input [56:0] input_69;
    input [56:0] input_70;
    input [56:0] input_71;
    input [56:0] input_72;
    input [56:0] input_73;
    input [56:0] input_74;
    input [56:0] input_75;
    input [56:0] input_76;
    input [56:0] input_77;
    input [56:0] input_78;
    input [56:0] input_79;
    input [56:0] input_80;
    input [56:0] input_81;
    input [56:0] input_82;
    input [56:0] input_83;
    input [56:0] input_84;
    input [56:0] input_85;
    input [56:0] input_86;
    input [56:0] input_87;
    input [56:0] input_88;
    input [56:0] input_89;
    input [56:0] input_90;
    input [56:0] input_91;
    input [56:0] input_92;
    input [56:0] input_93;
    input [56:0] input_94;
    input [56:0] input_95;
    input [56:0] input_96;
    input [56:0] input_97;
    input [56:0] input_98;
    input [56:0] input_99;
    input [56:0] input_100;
    input [56:0] input_101;
    input [56:0] input_102;
    input [56:0] input_103;
    input [56:0] input_104;
    input [56:0] input_105;
    input [56:0] input_106;
    input [56:0] input_107;
    input [56:0] input_108;
    input [56:0] input_109;
    input [56:0] input_110;
    input [56:0] input_111;
    input [56:0] input_112;
    input [56:0] input_113;
    input [56:0] input_114;
    input [56:0] input_115;
    input [56:0] input_116;
    input [56:0] input_117;
    input [56:0] input_118;
    input [56:0] input_119;
    input [56:0] input_120;
    input [56:0] input_121;
    input [56:0] input_122;
    input [56:0] input_123;
    input [56:0] input_124;
    input [56:0] input_125;
    input [56:0] input_126;
    input [56:0] input_127;
    input [56:0] input_128;
    input [56:0] input_129;
    input [56:0] input_130;
    input [56:0] input_131;
    input [56:0] input_132;
    input [56:0] input_133;
    input [56:0] input_134;
    input [56:0] input_135;
    input [56:0] input_136;
    input [56:0] input_137;
    input [56:0] input_138;
    input [56:0] input_139;
    input [56:0] input_140;
    input [56:0] input_141;
    input [56:0] input_142;
    input [56:0] input_143;
    input [56:0] input_144;
    input [56:0] input_145;
    input [56:0] input_146;
    input [56:0] input_147;
    input [56:0] input_148;
    input [56:0] input_149;
    input [56:0] input_150;
    input [56:0] input_151;
    input [56:0] input_152;
    input [56:0] input_153;
    input [56:0] input_154;
    input [56:0] input_155;
    input [56:0] input_156;
    input [56:0] input_157;
    input [56:0] input_158;
    input [56:0] input_159;
    input [56:0] input_160;
    input [56:0] input_161;
    input [56:0] input_162;
    input [56:0] input_163;
    input [56:0] input_164;
    input [56:0] input_165;
    input [56:0] input_166;
    input [56:0] input_167;
    input [56:0] input_168;
    input [56:0] input_169;
    input [56:0] input_170;
    input [56:0] input_171;
    input [56:0] input_172;
    input [56:0] input_173;
    input [56:0] input_174;
    input [56:0] input_175;
    input [56:0] input_176;
    input [56:0] input_177;
    input [56:0] input_178;
    input [56:0] input_179;
    input [56:0] input_180;
    input [56:0] input_181;
    input [56:0] input_182;
    input [56:0] input_183;
    input [56:0] input_184;
    input [56:0] input_185;
    input [56:0] input_186;
    input [56:0] input_187;
    input [56:0] input_188;
    input [56:0] input_189;
    input [56:0] input_190;
    input [56:0] input_191;
    input [56:0] input_192;
    input [56:0] input_193;
    input [56:0] input_194;
    input [56:0] input_195;
    input [56:0] input_196;
    input [56:0] input_197;
    input [56:0] input_198;
    input [56:0] input_199;
    input [56:0] input_200;
    input [56:0] input_201;
    input [56:0] input_202;
    input [56:0] input_203;
    input [56:0] input_204;
    input [56:0] input_205;
    input [56:0] input_206;
    input [56:0] input_207;
    input [56:0] input_208;
    input [56:0] input_209;
    input [56:0] input_210;
    input [56:0] input_211;
    input [56:0] input_212;
    input [56:0] input_213;
    input [56:0] input_214;
    input [56:0] input_215;
    input [56:0] input_216;
    input [56:0] input_217;
    input [56:0] input_218;
    input [56:0] input_219;
    input [56:0] input_220;
    input [56:0] input_221;
    input [56:0] input_222;
    input [56:0] input_223;
    input [56:0] input_224;
    input [56:0] input_225;
    input [56:0] input_226;
    input [56:0] input_227;
    input [56:0] input_228;
    input [56:0] input_229;
    input [56:0] input_230;
    input [56:0] input_231;
    input [56:0] input_232;
    input [56:0] input_233;
    input [56:0] input_234;
    input [56:0] input_235;
    input [56:0] input_236;
    input [56:0] input_237;
    input [56:0] input_238;
    input [56:0] input_239;
    input [56:0] input_240;
    input [56:0] input_241;
    input [56:0] input_242;
    input [56:0] input_243;
    input [56:0] input_244;
    input [56:0] input_245;
    input [56:0] input_246;
    input [56:0] input_247;
    input [56:0] input_248;
    input [56:0] input_249;
    input [56:0] input_250;
    input [56:0] input_251;
    input [56:0] input_252;
    input [56:0] input_253;
    input [56:0] input_254;
    input [56:0] input_255;
    input [56:0] input_256;
    input [56:0] input_257;
    input [56:0] input_258;
    input [56:0] input_259;
    input [56:0] input_260;
    input [56:0] input_261;
    input [56:0] input_262;
    input [56:0] input_263;
    input [56:0] input_264;
    input [56:0] input_265;
    input [56:0] input_266;
    input [56:0] input_267;
    input [56:0] input_268;
    input [56:0] input_269;
    input [56:0] input_270;
    input [56:0] input_271;
    input [56:0] input_272;
    input [56:0] input_273;
    input [56:0] input_274;
    input [56:0] input_275;
    input [56:0] input_276;
    input [56:0] input_277;
    input [56:0] input_278;
    input [56:0] input_279;
    input [56:0] input_280;
    input [56:0] input_281;
    input [56:0] input_282;
    input [56:0] input_283;
    input [56:0] input_284;
    input [56:0] input_285;
    input [56:0] input_286;
    input [56:0] input_287;
    input [56:0] input_288;
    input [56:0] input_289;
    input [56:0] input_290;
    input [56:0] input_291;
    input [56:0] input_292;
    input [56:0] input_293;
    input [56:0] input_294;
    input [56:0] input_295;
    input [56:0] input_296;
    input [56:0] input_297;
    input [56:0] input_298;
    input [56:0] input_299;
    input [56:0] input_300;
    input [56:0] input_301;
    input [56:0] input_302;
    input [56:0] input_303;
    input [56:0] input_304;
    input [56:0] input_305;
    input [56:0] input_306;
    input [56:0] input_307;
    input [56:0] input_308;
    input [56:0] input_309;
    input [56:0] input_310;
    input [56:0] input_311;
    input [56:0] input_312;
    input [56:0] input_313;
    input [56:0] input_314;
    input [56:0] input_315;
    input [56:0] input_316;
    input [56:0] input_317;
    input [56:0] input_318;
    input [56:0] input_319;
    input [56:0] input_320;
    input [56:0] input_321;
    input [56:0] input_322;
    input [56:0] input_323;
    input [56:0] input_324;
    input [56:0] input_325;
    input [56:0] input_326;
    input [56:0] input_327;
    input [56:0] input_328;
    input [56:0] input_329;
    input [56:0] input_330;
    input [56:0] input_331;
    input [56:0] input_332;
    input [56:0] input_333;
    input [56:0] input_334;
    input [56:0] input_335;
    input [56:0] input_336;
    input [56:0] input_337;
    input [56:0] input_338;
    input [56:0] input_339;
    input [56:0] input_340;
    input [56:0] input_341;
    input [56:0] input_342;
    input [56:0] input_343;
    input [56:0] input_344;
    input [56:0] input_345;
    input [56:0] input_346;
    input [56:0] input_347;
    input [56:0] input_348;
    input [56:0] input_349;
    input [56:0] input_350;
    input [56:0] input_351;
    input [56:0] input_352;
    input [56:0] input_353;
    input [56:0] input_354;
    input [56:0] input_355;
    input [56:0] input_356;
    input [56:0] input_357;
    input [56:0] input_358;
    input [56:0] input_359;
    input [56:0] input_360;
    input [56:0] input_361;
    input [56:0] input_362;
    input [56:0] input_363;
    input [56:0] input_364;
    input [56:0] input_365;
    input [56:0] input_366;
    input [56:0] input_367;
    input [56:0] input_368;
    input [56:0] input_369;
    input [56:0] input_370;
    input [56:0] input_371;
    input [56:0] input_372;
    input [56:0] input_373;
    input [56:0] input_374;
    input [56:0] input_375;
    input [56:0] input_376;
    input [56:0] input_377;
    input [56:0] input_378;
    input [56:0] input_379;
    input [56:0] input_380;
    input [56:0] input_381;
    input [56:0] input_382;
    input [56:0] input_383;
    input [56:0] input_384;
    input [56:0] input_385;
    input [56:0] input_386;
    input [56:0] input_387;
    input [56:0] input_388;
    input [56:0] input_389;
    input [56:0] input_390;
    input [56:0] input_391;
    input [56:0] input_392;
    input [56:0] input_393;
    input [56:0] input_394;
    input [56:0] input_395;
    input [56:0] input_396;
    input [56:0] input_397;
    input [56:0] input_398;
    input [56:0] input_399;
    input [56:0] input_400;
    input [56:0] input_401;
    input [56:0] input_402;
    input [56:0] input_403;
    input [56:0] input_404;
    input [56:0] input_405;
    input [56:0] input_406;
    input [56:0] input_407;
    input [56:0] input_408;
    input [56:0] input_409;
    input [56:0] input_410;
    input [56:0] input_411;
    input [56:0] input_412;
    input [56:0] input_413;
    input [56:0] input_414;
    input [56:0] input_415;
    input [56:0] input_416;
    input [56:0] input_417;
    input [56:0] input_418;
    input [56:0] input_419;
    input [56:0] input_420;
    input [56:0] input_421;
    input [56:0] input_422;
    input [56:0] input_423;
    input [56:0] input_424;
    input [56:0] input_425;
    input [56:0] input_426;
    input [56:0] input_427;
    input [56:0] input_428;
    input [56:0] input_429;
    input [56:0] input_430;
    input [56:0] input_431;
    input [56:0] input_432;
    input [56:0] input_433;
    input [56:0] input_434;
    input [56:0] input_435;
    input [56:0] input_436;
    input [56:0] input_437;
    input [56:0] input_438;
    input [56:0] input_439;
    input [56:0] input_440;
    input [56:0] input_441;
    input [56:0] input_442;
    input [56:0] input_443;
    input [56:0] input_444;
    input [56:0] input_445;
    input [56:0] input_446;
    input [56:0] input_447;
    input [56:0] input_448;
    input [56:0] input_449;
    input [56:0] input_450;
    input [56:0] input_451;
    input [56:0] input_452;
    input [56:0] input_453;
    input [56:0] input_454;
    input [56:0] input_455;
    input [56:0] input_456;
    input [56:0] input_457;
    input [56:0] input_458;
    input [56:0] input_459;
    input [56:0] input_460;
    input [56:0] input_461;
    input [56:0] input_462;
    input [56:0] input_463;
    input [56:0] input_464;
    input [56:0] input_465;
    input [56:0] input_466;
    input [56:0] input_467;
    input [56:0] input_468;
    input [56:0] input_469;
    input [56:0] input_470;
    input [56:0] input_471;
    input [56:0] input_472;
    input [56:0] input_473;
    input [56:0] input_474;
    input [56:0] input_475;
    input [56:0] input_476;
    input [56:0] input_477;
    input [56:0] input_478;
    input [56:0] input_479;
    input [56:0] input_480;
    input [56:0] input_481;
    input [56:0] input_482;
    input [56:0] input_483;
    input [56:0] input_484;
    input [56:0] input_485;
    input [56:0] input_486;
    input [56:0] input_487;
    input [56:0] input_488;
    input [56:0] input_489;
    input [56:0] input_490;
    input [56:0] input_491;
    input [56:0] input_492;
    input [56:0] input_493;
    input [56:0] input_494;
    input [56:0] input_495;
    input [56:0] input_496;
    input [56:0] input_497;
    input [56:0] input_498;
    input [56:0] input_499;
    input [56:0] input_500;
    input [56:0] input_501;
    input [56:0] input_502;
    input [56:0] input_503;
    input [56:0] input_504;
    input [56:0] input_505;
    input [56:0] input_506;
    input [56:0] input_507;
    input [56:0] input_508;
    input [56:0] input_509;
    input [56:0] input_510;
    input [56:0] input_511;
    input [56:0] input_512;
    input [56:0] input_513;
    input [56:0] input_514;
    input [56:0] input_515;
    input [56:0] input_516;
    input [56:0] input_517;
    input [56:0] input_518;
    input [56:0] input_519;
    input [56:0] input_520;
    input [56:0] input_521;
    input [56:0] input_522;
    input [56:0] input_523;
    input [56:0] input_524;
    input [56:0] input_525;
    input [56:0] input_526;
    input [56:0] input_527;
    input [56:0] input_528;
    input [56:0] input_529;
    input [56:0] input_530;
    input [56:0] input_531;
    input [56:0] input_532;
    input [56:0] input_533;
    input [56:0] input_534;
    input [56:0] input_535;
    input [56:0] input_536;
    input [56:0] input_537;
    input [56:0] input_538;
    input [56:0] input_539;
    input [56:0] input_540;
    input [56:0] input_541;
    input [56:0] input_542;
    input [56:0] input_543;
    input [56:0] input_544;
    input [56:0] input_545;
    input [56:0] input_546;
    input [56:0] input_547;
    input [56:0] input_548;
    input [56:0] input_549;
    input [56:0] input_550;
    input [56:0] input_551;
    input [56:0] input_552;
    input [56:0] input_553;
    input [56:0] input_554;
    input [56:0] input_555;
    input [56:0] input_556;
    input [56:0] input_557;
    input [56:0] input_558;
    input [56:0] input_559;
    input [56:0] input_560;
    input [56:0] input_561;
    input [56:0] input_562;
    input [56:0] input_563;
    input [56:0] input_564;
    input [56:0] input_565;
    input [56:0] input_566;
    input [56:0] input_567;
    input [56:0] input_568;
    input [56:0] input_569;
    input [56:0] input_570;
    input [56:0] input_571;
    input [56:0] input_572;
    input [56:0] input_573;
    input [56:0] input_574;
    input [56:0] input_575;
    input [56:0] input_576;
    input [56:0] input_577;
    input [56:0] input_578;
    input [56:0] input_579;
    input [56:0] input_580;
    input [56:0] input_581;
    input [56:0] input_582;
    input [56:0] input_583;
    input [56:0] input_584;
    input [56:0] input_585;
    input [56:0] input_586;
    input [56:0] input_587;
    input [56:0] input_588;
    input [56:0] input_589;
    input [56:0] input_590;
    input [56:0] input_591;
    input [56:0] input_592;
    input [56:0] input_593;
    input [56:0] input_594;
    input [56:0] input_595;
    input [56:0] input_596;
    input [56:0] input_597;
    input [56:0] input_598;
    input [56:0] input_599;
    input [56:0] input_600;
    input [56:0] input_601;
    input [56:0] input_602;
    input [56:0] input_603;
    input [56:0] input_604;
    input [56:0] input_605;
    input [56:0] input_606;
    input [56:0] input_607;
    input [56:0] input_608;
    input [56:0] input_609;
    input [56:0] input_610;
    input [56:0] input_611;
    input [56:0] input_612;
    input [56:0] input_613;
    input [56:0] input_614;
    input [56:0] input_615;
    input [56:0] input_616;
    input [56:0] input_617;
    input [56:0] input_618;
    input [56:0] input_619;
    input [56:0] input_620;
    input [56:0] input_621;
    input [56:0] input_622;
    input [56:0] input_623;
    input [56:0] input_624;
    input [56:0] input_625;
    input [56:0] input_626;
    input [56:0] input_627;
    input [56:0] input_628;
    input [56:0] input_629;
    input [56:0] input_630;
    input [56:0] input_631;
    input [56:0] input_632;
    input [56:0] input_633;
    input [56:0] input_634;
    input [56:0] input_635;
    input [56:0] input_636;
    input [56:0] input_637;
    input [56:0] input_638;
    input [56:0] input_639;
    input [56:0] input_640;
    input [56:0] input_641;
    input [56:0] input_642;
    input [56:0] input_643;
    input [56:0] input_644;
    input [56:0] input_645;
    input [56:0] input_646;
    input [56:0] input_647;
    input [56:0] input_648;
    input [56:0] input_649;
    input [56:0] input_650;
    input [56:0] input_651;
    input [56:0] input_652;
    input [56:0] input_653;
    input [56:0] input_654;
    input [56:0] input_655;
    input [56:0] input_656;
    input [56:0] input_657;
    input [56:0] input_658;
    input [56:0] input_659;
    input [56:0] input_660;
    input [56:0] input_661;
    input [56:0] input_662;
    input [56:0] input_663;
    input [56:0] input_664;
    input [56:0] input_665;
    input [56:0] input_666;
    input [56:0] input_667;
    input [56:0] input_668;
    input [56:0] input_669;
    input [56:0] input_670;
    input [56:0] input_671;
    input [56:0] input_672;
    input [56:0] input_673;
    input [56:0] input_674;
    input [56:0] input_675;
    input [56:0] input_676;
    input [56:0] input_677;
    input [56:0] input_678;
    input [56:0] input_679;
    input [56:0] input_680;
    input [56:0] input_681;
    input [56:0] input_682;
    input [56:0] input_683;
    input [56:0] input_684;
    input [56:0] input_685;
    input [56:0] input_686;
    input [56:0] input_687;
    input [56:0] input_688;
    input [56:0] input_689;
    input [56:0] input_690;
    input [56:0] input_691;
    input [56:0] input_692;
    input [56:0] input_693;
    input [56:0] input_694;
    input [56:0] input_695;
    input [56:0] input_696;
    input [56:0] input_697;
    input [56:0] input_698;
    input [56:0] input_699;
    input [56:0] input_700;
    input [56:0] input_701;
    input [56:0] input_702;
    input [56:0] input_703;
    input [56:0] input_704;
    input [56:0] input_705;
    input [56:0] input_706;
    input [56:0] input_707;
    input [56:0] input_708;
    input [56:0] input_709;
    input [56:0] input_710;
    input [56:0] input_711;
    input [56:0] input_712;
    input [56:0] input_713;
    input [56:0] input_714;
    input [56:0] input_715;
    input [56:0] input_716;
    input [56:0] input_717;
    input [56:0] input_718;
    input [56:0] input_719;
    input [56:0] input_720;
    input [56:0] input_721;
    input [56:0] input_722;
    input [56:0] input_723;
    input [56:0] input_724;
    input [56:0] input_725;
    input [56:0] input_726;
    input [56:0] input_727;
    input [56:0] input_728;
    input [56:0] input_729;
    input [56:0] input_730;
    input [56:0] input_731;
    input [56:0] input_732;
    input [56:0] input_733;
    input [56:0] input_734;
    input [56:0] input_735;
    input [56:0] input_736;
    input [56:0] input_737;
    input [56:0] input_738;
    input [56:0] input_739;
    input [56:0] input_740;
    input [56:0] input_741;
    input [56:0] input_742;
    input [56:0] input_743;
    input [56:0] input_744;
    input [56:0] input_745;
    input [56:0] input_746;
    input [56:0] input_747;
    input [56:0] input_748;
    input [56:0] input_749;
    input [56:0] input_750;
    input [56:0] input_751;
    input [56:0] input_752;
    input [56:0] input_753;
    input [56:0] input_754;
    input [56:0] input_755;
    input [56:0] input_756;
    input [56:0] input_757;
    input [56:0] input_758;
    input [56:0] input_759;
    input [56:0] input_760;
    input [56:0] input_761;
    input [56:0] input_762;
    input [56:0] input_763;
    input [56:0] input_764;
    input [56:0] input_765;
    input [56:0] input_766;
    input [56:0] input_767;
    input [56:0] input_768;
    input [56:0] input_769;
    input [56:0] input_770;
    input [56:0] input_771;
    input [56:0] input_772;
    input [56:0] input_773;
    input [56:0] input_774;
    input [56:0] input_775;
    input [56:0] input_776;
    input [56:0] input_777;
    input [56:0] input_778;
    input [56:0] input_779;
    input [56:0] input_780;
    input [56:0] input_781;
    input [56:0] input_782;
    input [56:0] input_783;
    input [56:0] input_784;
    input [56:0] input_785;
    input [56:0] input_786;
    input [56:0] input_787;
    input [56:0] input_788;
    input [56:0] input_789;
    input [56:0] input_790;
    input [56:0] input_791;
    input [56:0] input_792;
    input [56:0] input_793;
    input [56:0] input_794;
    input [56:0] input_795;
    input [56:0] input_796;
    input [56:0] input_797;
    input [56:0] input_798;
    input [56:0] input_799;
    input [56:0] input_800;
    input [56:0] input_801;
    input [56:0] input_802;
    input [56:0] input_803;
    input [56:0] input_804;
    input [56:0] input_805;
    input [56:0] input_806;
    input [56:0] input_807;
    input [56:0] input_808;
    input [56:0] input_809;
    input [56:0] input_810;
    input [56:0] input_811;
    input [56:0] input_812;
    input [56:0] input_813;
    input [56:0] input_814;
    input [56:0] input_815;
    input [56:0] input_816;
    input [56:0] input_817;
    input [56:0] input_818;
    input [56:0] input_819;
    input [56:0] input_820;
    input [56:0] input_821;
    input [56:0] input_822;
    input [56:0] input_823;
    input [56:0] input_824;
    input [56:0] input_825;
    input [56:0] input_826;
    input [56:0] input_827;
    input [56:0] input_828;
    input [56:0] input_829;
    input [56:0] input_830;
    input [56:0] input_831;
    input [56:0] input_832;
    input [56:0] input_833;
    input [56:0] input_834;
    input [56:0] input_835;
    input [56:0] input_836;
    input [56:0] input_837;
    input [56:0] input_838;
    input [56:0] input_839;
    input [56:0] input_840;
    input [56:0] input_841;
    input [56:0] input_842;
    input [56:0] input_843;
    input [56:0] input_844;
    input [56:0] input_845;
    input [56:0] input_846;
    input [56:0] input_847;
    input [56:0] input_848;
    input [56:0] input_849;
    input [56:0] input_850;
    input [56:0] input_851;
    input [56:0] input_852;
    input [56:0] input_853;
    input [56:0] input_854;
    input [56:0] input_855;
    input [56:0] input_856;
    input [56:0] input_857;
    input [56:0] input_858;
    input [56:0] input_859;
    input [56:0] input_860;
    input [56:0] input_861;
    input [56:0] input_862;
    input [56:0] input_863;
    input [56:0] input_864;
    input [56:0] input_865;
    input [56:0] input_866;
    input [56:0] input_867;
    input [56:0] input_868;
    input [56:0] input_869;
    input [56:0] input_870;
    input [56:0] input_871;
    input [56:0] input_872;
    input [56:0] input_873;
    input [56:0] input_874;
    input [56:0] input_875;
    input [56:0] input_876;
    input [56:0] input_877;
    input [56:0] input_878;
    input [56:0] input_879;
    input [56:0] input_880;
    input [56:0] input_881;
    input [56:0] input_882;
    input [56:0] input_883;
    input [56:0] input_884;
    input [56:0] input_885;
    input [56:0] input_886;
    input [56:0] input_887;
    input [56:0] input_888;
    input [56:0] input_889;
    input [56:0] input_890;
    input [56:0] input_891;
    input [56:0] input_892;
    input [56:0] input_893;
    input [56:0] input_894;
    input [56:0] input_895;
    input [56:0] input_896;
    input [56:0] input_897;
    input [56:0] input_898;
    input [56:0] input_899;
    input [56:0] input_900;
    input [56:0] input_901;
    input [56:0] input_902;
    input [56:0] input_903;
    input [56:0] input_904;
    input [56:0] input_905;
    input [56:0] input_906;
    input [56:0] input_907;
    input [56:0] input_908;
    input [56:0] input_909;
    input [56:0] input_910;
    input [56:0] input_911;
    input [56:0] input_912;
    input [56:0] input_913;
    input [56:0] input_914;
    input [56:0] input_915;
    input [56:0] input_916;
    input [56:0] input_917;
    input [56:0] input_918;
    input [56:0] input_919;
    input [56:0] input_920;
    input [56:0] input_921;
    input [56:0] input_922;
    input [56:0] input_923;
    input [56:0] input_924;
    input [56:0] input_925;
    input [56:0] input_926;
    input [56:0] input_927;
    input [56:0] input_928;
    input [56:0] input_929;
    input [56:0] input_930;
    input [56:0] input_931;
    input [56:0] input_932;
    input [56:0] input_933;
    input [56:0] input_934;
    input [56:0] input_935;
    input [56:0] input_936;
    input [56:0] input_937;
    input [56:0] input_938;
    input [56:0] input_939;
    input [56:0] input_940;
    input [56:0] input_941;
    input [56:0] input_942;
    input [56:0] input_943;
    input [56:0] input_944;
    input [56:0] input_945;
    input [56:0] input_946;
    input [56:0] input_947;
    input [56:0] input_948;
    input [56:0] input_949;
    input [56:0] input_950;
    input [56:0] input_951;
    input [56:0] input_952;
    input [56:0] input_953;
    input [56:0] input_954;
    input [56:0] input_955;
    input [56:0] input_956;
    input [56:0] input_957;
    input [56:0] input_958;
    input [56:0] input_959;
    input [56:0] input_960;
    input [56:0] input_961;
    input [56:0] input_962;
    input [56:0] input_963;
    input [56:0] input_964;
    input [56:0] input_965;
    input [56:0] input_966;
    input [56:0] input_967;
    input [56:0] input_968;
    input [56:0] input_969;
    input [56:0] input_970;
    input [56:0] input_971;
    input [56:0] input_972;
    input [56:0] input_973;
    input [56:0] input_974;
    input [56:0] input_975;
    input [56:0] input_976;
    input [56:0] input_977;
    input [56:0] input_978;
    input [56:0] input_979;
    input [56:0] input_980;
    input [56:0] input_981;
    input [56:0] input_982;
    input [56:0] input_983;
    input [56:0] input_984;
    input [56:0] input_985;
    input [56:0] input_986;
    input [56:0] input_987;
    input [56:0] input_988;
    input [56:0] input_989;
    input [56:0] input_990;
    input [56:0] input_991;
    input [56:0] input_992;
    input [56:0] input_993;
    input [56:0] input_994;
    input [56:0] input_995;
    input [56:0] input_996;
    input [56:0] input_997;
    input [56:0] input_998;
    input [56:0] input_999;
    input [56:0] input_1000;
    input [56:0] input_1001;
    input [56:0] input_1002;
    input [56:0] input_1003;
    input [56:0] input_1004;
    input [56:0] input_1005;
    input [56:0] input_1006;
    input [56:0] input_1007;
    input [56:0] input_1008;
    input [56:0] input_1009;
    input [56:0] input_1010;
    input [56:0] input_1011;
    input [56:0] input_1012;
    input [56:0] input_1013;
    input [56:0] input_1014;
    input [56:0] input_1015;
    input [56:0] input_1016;
    input [56:0] input_1017;
    input [56:0] input_1018;
    input [56:0] input_1019;
    input [56:0] input_1020;
    input [56:0] input_1021;
    input [56:0] input_1022;
    input [56:0] input_1023;
    input [9:0] sel;
    reg [56:0] result;
  begin
    case (sel)
      10'b0000000000 : begin
        result = input_0;
      end
      10'b0000000001 : begin
        result = input_1;
      end
      10'b0000000010 : begin
        result = input_2;
      end
      10'b0000000011 : begin
        result = input_3;
      end
      10'b0000000100 : begin
        result = input_4;
      end
      10'b0000000101 : begin
        result = input_5;
      end
      10'b0000000110 : begin
        result = input_6;
      end
      10'b0000000111 : begin
        result = input_7;
      end
      10'b0000001000 : begin
        result = input_8;
      end
      10'b0000001001 : begin
        result = input_9;
      end
      10'b0000001010 : begin
        result = input_10;
      end
      10'b0000001011 : begin
        result = input_11;
      end
      10'b0000001100 : begin
        result = input_12;
      end
      10'b0000001101 : begin
        result = input_13;
      end
      10'b0000001110 : begin
        result = input_14;
      end
      10'b0000001111 : begin
        result = input_15;
      end
      10'b0000010000 : begin
        result = input_16;
      end
      10'b0000010001 : begin
        result = input_17;
      end
      10'b0000010010 : begin
        result = input_18;
      end
      10'b0000010011 : begin
        result = input_19;
      end
      10'b0000010100 : begin
        result = input_20;
      end
      10'b0000010101 : begin
        result = input_21;
      end
      10'b0000010110 : begin
        result = input_22;
      end
      10'b0000010111 : begin
        result = input_23;
      end
      10'b0000011000 : begin
        result = input_24;
      end
      10'b0000011001 : begin
        result = input_25;
      end
      10'b0000011010 : begin
        result = input_26;
      end
      10'b0000011011 : begin
        result = input_27;
      end
      10'b0000011100 : begin
        result = input_28;
      end
      10'b0000011101 : begin
        result = input_29;
      end
      10'b0000011110 : begin
        result = input_30;
      end
      10'b0000011111 : begin
        result = input_31;
      end
      10'b0000100000 : begin
        result = input_32;
      end
      10'b0000100001 : begin
        result = input_33;
      end
      10'b0000100010 : begin
        result = input_34;
      end
      10'b0000100011 : begin
        result = input_35;
      end
      10'b0000100100 : begin
        result = input_36;
      end
      10'b0000100101 : begin
        result = input_37;
      end
      10'b0000100110 : begin
        result = input_38;
      end
      10'b0000100111 : begin
        result = input_39;
      end
      10'b0000101000 : begin
        result = input_40;
      end
      10'b0000101001 : begin
        result = input_41;
      end
      10'b0000101010 : begin
        result = input_42;
      end
      10'b0000101011 : begin
        result = input_43;
      end
      10'b0000101100 : begin
        result = input_44;
      end
      10'b0000101101 : begin
        result = input_45;
      end
      10'b0000101110 : begin
        result = input_46;
      end
      10'b0000101111 : begin
        result = input_47;
      end
      10'b0000110000 : begin
        result = input_48;
      end
      10'b0000110001 : begin
        result = input_49;
      end
      10'b0000110010 : begin
        result = input_50;
      end
      10'b0000110011 : begin
        result = input_51;
      end
      10'b0000110100 : begin
        result = input_52;
      end
      10'b0000110101 : begin
        result = input_53;
      end
      10'b0000110110 : begin
        result = input_54;
      end
      10'b0000110111 : begin
        result = input_55;
      end
      10'b0000111000 : begin
        result = input_56;
      end
      10'b0000111001 : begin
        result = input_57;
      end
      10'b0000111010 : begin
        result = input_58;
      end
      10'b0000111011 : begin
        result = input_59;
      end
      10'b0000111100 : begin
        result = input_60;
      end
      10'b0000111101 : begin
        result = input_61;
      end
      10'b0000111110 : begin
        result = input_62;
      end
      10'b0000111111 : begin
        result = input_63;
      end
      10'b0001000000 : begin
        result = input_64;
      end
      10'b0001000001 : begin
        result = input_65;
      end
      10'b0001000010 : begin
        result = input_66;
      end
      10'b0001000011 : begin
        result = input_67;
      end
      10'b0001000100 : begin
        result = input_68;
      end
      10'b0001000101 : begin
        result = input_69;
      end
      10'b0001000110 : begin
        result = input_70;
      end
      10'b0001000111 : begin
        result = input_71;
      end
      10'b0001001000 : begin
        result = input_72;
      end
      10'b0001001001 : begin
        result = input_73;
      end
      10'b0001001010 : begin
        result = input_74;
      end
      10'b0001001011 : begin
        result = input_75;
      end
      10'b0001001100 : begin
        result = input_76;
      end
      10'b0001001101 : begin
        result = input_77;
      end
      10'b0001001110 : begin
        result = input_78;
      end
      10'b0001001111 : begin
        result = input_79;
      end
      10'b0001010000 : begin
        result = input_80;
      end
      10'b0001010001 : begin
        result = input_81;
      end
      10'b0001010010 : begin
        result = input_82;
      end
      10'b0001010011 : begin
        result = input_83;
      end
      10'b0001010100 : begin
        result = input_84;
      end
      10'b0001010101 : begin
        result = input_85;
      end
      10'b0001010110 : begin
        result = input_86;
      end
      10'b0001010111 : begin
        result = input_87;
      end
      10'b0001011000 : begin
        result = input_88;
      end
      10'b0001011001 : begin
        result = input_89;
      end
      10'b0001011010 : begin
        result = input_90;
      end
      10'b0001011011 : begin
        result = input_91;
      end
      10'b0001011100 : begin
        result = input_92;
      end
      10'b0001011101 : begin
        result = input_93;
      end
      10'b0001011110 : begin
        result = input_94;
      end
      10'b0001011111 : begin
        result = input_95;
      end
      10'b0001100000 : begin
        result = input_96;
      end
      10'b0001100001 : begin
        result = input_97;
      end
      10'b0001100010 : begin
        result = input_98;
      end
      10'b0001100011 : begin
        result = input_99;
      end
      10'b0001100100 : begin
        result = input_100;
      end
      10'b0001100101 : begin
        result = input_101;
      end
      10'b0001100110 : begin
        result = input_102;
      end
      10'b0001100111 : begin
        result = input_103;
      end
      10'b0001101000 : begin
        result = input_104;
      end
      10'b0001101001 : begin
        result = input_105;
      end
      10'b0001101010 : begin
        result = input_106;
      end
      10'b0001101011 : begin
        result = input_107;
      end
      10'b0001101100 : begin
        result = input_108;
      end
      10'b0001101101 : begin
        result = input_109;
      end
      10'b0001101110 : begin
        result = input_110;
      end
      10'b0001101111 : begin
        result = input_111;
      end
      10'b0001110000 : begin
        result = input_112;
      end
      10'b0001110001 : begin
        result = input_113;
      end
      10'b0001110010 : begin
        result = input_114;
      end
      10'b0001110011 : begin
        result = input_115;
      end
      10'b0001110100 : begin
        result = input_116;
      end
      10'b0001110101 : begin
        result = input_117;
      end
      10'b0001110110 : begin
        result = input_118;
      end
      10'b0001110111 : begin
        result = input_119;
      end
      10'b0001111000 : begin
        result = input_120;
      end
      10'b0001111001 : begin
        result = input_121;
      end
      10'b0001111010 : begin
        result = input_122;
      end
      10'b0001111011 : begin
        result = input_123;
      end
      10'b0001111100 : begin
        result = input_124;
      end
      10'b0001111101 : begin
        result = input_125;
      end
      10'b0001111110 : begin
        result = input_126;
      end
      10'b0001111111 : begin
        result = input_127;
      end
      10'b0010000000 : begin
        result = input_128;
      end
      10'b0010000001 : begin
        result = input_129;
      end
      10'b0010000010 : begin
        result = input_130;
      end
      10'b0010000011 : begin
        result = input_131;
      end
      10'b0010000100 : begin
        result = input_132;
      end
      10'b0010000101 : begin
        result = input_133;
      end
      10'b0010000110 : begin
        result = input_134;
      end
      10'b0010000111 : begin
        result = input_135;
      end
      10'b0010001000 : begin
        result = input_136;
      end
      10'b0010001001 : begin
        result = input_137;
      end
      10'b0010001010 : begin
        result = input_138;
      end
      10'b0010001011 : begin
        result = input_139;
      end
      10'b0010001100 : begin
        result = input_140;
      end
      10'b0010001101 : begin
        result = input_141;
      end
      10'b0010001110 : begin
        result = input_142;
      end
      10'b0010001111 : begin
        result = input_143;
      end
      10'b0010010000 : begin
        result = input_144;
      end
      10'b0010010001 : begin
        result = input_145;
      end
      10'b0010010010 : begin
        result = input_146;
      end
      10'b0010010011 : begin
        result = input_147;
      end
      10'b0010010100 : begin
        result = input_148;
      end
      10'b0010010101 : begin
        result = input_149;
      end
      10'b0010010110 : begin
        result = input_150;
      end
      10'b0010010111 : begin
        result = input_151;
      end
      10'b0010011000 : begin
        result = input_152;
      end
      10'b0010011001 : begin
        result = input_153;
      end
      10'b0010011010 : begin
        result = input_154;
      end
      10'b0010011011 : begin
        result = input_155;
      end
      10'b0010011100 : begin
        result = input_156;
      end
      10'b0010011101 : begin
        result = input_157;
      end
      10'b0010011110 : begin
        result = input_158;
      end
      10'b0010011111 : begin
        result = input_159;
      end
      10'b0010100000 : begin
        result = input_160;
      end
      10'b0010100001 : begin
        result = input_161;
      end
      10'b0010100010 : begin
        result = input_162;
      end
      10'b0010100011 : begin
        result = input_163;
      end
      10'b0010100100 : begin
        result = input_164;
      end
      10'b0010100101 : begin
        result = input_165;
      end
      10'b0010100110 : begin
        result = input_166;
      end
      10'b0010100111 : begin
        result = input_167;
      end
      10'b0010101000 : begin
        result = input_168;
      end
      10'b0010101001 : begin
        result = input_169;
      end
      10'b0010101010 : begin
        result = input_170;
      end
      10'b0010101011 : begin
        result = input_171;
      end
      10'b0010101100 : begin
        result = input_172;
      end
      10'b0010101101 : begin
        result = input_173;
      end
      10'b0010101110 : begin
        result = input_174;
      end
      10'b0010101111 : begin
        result = input_175;
      end
      10'b0010110000 : begin
        result = input_176;
      end
      10'b0010110001 : begin
        result = input_177;
      end
      10'b0010110010 : begin
        result = input_178;
      end
      10'b0010110011 : begin
        result = input_179;
      end
      10'b0010110100 : begin
        result = input_180;
      end
      10'b0010110101 : begin
        result = input_181;
      end
      10'b0010110110 : begin
        result = input_182;
      end
      10'b0010110111 : begin
        result = input_183;
      end
      10'b0010111000 : begin
        result = input_184;
      end
      10'b0010111001 : begin
        result = input_185;
      end
      10'b0010111010 : begin
        result = input_186;
      end
      10'b0010111011 : begin
        result = input_187;
      end
      10'b0010111100 : begin
        result = input_188;
      end
      10'b0010111101 : begin
        result = input_189;
      end
      10'b0010111110 : begin
        result = input_190;
      end
      10'b0010111111 : begin
        result = input_191;
      end
      10'b0011000000 : begin
        result = input_192;
      end
      10'b0011000001 : begin
        result = input_193;
      end
      10'b0011000010 : begin
        result = input_194;
      end
      10'b0011000011 : begin
        result = input_195;
      end
      10'b0011000100 : begin
        result = input_196;
      end
      10'b0011000101 : begin
        result = input_197;
      end
      10'b0011000110 : begin
        result = input_198;
      end
      10'b0011000111 : begin
        result = input_199;
      end
      10'b0011001000 : begin
        result = input_200;
      end
      10'b0011001001 : begin
        result = input_201;
      end
      10'b0011001010 : begin
        result = input_202;
      end
      10'b0011001011 : begin
        result = input_203;
      end
      10'b0011001100 : begin
        result = input_204;
      end
      10'b0011001101 : begin
        result = input_205;
      end
      10'b0011001110 : begin
        result = input_206;
      end
      10'b0011001111 : begin
        result = input_207;
      end
      10'b0011010000 : begin
        result = input_208;
      end
      10'b0011010001 : begin
        result = input_209;
      end
      10'b0011010010 : begin
        result = input_210;
      end
      10'b0011010011 : begin
        result = input_211;
      end
      10'b0011010100 : begin
        result = input_212;
      end
      10'b0011010101 : begin
        result = input_213;
      end
      10'b0011010110 : begin
        result = input_214;
      end
      10'b0011010111 : begin
        result = input_215;
      end
      10'b0011011000 : begin
        result = input_216;
      end
      10'b0011011001 : begin
        result = input_217;
      end
      10'b0011011010 : begin
        result = input_218;
      end
      10'b0011011011 : begin
        result = input_219;
      end
      10'b0011011100 : begin
        result = input_220;
      end
      10'b0011011101 : begin
        result = input_221;
      end
      10'b0011011110 : begin
        result = input_222;
      end
      10'b0011011111 : begin
        result = input_223;
      end
      10'b0011100000 : begin
        result = input_224;
      end
      10'b0011100001 : begin
        result = input_225;
      end
      10'b0011100010 : begin
        result = input_226;
      end
      10'b0011100011 : begin
        result = input_227;
      end
      10'b0011100100 : begin
        result = input_228;
      end
      10'b0011100101 : begin
        result = input_229;
      end
      10'b0011100110 : begin
        result = input_230;
      end
      10'b0011100111 : begin
        result = input_231;
      end
      10'b0011101000 : begin
        result = input_232;
      end
      10'b0011101001 : begin
        result = input_233;
      end
      10'b0011101010 : begin
        result = input_234;
      end
      10'b0011101011 : begin
        result = input_235;
      end
      10'b0011101100 : begin
        result = input_236;
      end
      10'b0011101101 : begin
        result = input_237;
      end
      10'b0011101110 : begin
        result = input_238;
      end
      10'b0011101111 : begin
        result = input_239;
      end
      10'b0011110000 : begin
        result = input_240;
      end
      10'b0011110001 : begin
        result = input_241;
      end
      10'b0011110010 : begin
        result = input_242;
      end
      10'b0011110011 : begin
        result = input_243;
      end
      10'b0011110100 : begin
        result = input_244;
      end
      10'b0011110101 : begin
        result = input_245;
      end
      10'b0011110110 : begin
        result = input_246;
      end
      10'b0011110111 : begin
        result = input_247;
      end
      10'b0011111000 : begin
        result = input_248;
      end
      10'b0011111001 : begin
        result = input_249;
      end
      10'b0011111010 : begin
        result = input_250;
      end
      10'b0011111011 : begin
        result = input_251;
      end
      10'b0011111100 : begin
        result = input_252;
      end
      10'b0011111101 : begin
        result = input_253;
      end
      10'b0011111110 : begin
        result = input_254;
      end
      10'b0011111111 : begin
        result = input_255;
      end
      10'b0100000000 : begin
        result = input_256;
      end
      10'b0100000001 : begin
        result = input_257;
      end
      10'b0100000010 : begin
        result = input_258;
      end
      10'b0100000011 : begin
        result = input_259;
      end
      10'b0100000100 : begin
        result = input_260;
      end
      10'b0100000101 : begin
        result = input_261;
      end
      10'b0100000110 : begin
        result = input_262;
      end
      10'b0100000111 : begin
        result = input_263;
      end
      10'b0100001000 : begin
        result = input_264;
      end
      10'b0100001001 : begin
        result = input_265;
      end
      10'b0100001010 : begin
        result = input_266;
      end
      10'b0100001011 : begin
        result = input_267;
      end
      10'b0100001100 : begin
        result = input_268;
      end
      10'b0100001101 : begin
        result = input_269;
      end
      10'b0100001110 : begin
        result = input_270;
      end
      10'b0100001111 : begin
        result = input_271;
      end
      10'b0100010000 : begin
        result = input_272;
      end
      10'b0100010001 : begin
        result = input_273;
      end
      10'b0100010010 : begin
        result = input_274;
      end
      10'b0100010011 : begin
        result = input_275;
      end
      10'b0100010100 : begin
        result = input_276;
      end
      10'b0100010101 : begin
        result = input_277;
      end
      10'b0100010110 : begin
        result = input_278;
      end
      10'b0100010111 : begin
        result = input_279;
      end
      10'b0100011000 : begin
        result = input_280;
      end
      10'b0100011001 : begin
        result = input_281;
      end
      10'b0100011010 : begin
        result = input_282;
      end
      10'b0100011011 : begin
        result = input_283;
      end
      10'b0100011100 : begin
        result = input_284;
      end
      10'b0100011101 : begin
        result = input_285;
      end
      10'b0100011110 : begin
        result = input_286;
      end
      10'b0100011111 : begin
        result = input_287;
      end
      10'b0100100000 : begin
        result = input_288;
      end
      10'b0100100001 : begin
        result = input_289;
      end
      10'b0100100010 : begin
        result = input_290;
      end
      10'b0100100011 : begin
        result = input_291;
      end
      10'b0100100100 : begin
        result = input_292;
      end
      10'b0100100101 : begin
        result = input_293;
      end
      10'b0100100110 : begin
        result = input_294;
      end
      10'b0100100111 : begin
        result = input_295;
      end
      10'b0100101000 : begin
        result = input_296;
      end
      10'b0100101001 : begin
        result = input_297;
      end
      10'b0100101010 : begin
        result = input_298;
      end
      10'b0100101011 : begin
        result = input_299;
      end
      10'b0100101100 : begin
        result = input_300;
      end
      10'b0100101101 : begin
        result = input_301;
      end
      10'b0100101110 : begin
        result = input_302;
      end
      10'b0100101111 : begin
        result = input_303;
      end
      10'b0100110000 : begin
        result = input_304;
      end
      10'b0100110001 : begin
        result = input_305;
      end
      10'b0100110010 : begin
        result = input_306;
      end
      10'b0100110011 : begin
        result = input_307;
      end
      10'b0100110100 : begin
        result = input_308;
      end
      10'b0100110101 : begin
        result = input_309;
      end
      10'b0100110110 : begin
        result = input_310;
      end
      10'b0100110111 : begin
        result = input_311;
      end
      10'b0100111000 : begin
        result = input_312;
      end
      10'b0100111001 : begin
        result = input_313;
      end
      10'b0100111010 : begin
        result = input_314;
      end
      10'b0100111011 : begin
        result = input_315;
      end
      10'b0100111100 : begin
        result = input_316;
      end
      10'b0100111101 : begin
        result = input_317;
      end
      10'b0100111110 : begin
        result = input_318;
      end
      10'b0100111111 : begin
        result = input_319;
      end
      10'b0101000000 : begin
        result = input_320;
      end
      10'b0101000001 : begin
        result = input_321;
      end
      10'b0101000010 : begin
        result = input_322;
      end
      10'b0101000011 : begin
        result = input_323;
      end
      10'b0101000100 : begin
        result = input_324;
      end
      10'b0101000101 : begin
        result = input_325;
      end
      10'b0101000110 : begin
        result = input_326;
      end
      10'b0101000111 : begin
        result = input_327;
      end
      10'b0101001000 : begin
        result = input_328;
      end
      10'b0101001001 : begin
        result = input_329;
      end
      10'b0101001010 : begin
        result = input_330;
      end
      10'b0101001011 : begin
        result = input_331;
      end
      10'b0101001100 : begin
        result = input_332;
      end
      10'b0101001101 : begin
        result = input_333;
      end
      10'b0101001110 : begin
        result = input_334;
      end
      10'b0101001111 : begin
        result = input_335;
      end
      10'b0101010000 : begin
        result = input_336;
      end
      10'b0101010001 : begin
        result = input_337;
      end
      10'b0101010010 : begin
        result = input_338;
      end
      10'b0101010011 : begin
        result = input_339;
      end
      10'b0101010100 : begin
        result = input_340;
      end
      10'b0101010101 : begin
        result = input_341;
      end
      10'b0101010110 : begin
        result = input_342;
      end
      10'b0101010111 : begin
        result = input_343;
      end
      10'b0101011000 : begin
        result = input_344;
      end
      10'b0101011001 : begin
        result = input_345;
      end
      10'b0101011010 : begin
        result = input_346;
      end
      10'b0101011011 : begin
        result = input_347;
      end
      10'b0101011100 : begin
        result = input_348;
      end
      10'b0101011101 : begin
        result = input_349;
      end
      10'b0101011110 : begin
        result = input_350;
      end
      10'b0101011111 : begin
        result = input_351;
      end
      10'b0101100000 : begin
        result = input_352;
      end
      10'b0101100001 : begin
        result = input_353;
      end
      10'b0101100010 : begin
        result = input_354;
      end
      10'b0101100011 : begin
        result = input_355;
      end
      10'b0101100100 : begin
        result = input_356;
      end
      10'b0101100101 : begin
        result = input_357;
      end
      10'b0101100110 : begin
        result = input_358;
      end
      10'b0101100111 : begin
        result = input_359;
      end
      10'b0101101000 : begin
        result = input_360;
      end
      10'b0101101001 : begin
        result = input_361;
      end
      10'b0101101010 : begin
        result = input_362;
      end
      10'b0101101011 : begin
        result = input_363;
      end
      10'b0101101100 : begin
        result = input_364;
      end
      10'b0101101101 : begin
        result = input_365;
      end
      10'b0101101110 : begin
        result = input_366;
      end
      10'b0101101111 : begin
        result = input_367;
      end
      10'b0101110000 : begin
        result = input_368;
      end
      10'b0101110001 : begin
        result = input_369;
      end
      10'b0101110010 : begin
        result = input_370;
      end
      10'b0101110011 : begin
        result = input_371;
      end
      10'b0101110100 : begin
        result = input_372;
      end
      10'b0101110101 : begin
        result = input_373;
      end
      10'b0101110110 : begin
        result = input_374;
      end
      10'b0101110111 : begin
        result = input_375;
      end
      10'b0101111000 : begin
        result = input_376;
      end
      10'b0101111001 : begin
        result = input_377;
      end
      10'b0101111010 : begin
        result = input_378;
      end
      10'b0101111011 : begin
        result = input_379;
      end
      10'b0101111100 : begin
        result = input_380;
      end
      10'b0101111101 : begin
        result = input_381;
      end
      10'b0101111110 : begin
        result = input_382;
      end
      10'b0101111111 : begin
        result = input_383;
      end
      10'b0110000000 : begin
        result = input_384;
      end
      10'b0110000001 : begin
        result = input_385;
      end
      10'b0110000010 : begin
        result = input_386;
      end
      10'b0110000011 : begin
        result = input_387;
      end
      10'b0110000100 : begin
        result = input_388;
      end
      10'b0110000101 : begin
        result = input_389;
      end
      10'b0110000110 : begin
        result = input_390;
      end
      10'b0110000111 : begin
        result = input_391;
      end
      10'b0110001000 : begin
        result = input_392;
      end
      10'b0110001001 : begin
        result = input_393;
      end
      10'b0110001010 : begin
        result = input_394;
      end
      10'b0110001011 : begin
        result = input_395;
      end
      10'b0110001100 : begin
        result = input_396;
      end
      10'b0110001101 : begin
        result = input_397;
      end
      10'b0110001110 : begin
        result = input_398;
      end
      10'b0110001111 : begin
        result = input_399;
      end
      10'b0110010000 : begin
        result = input_400;
      end
      10'b0110010001 : begin
        result = input_401;
      end
      10'b0110010010 : begin
        result = input_402;
      end
      10'b0110010011 : begin
        result = input_403;
      end
      10'b0110010100 : begin
        result = input_404;
      end
      10'b0110010101 : begin
        result = input_405;
      end
      10'b0110010110 : begin
        result = input_406;
      end
      10'b0110010111 : begin
        result = input_407;
      end
      10'b0110011000 : begin
        result = input_408;
      end
      10'b0110011001 : begin
        result = input_409;
      end
      10'b0110011010 : begin
        result = input_410;
      end
      10'b0110011011 : begin
        result = input_411;
      end
      10'b0110011100 : begin
        result = input_412;
      end
      10'b0110011101 : begin
        result = input_413;
      end
      10'b0110011110 : begin
        result = input_414;
      end
      10'b0110011111 : begin
        result = input_415;
      end
      10'b0110100000 : begin
        result = input_416;
      end
      10'b0110100001 : begin
        result = input_417;
      end
      10'b0110100010 : begin
        result = input_418;
      end
      10'b0110100011 : begin
        result = input_419;
      end
      10'b0110100100 : begin
        result = input_420;
      end
      10'b0110100101 : begin
        result = input_421;
      end
      10'b0110100110 : begin
        result = input_422;
      end
      10'b0110100111 : begin
        result = input_423;
      end
      10'b0110101000 : begin
        result = input_424;
      end
      10'b0110101001 : begin
        result = input_425;
      end
      10'b0110101010 : begin
        result = input_426;
      end
      10'b0110101011 : begin
        result = input_427;
      end
      10'b0110101100 : begin
        result = input_428;
      end
      10'b0110101101 : begin
        result = input_429;
      end
      10'b0110101110 : begin
        result = input_430;
      end
      10'b0110101111 : begin
        result = input_431;
      end
      10'b0110110000 : begin
        result = input_432;
      end
      10'b0110110001 : begin
        result = input_433;
      end
      10'b0110110010 : begin
        result = input_434;
      end
      10'b0110110011 : begin
        result = input_435;
      end
      10'b0110110100 : begin
        result = input_436;
      end
      10'b0110110101 : begin
        result = input_437;
      end
      10'b0110110110 : begin
        result = input_438;
      end
      10'b0110110111 : begin
        result = input_439;
      end
      10'b0110111000 : begin
        result = input_440;
      end
      10'b0110111001 : begin
        result = input_441;
      end
      10'b0110111010 : begin
        result = input_442;
      end
      10'b0110111011 : begin
        result = input_443;
      end
      10'b0110111100 : begin
        result = input_444;
      end
      10'b0110111101 : begin
        result = input_445;
      end
      10'b0110111110 : begin
        result = input_446;
      end
      10'b0110111111 : begin
        result = input_447;
      end
      10'b0111000000 : begin
        result = input_448;
      end
      10'b0111000001 : begin
        result = input_449;
      end
      10'b0111000010 : begin
        result = input_450;
      end
      10'b0111000011 : begin
        result = input_451;
      end
      10'b0111000100 : begin
        result = input_452;
      end
      10'b0111000101 : begin
        result = input_453;
      end
      10'b0111000110 : begin
        result = input_454;
      end
      10'b0111000111 : begin
        result = input_455;
      end
      10'b0111001000 : begin
        result = input_456;
      end
      10'b0111001001 : begin
        result = input_457;
      end
      10'b0111001010 : begin
        result = input_458;
      end
      10'b0111001011 : begin
        result = input_459;
      end
      10'b0111001100 : begin
        result = input_460;
      end
      10'b0111001101 : begin
        result = input_461;
      end
      10'b0111001110 : begin
        result = input_462;
      end
      10'b0111001111 : begin
        result = input_463;
      end
      10'b0111010000 : begin
        result = input_464;
      end
      10'b0111010001 : begin
        result = input_465;
      end
      10'b0111010010 : begin
        result = input_466;
      end
      10'b0111010011 : begin
        result = input_467;
      end
      10'b0111010100 : begin
        result = input_468;
      end
      10'b0111010101 : begin
        result = input_469;
      end
      10'b0111010110 : begin
        result = input_470;
      end
      10'b0111010111 : begin
        result = input_471;
      end
      10'b0111011000 : begin
        result = input_472;
      end
      10'b0111011001 : begin
        result = input_473;
      end
      10'b0111011010 : begin
        result = input_474;
      end
      10'b0111011011 : begin
        result = input_475;
      end
      10'b0111011100 : begin
        result = input_476;
      end
      10'b0111011101 : begin
        result = input_477;
      end
      10'b0111011110 : begin
        result = input_478;
      end
      10'b0111011111 : begin
        result = input_479;
      end
      10'b0111100000 : begin
        result = input_480;
      end
      10'b0111100001 : begin
        result = input_481;
      end
      10'b0111100010 : begin
        result = input_482;
      end
      10'b0111100011 : begin
        result = input_483;
      end
      10'b0111100100 : begin
        result = input_484;
      end
      10'b0111100101 : begin
        result = input_485;
      end
      10'b0111100110 : begin
        result = input_486;
      end
      10'b0111100111 : begin
        result = input_487;
      end
      10'b0111101000 : begin
        result = input_488;
      end
      10'b0111101001 : begin
        result = input_489;
      end
      10'b0111101010 : begin
        result = input_490;
      end
      10'b0111101011 : begin
        result = input_491;
      end
      10'b0111101100 : begin
        result = input_492;
      end
      10'b0111101101 : begin
        result = input_493;
      end
      10'b0111101110 : begin
        result = input_494;
      end
      10'b0111101111 : begin
        result = input_495;
      end
      10'b0111110000 : begin
        result = input_496;
      end
      10'b0111110001 : begin
        result = input_497;
      end
      10'b0111110010 : begin
        result = input_498;
      end
      10'b0111110011 : begin
        result = input_499;
      end
      10'b0111110100 : begin
        result = input_500;
      end
      10'b0111110101 : begin
        result = input_501;
      end
      10'b0111110110 : begin
        result = input_502;
      end
      10'b0111110111 : begin
        result = input_503;
      end
      10'b0111111000 : begin
        result = input_504;
      end
      10'b0111111001 : begin
        result = input_505;
      end
      10'b0111111010 : begin
        result = input_506;
      end
      10'b0111111011 : begin
        result = input_507;
      end
      10'b0111111100 : begin
        result = input_508;
      end
      10'b0111111101 : begin
        result = input_509;
      end
      10'b0111111110 : begin
        result = input_510;
      end
      10'b0111111111 : begin
        result = input_511;
      end
      10'b1000000000 : begin
        result = input_512;
      end
      10'b1000000001 : begin
        result = input_513;
      end
      10'b1000000010 : begin
        result = input_514;
      end
      10'b1000000011 : begin
        result = input_515;
      end
      10'b1000000100 : begin
        result = input_516;
      end
      10'b1000000101 : begin
        result = input_517;
      end
      10'b1000000110 : begin
        result = input_518;
      end
      10'b1000000111 : begin
        result = input_519;
      end
      10'b1000001000 : begin
        result = input_520;
      end
      10'b1000001001 : begin
        result = input_521;
      end
      10'b1000001010 : begin
        result = input_522;
      end
      10'b1000001011 : begin
        result = input_523;
      end
      10'b1000001100 : begin
        result = input_524;
      end
      10'b1000001101 : begin
        result = input_525;
      end
      10'b1000001110 : begin
        result = input_526;
      end
      10'b1000001111 : begin
        result = input_527;
      end
      10'b1000010000 : begin
        result = input_528;
      end
      10'b1000010001 : begin
        result = input_529;
      end
      10'b1000010010 : begin
        result = input_530;
      end
      10'b1000010011 : begin
        result = input_531;
      end
      10'b1000010100 : begin
        result = input_532;
      end
      10'b1000010101 : begin
        result = input_533;
      end
      10'b1000010110 : begin
        result = input_534;
      end
      10'b1000010111 : begin
        result = input_535;
      end
      10'b1000011000 : begin
        result = input_536;
      end
      10'b1000011001 : begin
        result = input_537;
      end
      10'b1000011010 : begin
        result = input_538;
      end
      10'b1000011011 : begin
        result = input_539;
      end
      10'b1000011100 : begin
        result = input_540;
      end
      10'b1000011101 : begin
        result = input_541;
      end
      10'b1000011110 : begin
        result = input_542;
      end
      10'b1000011111 : begin
        result = input_543;
      end
      10'b1000100000 : begin
        result = input_544;
      end
      10'b1000100001 : begin
        result = input_545;
      end
      10'b1000100010 : begin
        result = input_546;
      end
      10'b1000100011 : begin
        result = input_547;
      end
      10'b1000100100 : begin
        result = input_548;
      end
      10'b1000100101 : begin
        result = input_549;
      end
      10'b1000100110 : begin
        result = input_550;
      end
      10'b1000100111 : begin
        result = input_551;
      end
      10'b1000101000 : begin
        result = input_552;
      end
      10'b1000101001 : begin
        result = input_553;
      end
      10'b1000101010 : begin
        result = input_554;
      end
      10'b1000101011 : begin
        result = input_555;
      end
      10'b1000101100 : begin
        result = input_556;
      end
      10'b1000101101 : begin
        result = input_557;
      end
      10'b1000101110 : begin
        result = input_558;
      end
      10'b1000101111 : begin
        result = input_559;
      end
      10'b1000110000 : begin
        result = input_560;
      end
      10'b1000110001 : begin
        result = input_561;
      end
      10'b1000110010 : begin
        result = input_562;
      end
      10'b1000110011 : begin
        result = input_563;
      end
      10'b1000110100 : begin
        result = input_564;
      end
      10'b1000110101 : begin
        result = input_565;
      end
      10'b1000110110 : begin
        result = input_566;
      end
      10'b1000110111 : begin
        result = input_567;
      end
      10'b1000111000 : begin
        result = input_568;
      end
      10'b1000111001 : begin
        result = input_569;
      end
      10'b1000111010 : begin
        result = input_570;
      end
      10'b1000111011 : begin
        result = input_571;
      end
      10'b1000111100 : begin
        result = input_572;
      end
      10'b1000111101 : begin
        result = input_573;
      end
      10'b1000111110 : begin
        result = input_574;
      end
      10'b1000111111 : begin
        result = input_575;
      end
      10'b1001000000 : begin
        result = input_576;
      end
      10'b1001000001 : begin
        result = input_577;
      end
      10'b1001000010 : begin
        result = input_578;
      end
      10'b1001000011 : begin
        result = input_579;
      end
      10'b1001000100 : begin
        result = input_580;
      end
      10'b1001000101 : begin
        result = input_581;
      end
      10'b1001000110 : begin
        result = input_582;
      end
      10'b1001000111 : begin
        result = input_583;
      end
      10'b1001001000 : begin
        result = input_584;
      end
      10'b1001001001 : begin
        result = input_585;
      end
      10'b1001001010 : begin
        result = input_586;
      end
      10'b1001001011 : begin
        result = input_587;
      end
      10'b1001001100 : begin
        result = input_588;
      end
      10'b1001001101 : begin
        result = input_589;
      end
      10'b1001001110 : begin
        result = input_590;
      end
      10'b1001001111 : begin
        result = input_591;
      end
      10'b1001010000 : begin
        result = input_592;
      end
      10'b1001010001 : begin
        result = input_593;
      end
      10'b1001010010 : begin
        result = input_594;
      end
      10'b1001010011 : begin
        result = input_595;
      end
      10'b1001010100 : begin
        result = input_596;
      end
      10'b1001010101 : begin
        result = input_597;
      end
      10'b1001010110 : begin
        result = input_598;
      end
      10'b1001010111 : begin
        result = input_599;
      end
      10'b1001011000 : begin
        result = input_600;
      end
      10'b1001011001 : begin
        result = input_601;
      end
      10'b1001011010 : begin
        result = input_602;
      end
      10'b1001011011 : begin
        result = input_603;
      end
      10'b1001011100 : begin
        result = input_604;
      end
      10'b1001011101 : begin
        result = input_605;
      end
      10'b1001011110 : begin
        result = input_606;
      end
      10'b1001011111 : begin
        result = input_607;
      end
      10'b1001100000 : begin
        result = input_608;
      end
      10'b1001100001 : begin
        result = input_609;
      end
      10'b1001100010 : begin
        result = input_610;
      end
      10'b1001100011 : begin
        result = input_611;
      end
      10'b1001100100 : begin
        result = input_612;
      end
      10'b1001100101 : begin
        result = input_613;
      end
      10'b1001100110 : begin
        result = input_614;
      end
      10'b1001100111 : begin
        result = input_615;
      end
      10'b1001101000 : begin
        result = input_616;
      end
      10'b1001101001 : begin
        result = input_617;
      end
      10'b1001101010 : begin
        result = input_618;
      end
      10'b1001101011 : begin
        result = input_619;
      end
      10'b1001101100 : begin
        result = input_620;
      end
      10'b1001101101 : begin
        result = input_621;
      end
      10'b1001101110 : begin
        result = input_622;
      end
      10'b1001101111 : begin
        result = input_623;
      end
      10'b1001110000 : begin
        result = input_624;
      end
      10'b1001110001 : begin
        result = input_625;
      end
      10'b1001110010 : begin
        result = input_626;
      end
      10'b1001110011 : begin
        result = input_627;
      end
      10'b1001110100 : begin
        result = input_628;
      end
      10'b1001110101 : begin
        result = input_629;
      end
      10'b1001110110 : begin
        result = input_630;
      end
      10'b1001110111 : begin
        result = input_631;
      end
      10'b1001111000 : begin
        result = input_632;
      end
      10'b1001111001 : begin
        result = input_633;
      end
      10'b1001111010 : begin
        result = input_634;
      end
      10'b1001111011 : begin
        result = input_635;
      end
      10'b1001111100 : begin
        result = input_636;
      end
      10'b1001111101 : begin
        result = input_637;
      end
      10'b1001111110 : begin
        result = input_638;
      end
      10'b1001111111 : begin
        result = input_639;
      end
      10'b1010000000 : begin
        result = input_640;
      end
      10'b1010000001 : begin
        result = input_641;
      end
      10'b1010000010 : begin
        result = input_642;
      end
      10'b1010000011 : begin
        result = input_643;
      end
      10'b1010000100 : begin
        result = input_644;
      end
      10'b1010000101 : begin
        result = input_645;
      end
      10'b1010000110 : begin
        result = input_646;
      end
      10'b1010000111 : begin
        result = input_647;
      end
      10'b1010001000 : begin
        result = input_648;
      end
      10'b1010001001 : begin
        result = input_649;
      end
      10'b1010001010 : begin
        result = input_650;
      end
      10'b1010001011 : begin
        result = input_651;
      end
      10'b1010001100 : begin
        result = input_652;
      end
      10'b1010001101 : begin
        result = input_653;
      end
      10'b1010001110 : begin
        result = input_654;
      end
      10'b1010001111 : begin
        result = input_655;
      end
      10'b1010010000 : begin
        result = input_656;
      end
      10'b1010010001 : begin
        result = input_657;
      end
      10'b1010010010 : begin
        result = input_658;
      end
      10'b1010010011 : begin
        result = input_659;
      end
      10'b1010010100 : begin
        result = input_660;
      end
      10'b1010010101 : begin
        result = input_661;
      end
      10'b1010010110 : begin
        result = input_662;
      end
      10'b1010010111 : begin
        result = input_663;
      end
      10'b1010011000 : begin
        result = input_664;
      end
      10'b1010011001 : begin
        result = input_665;
      end
      10'b1010011010 : begin
        result = input_666;
      end
      10'b1010011011 : begin
        result = input_667;
      end
      10'b1010011100 : begin
        result = input_668;
      end
      10'b1010011101 : begin
        result = input_669;
      end
      10'b1010011110 : begin
        result = input_670;
      end
      10'b1010011111 : begin
        result = input_671;
      end
      10'b1010100000 : begin
        result = input_672;
      end
      10'b1010100001 : begin
        result = input_673;
      end
      10'b1010100010 : begin
        result = input_674;
      end
      10'b1010100011 : begin
        result = input_675;
      end
      10'b1010100100 : begin
        result = input_676;
      end
      10'b1010100101 : begin
        result = input_677;
      end
      10'b1010100110 : begin
        result = input_678;
      end
      10'b1010100111 : begin
        result = input_679;
      end
      10'b1010101000 : begin
        result = input_680;
      end
      10'b1010101001 : begin
        result = input_681;
      end
      10'b1010101010 : begin
        result = input_682;
      end
      10'b1010101011 : begin
        result = input_683;
      end
      10'b1010101100 : begin
        result = input_684;
      end
      10'b1010101101 : begin
        result = input_685;
      end
      10'b1010101110 : begin
        result = input_686;
      end
      10'b1010101111 : begin
        result = input_687;
      end
      10'b1010110000 : begin
        result = input_688;
      end
      10'b1010110001 : begin
        result = input_689;
      end
      10'b1010110010 : begin
        result = input_690;
      end
      10'b1010110011 : begin
        result = input_691;
      end
      10'b1010110100 : begin
        result = input_692;
      end
      10'b1010110101 : begin
        result = input_693;
      end
      10'b1010110110 : begin
        result = input_694;
      end
      10'b1010110111 : begin
        result = input_695;
      end
      10'b1010111000 : begin
        result = input_696;
      end
      10'b1010111001 : begin
        result = input_697;
      end
      10'b1010111010 : begin
        result = input_698;
      end
      10'b1010111011 : begin
        result = input_699;
      end
      10'b1010111100 : begin
        result = input_700;
      end
      10'b1010111101 : begin
        result = input_701;
      end
      10'b1010111110 : begin
        result = input_702;
      end
      10'b1010111111 : begin
        result = input_703;
      end
      10'b1011000000 : begin
        result = input_704;
      end
      10'b1011000001 : begin
        result = input_705;
      end
      10'b1011000010 : begin
        result = input_706;
      end
      10'b1011000011 : begin
        result = input_707;
      end
      10'b1011000100 : begin
        result = input_708;
      end
      10'b1011000101 : begin
        result = input_709;
      end
      10'b1011000110 : begin
        result = input_710;
      end
      10'b1011000111 : begin
        result = input_711;
      end
      10'b1011001000 : begin
        result = input_712;
      end
      10'b1011001001 : begin
        result = input_713;
      end
      10'b1011001010 : begin
        result = input_714;
      end
      10'b1011001011 : begin
        result = input_715;
      end
      10'b1011001100 : begin
        result = input_716;
      end
      10'b1011001101 : begin
        result = input_717;
      end
      10'b1011001110 : begin
        result = input_718;
      end
      10'b1011001111 : begin
        result = input_719;
      end
      10'b1011010000 : begin
        result = input_720;
      end
      10'b1011010001 : begin
        result = input_721;
      end
      10'b1011010010 : begin
        result = input_722;
      end
      10'b1011010011 : begin
        result = input_723;
      end
      10'b1011010100 : begin
        result = input_724;
      end
      10'b1011010101 : begin
        result = input_725;
      end
      10'b1011010110 : begin
        result = input_726;
      end
      10'b1011010111 : begin
        result = input_727;
      end
      10'b1011011000 : begin
        result = input_728;
      end
      10'b1011011001 : begin
        result = input_729;
      end
      10'b1011011010 : begin
        result = input_730;
      end
      10'b1011011011 : begin
        result = input_731;
      end
      10'b1011011100 : begin
        result = input_732;
      end
      10'b1011011101 : begin
        result = input_733;
      end
      10'b1011011110 : begin
        result = input_734;
      end
      10'b1011011111 : begin
        result = input_735;
      end
      10'b1011100000 : begin
        result = input_736;
      end
      10'b1011100001 : begin
        result = input_737;
      end
      10'b1011100010 : begin
        result = input_738;
      end
      10'b1011100011 : begin
        result = input_739;
      end
      10'b1011100100 : begin
        result = input_740;
      end
      10'b1011100101 : begin
        result = input_741;
      end
      10'b1011100110 : begin
        result = input_742;
      end
      10'b1011100111 : begin
        result = input_743;
      end
      10'b1011101000 : begin
        result = input_744;
      end
      10'b1011101001 : begin
        result = input_745;
      end
      10'b1011101010 : begin
        result = input_746;
      end
      10'b1011101011 : begin
        result = input_747;
      end
      10'b1011101100 : begin
        result = input_748;
      end
      10'b1011101101 : begin
        result = input_749;
      end
      10'b1011101110 : begin
        result = input_750;
      end
      10'b1011101111 : begin
        result = input_751;
      end
      10'b1011110000 : begin
        result = input_752;
      end
      10'b1011110001 : begin
        result = input_753;
      end
      10'b1011110010 : begin
        result = input_754;
      end
      10'b1011110011 : begin
        result = input_755;
      end
      10'b1011110100 : begin
        result = input_756;
      end
      10'b1011110101 : begin
        result = input_757;
      end
      10'b1011110110 : begin
        result = input_758;
      end
      10'b1011110111 : begin
        result = input_759;
      end
      10'b1011111000 : begin
        result = input_760;
      end
      10'b1011111001 : begin
        result = input_761;
      end
      10'b1011111010 : begin
        result = input_762;
      end
      10'b1011111011 : begin
        result = input_763;
      end
      10'b1011111100 : begin
        result = input_764;
      end
      10'b1011111101 : begin
        result = input_765;
      end
      10'b1011111110 : begin
        result = input_766;
      end
      10'b1011111111 : begin
        result = input_767;
      end
      10'b1100000000 : begin
        result = input_768;
      end
      10'b1100000001 : begin
        result = input_769;
      end
      10'b1100000010 : begin
        result = input_770;
      end
      10'b1100000011 : begin
        result = input_771;
      end
      10'b1100000100 : begin
        result = input_772;
      end
      10'b1100000101 : begin
        result = input_773;
      end
      10'b1100000110 : begin
        result = input_774;
      end
      10'b1100000111 : begin
        result = input_775;
      end
      10'b1100001000 : begin
        result = input_776;
      end
      10'b1100001001 : begin
        result = input_777;
      end
      10'b1100001010 : begin
        result = input_778;
      end
      10'b1100001011 : begin
        result = input_779;
      end
      10'b1100001100 : begin
        result = input_780;
      end
      10'b1100001101 : begin
        result = input_781;
      end
      10'b1100001110 : begin
        result = input_782;
      end
      10'b1100001111 : begin
        result = input_783;
      end
      10'b1100010000 : begin
        result = input_784;
      end
      10'b1100010001 : begin
        result = input_785;
      end
      10'b1100010010 : begin
        result = input_786;
      end
      10'b1100010011 : begin
        result = input_787;
      end
      10'b1100010100 : begin
        result = input_788;
      end
      10'b1100010101 : begin
        result = input_789;
      end
      10'b1100010110 : begin
        result = input_790;
      end
      10'b1100010111 : begin
        result = input_791;
      end
      10'b1100011000 : begin
        result = input_792;
      end
      10'b1100011001 : begin
        result = input_793;
      end
      10'b1100011010 : begin
        result = input_794;
      end
      10'b1100011011 : begin
        result = input_795;
      end
      10'b1100011100 : begin
        result = input_796;
      end
      10'b1100011101 : begin
        result = input_797;
      end
      10'b1100011110 : begin
        result = input_798;
      end
      10'b1100011111 : begin
        result = input_799;
      end
      10'b1100100000 : begin
        result = input_800;
      end
      10'b1100100001 : begin
        result = input_801;
      end
      10'b1100100010 : begin
        result = input_802;
      end
      10'b1100100011 : begin
        result = input_803;
      end
      10'b1100100100 : begin
        result = input_804;
      end
      10'b1100100101 : begin
        result = input_805;
      end
      10'b1100100110 : begin
        result = input_806;
      end
      10'b1100100111 : begin
        result = input_807;
      end
      10'b1100101000 : begin
        result = input_808;
      end
      10'b1100101001 : begin
        result = input_809;
      end
      10'b1100101010 : begin
        result = input_810;
      end
      10'b1100101011 : begin
        result = input_811;
      end
      10'b1100101100 : begin
        result = input_812;
      end
      10'b1100101101 : begin
        result = input_813;
      end
      10'b1100101110 : begin
        result = input_814;
      end
      10'b1100101111 : begin
        result = input_815;
      end
      10'b1100110000 : begin
        result = input_816;
      end
      10'b1100110001 : begin
        result = input_817;
      end
      10'b1100110010 : begin
        result = input_818;
      end
      10'b1100110011 : begin
        result = input_819;
      end
      10'b1100110100 : begin
        result = input_820;
      end
      10'b1100110101 : begin
        result = input_821;
      end
      10'b1100110110 : begin
        result = input_822;
      end
      10'b1100110111 : begin
        result = input_823;
      end
      10'b1100111000 : begin
        result = input_824;
      end
      10'b1100111001 : begin
        result = input_825;
      end
      10'b1100111010 : begin
        result = input_826;
      end
      10'b1100111011 : begin
        result = input_827;
      end
      10'b1100111100 : begin
        result = input_828;
      end
      10'b1100111101 : begin
        result = input_829;
      end
      10'b1100111110 : begin
        result = input_830;
      end
      10'b1100111111 : begin
        result = input_831;
      end
      10'b1101000000 : begin
        result = input_832;
      end
      10'b1101000001 : begin
        result = input_833;
      end
      10'b1101000010 : begin
        result = input_834;
      end
      10'b1101000011 : begin
        result = input_835;
      end
      10'b1101000100 : begin
        result = input_836;
      end
      10'b1101000101 : begin
        result = input_837;
      end
      10'b1101000110 : begin
        result = input_838;
      end
      10'b1101000111 : begin
        result = input_839;
      end
      10'b1101001000 : begin
        result = input_840;
      end
      10'b1101001001 : begin
        result = input_841;
      end
      10'b1101001010 : begin
        result = input_842;
      end
      10'b1101001011 : begin
        result = input_843;
      end
      10'b1101001100 : begin
        result = input_844;
      end
      10'b1101001101 : begin
        result = input_845;
      end
      10'b1101001110 : begin
        result = input_846;
      end
      10'b1101001111 : begin
        result = input_847;
      end
      10'b1101010000 : begin
        result = input_848;
      end
      10'b1101010001 : begin
        result = input_849;
      end
      10'b1101010010 : begin
        result = input_850;
      end
      10'b1101010011 : begin
        result = input_851;
      end
      10'b1101010100 : begin
        result = input_852;
      end
      10'b1101010101 : begin
        result = input_853;
      end
      10'b1101010110 : begin
        result = input_854;
      end
      10'b1101010111 : begin
        result = input_855;
      end
      10'b1101011000 : begin
        result = input_856;
      end
      10'b1101011001 : begin
        result = input_857;
      end
      10'b1101011010 : begin
        result = input_858;
      end
      10'b1101011011 : begin
        result = input_859;
      end
      10'b1101011100 : begin
        result = input_860;
      end
      10'b1101011101 : begin
        result = input_861;
      end
      10'b1101011110 : begin
        result = input_862;
      end
      10'b1101011111 : begin
        result = input_863;
      end
      10'b1101100000 : begin
        result = input_864;
      end
      10'b1101100001 : begin
        result = input_865;
      end
      10'b1101100010 : begin
        result = input_866;
      end
      10'b1101100011 : begin
        result = input_867;
      end
      10'b1101100100 : begin
        result = input_868;
      end
      10'b1101100101 : begin
        result = input_869;
      end
      10'b1101100110 : begin
        result = input_870;
      end
      10'b1101100111 : begin
        result = input_871;
      end
      10'b1101101000 : begin
        result = input_872;
      end
      10'b1101101001 : begin
        result = input_873;
      end
      10'b1101101010 : begin
        result = input_874;
      end
      10'b1101101011 : begin
        result = input_875;
      end
      10'b1101101100 : begin
        result = input_876;
      end
      10'b1101101101 : begin
        result = input_877;
      end
      10'b1101101110 : begin
        result = input_878;
      end
      10'b1101101111 : begin
        result = input_879;
      end
      10'b1101110000 : begin
        result = input_880;
      end
      10'b1101110001 : begin
        result = input_881;
      end
      10'b1101110010 : begin
        result = input_882;
      end
      10'b1101110011 : begin
        result = input_883;
      end
      10'b1101110100 : begin
        result = input_884;
      end
      10'b1101110101 : begin
        result = input_885;
      end
      10'b1101110110 : begin
        result = input_886;
      end
      10'b1101110111 : begin
        result = input_887;
      end
      10'b1101111000 : begin
        result = input_888;
      end
      10'b1101111001 : begin
        result = input_889;
      end
      10'b1101111010 : begin
        result = input_890;
      end
      10'b1101111011 : begin
        result = input_891;
      end
      10'b1101111100 : begin
        result = input_892;
      end
      10'b1101111101 : begin
        result = input_893;
      end
      10'b1101111110 : begin
        result = input_894;
      end
      10'b1101111111 : begin
        result = input_895;
      end
      10'b1110000000 : begin
        result = input_896;
      end
      10'b1110000001 : begin
        result = input_897;
      end
      10'b1110000010 : begin
        result = input_898;
      end
      10'b1110000011 : begin
        result = input_899;
      end
      10'b1110000100 : begin
        result = input_900;
      end
      10'b1110000101 : begin
        result = input_901;
      end
      10'b1110000110 : begin
        result = input_902;
      end
      10'b1110000111 : begin
        result = input_903;
      end
      10'b1110001000 : begin
        result = input_904;
      end
      10'b1110001001 : begin
        result = input_905;
      end
      10'b1110001010 : begin
        result = input_906;
      end
      10'b1110001011 : begin
        result = input_907;
      end
      10'b1110001100 : begin
        result = input_908;
      end
      10'b1110001101 : begin
        result = input_909;
      end
      10'b1110001110 : begin
        result = input_910;
      end
      10'b1110001111 : begin
        result = input_911;
      end
      10'b1110010000 : begin
        result = input_912;
      end
      10'b1110010001 : begin
        result = input_913;
      end
      10'b1110010010 : begin
        result = input_914;
      end
      10'b1110010011 : begin
        result = input_915;
      end
      10'b1110010100 : begin
        result = input_916;
      end
      10'b1110010101 : begin
        result = input_917;
      end
      10'b1110010110 : begin
        result = input_918;
      end
      10'b1110010111 : begin
        result = input_919;
      end
      10'b1110011000 : begin
        result = input_920;
      end
      10'b1110011001 : begin
        result = input_921;
      end
      10'b1110011010 : begin
        result = input_922;
      end
      10'b1110011011 : begin
        result = input_923;
      end
      10'b1110011100 : begin
        result = input_924;
      end
      10'b1110011101 : begin
        result = input_925;
      end
      10'b1110011110 : begin
        result = input_926;
      end
      10'b1110011111 : begin
        result = input_927;
      end
      10'b1110100000 : begin
        result = input_928;
      end
      10'b1110100001 : begin
        result = input_929;
      end
      10'b1110100010 : begin
        result = input_930;
      end
      10'b1110100011 : begin
        result = input_931;
      end
      10'b1110100100 : begin
        result = input_932;
      end
      10'b1110100101 : begin
        result = input_933;
      end
      10'b1110100110 : begin
        result = input_934;
      end
      10'b1110100111 : begin
        result = input_935;
      end
      10'b1110101000 : begin
        result = input_936;
      end
      10'b1110101001 : begin
        result = input_937;
      end
      10'b1110101010 : begin
        result = input_938;
      end
      10'b1110101011 : begin
        result = input_939;
      end
      10'b1110101100 : begin
        result = input_940;
      end
      10'b1110101101 : begin
        result = input_941;
      end
      10'b1110101110 : begin
        result = input_942;
      end
      10'b1110101111 : begin
        result = input_943;
      end
      10'b1110110000 : begin
        result = input_944;
      end
      10'b1110110001 : begin
        result = input_945;
      end
      10'b1110110010 : begin
        result = input_946;
      end
      10'b1110110011 : begin
        result = input_947;
      end
      10'b1110110100 : begin
        result = input_948;
      end
      10'b1110110101 : begin
        result = input_949;
      end
      10'b1110110110 : begin
        result = input_950;
      end
      10'b1110110111 : begin
        result = input_951;
      end
      10'b1110111000 : begin
        result = input_952;
      end
      10'b1110111001 : begin
        result = input_953;
      end
      10'b1110111010 : begin
        result = input_954;
      end
      10'b1110111011 : begin
        result = input_955;
      end
      10'b1110111100 : begin
        result = input_956;
      end
      10'b1110111101 : begin
        result = input_957;
      end
      10'b1110111110 : begin
        result = input_958;
      end
      10'b1110111111 : begin
        result = input_959;
      end
      10'b1111000000 : begin
        result = input_960;
      end
      10'b1111000001 : begin
        result = input_961;
      end
      10'b1111000010 : begin
        result = input_962;
      end
      10'b1111000011 : begin
        result = input_963;
      end
      10'b1111000100 : begin
        result = input_964;
      end
      10'b1111000101 : begin
        result = input_965;
      end
      10'b1111000110 : begin
        result = input_966;
      end
      10'b1111000111 : begin
        result = input_967;
      end
      10'b1111001000 : begin
        result = input_968;
      end
      10'b1111001001 : begin
        result = input_969;
      end
      10'b1111001010 : begin
        result = input_970;
      end
      10'b1111001011 : begin
        result = input_971;
      end
      10'b1111001100 : begin
        result = input_972;
      end
      10'b1111001101 : begin
        result = input_973;
      end
      10'b1111001110 : begin
        result = input_974;
      end
      10'b1111001111 : begin
        result = input_975;
      end
      10'b1111010000 : begin
        result = input_976;
      end
      10'b1111010001 : begin
        result = input_977;
      end
      10'b1111010010 : begin
        result = input_978;
      end
      10'b1111010011 : begin
        result = input_979;
      end
      10'b1111010100 : begin
        result = input_980;
      end
      10'b1111010101 : begin
        result = input_981;
      end
      10'b1111010110 : begin
        result = input_982;
      end
      10'b1111010111 : begin
        result = input_983;
      end
      10'b1111011000 : begin
        result = input_984;
      end
      10'b1111011001 : begin
        result = input_985;
      end
      10'b1111011010 : begin
        result = input_986;
      end
      10'b1111011011 : begin
        result = input_987;
      end
      10'b1111011100 : begin
        result = input_988;
      end
      10'b1111011101 : begin
        result = input_989;
      end
      10'b1111011110 : begin
        result = input_990;
      end
      10'b1111011111 : begin
        result = input_991;
      end
      10'b1111100000 : begin
        result = input_992;
      end
      10'b1111100001 : begin
        result = input_993;
      end
      10'b1111100010 : begin
        result = input_994;
      end
      10'b1111100011 : begin
        result = input_995;
      end
      10'b1111100100 : begin
        result = input_996;
      end
      10'b1111100101 : begin
        result = input_997;
      end
      10'b1111100110 : begin
        result = input_998;
      end
      10'b1111100111 : begin
        result = input_999;
      end
      10'b1111101000 : begin
        result = input_1000;
      end
      10'b1111101001 : begin
        result = input_1001;
      end
      10'b1111101010 : begin
        result = input_1002;
      end
      10'b1111101011 : begin
        result = input_1003;
      end
      10'b1111101100 : begin
        result = input_1004;
      end
      10'b1111101101 : begin
        result = input_1005;
      end
      10'b1111101110 : begin
        result = input_1006;
      end
      10'b1111101111 : begin
        result = input_1007;
      end
      10'b1111110000 : begin
        result = input_1008;
      end
      10'b1111110001 : begin
        result = input_1009;
      end
      10'b1111110010 : begin
        result = input_1010;
      end
      10'b1111110011 : begin
        result = input_1011;
      end
      10'b1111110100 : begin
        result = input_1012;
      end
      10'b1111110101 : begin
        result = input_1013;
      end
      10'b1111110110 : begin
        result = input_1014;
      end
      10'b1111110111 : begin
        result = input_1015;
      end
      10'b1111111000 : begin
        result = input_1016;
      end
      10'b1111111001 : begin
        result = input_1017;
      end
      10'b1111111010 : begin
        result = input_1018;
      end
      10'b1111111011 : begin
        result = input_1019;
      end
      10'b1111111100 : begin
        result = input_1020;
      end
      10'b1111111101 : begin
        result = input_1021;
      end
      10'b1111111110 : begin
        result = input_1022;
      end
      default : begin
        result = input_1023;
      end
    endcase
    MUX_v_57_1024_2 = result;
  end
  endfunction


  function automatic [61:0] signext_62_57;
    input [56:0] vector;
  begin
    signext_62_57= {{5{vector[56]}}, vector};
  end
  endfunction

endmodule




//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ../td_ccore_solutions/leading_sign_57_0_1_0_86bc929c751c44a7dedde748d1abc423b086_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Mon May 27 10:59:57 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_57_0_1_0
// ------------------------------------------------------------------


module leading_sign_57_0_1_0 (
  mantissa, all_same, rtn
);
  input [56:0] mantissa;
  output all_same;
  output [5:0] rtn;


  // Interconnect Declarations
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_18_3_sdt_3;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_42_4_sdt_4;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_62_3_sdt_3;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_90_5_sdt_5;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_110_3_sdt_3;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_134_4_sdt_4;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_2;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_154_3_sdt_3;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_168_6_sdt_6;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_14_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_34_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_58_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_78_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_106_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_126_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_1;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_150_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_24;
  wire c_h_1_25;
  wire c_h_1_26;
  wire c_h_1_27;

  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_and_221_nl;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_and_219_nl;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_nl;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_or_4_nl;

  // Interconnect Declarations for Component Instantiations 
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_2 = ~((mantissa[54:53]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_1 = ~((mantissa[56:55]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_14_2_sdt_1 = ~((mantissa[52:51]!=2'b00));
  assign c_h_1_2 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_2;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_18_3_sdt_3 = (mantissa[50:49]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_14_2_sdt_1;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_2 = ~((mantissa[46:45]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_1 = ~((mantissa[48:47]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_34_2_sdt_1 = ~((mantissa[44:43]!=2'b00));
  assign c_h_1_5 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_18_3_sdt_3;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_42_4_sdt_4 = (mantissa[42:41]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_34_2_sdt_1 & c_h_1_5;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_2 = ~((mantissa[38:37]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_1 = ~((mantissa[40:39]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_58_2_sdt_1 = ~((mantissa[36:35]!=2'b00));
  assign c_h_1_9 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_2;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_62_3_sdt_3 = (mantissa[34:33]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_58_2_sdt_1;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_2 = ~((mantissa[30:29]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_1 = ~((mantissa[32:31]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_78_2_sdt_1 = ~((mantissa[28:27]!=2'b00));
  assign c_h_1_12 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_42_4_sdt_4;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_90_5_sdt_5 = (mantissa[26:25]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_78_2_sdt_1 & c_h_1_12
      & c_h_1_13;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_2 = ~((mantissa[22:21]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_1 = ~((mantissa[24:23]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_106_2_sdt_1 = ~((mantissa[20:19]!=2'b00));
  assign c_h_1_17 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_2;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_110_3_sdt_3 = (mantissa[18:17]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_106_2_sdt_1;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_2 = ~((mantissa[14:13]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_1 = ~((mantissa[16:15]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_126_2_sdt_1 = ~((mantissa[12:11]!=2'b00));
  assign c_h_1_20 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_110_3_sdt_3;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_134_4_sdt_4 = (mantissa[10:9]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_126_2_sdt_1 & c_h_1_20;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_2 = ~((mantissa[6:5]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_1 = ~((mantissa[8:7]!=2'b00));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_150_2_sdt_1 = ~((mantissa[4:3]!=2'b00));
  assign c_h_1_24 = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_1
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_2;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_154_3_sdt_3 = (mantissa[2:1]==2'b00)
      & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_150_2_sdt_1;
  assign c_h_1_25 = c_h_1_24 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_154_3_sdt_3;
  assign c_h_1_26 = c_h_1_21 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_134_4_sdt_4;
  assign c_h_1_27 = c_h_1_14 & return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_90_5_sdt_5;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_168_6_sdt_6 = (~
      (mantissa[0])) & c_h_1_25 & c_h_1_26 & c_h_1_27;
  assign all_same = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_168_6_sdt_6;
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_and_221_nl = c_h_1_14 &
      (c_h_1_26 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_90_5_sdt_5));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_and_219_nl = c_h_1_6 &
      (c_h_1_13 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_42_4_sdt_4))
      & (~((~(c_h_1_21 & (c_h_1_25 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_134_4_sdt_4))))
      & c_h_1_27));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_nl
      = c_h_1_2 & (c_h_1_5 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_18_3_sdt_3))
      & (~((~(c_h_1_9 & (c_h_1_12 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~((~(c_h_1_17 & (c_h_1_20 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_110_3_sdt_3))
      & (~((~(c_h_1_24 & (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_154_3_sdt_3)))
      & c_h_1_26)))) & c_h_1_27));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_1_nl
      = return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_1 & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_14_2_sdt_1
      | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_6_2_sdt_2)) & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_34_2_sdt_1 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_58_2_sdt_1 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_50_2_sdt_2))
      & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_1 &
      (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_78_2_sdt_1 | (~ return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_106_2_sdt_1 | (~
      return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_98_2_sdt_2)) & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_126_2_sdt_1 | (~
      return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_118_2_sdt_2)))) & c_h_1_21))
      & (~((~(return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_1
      & (return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_150_2_sdt_1 | (~
      return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_142_2_sdt_2)) & (~ c_h_1_25)))
      & c_h_1_26)))) & c_h_1_27));
  assign return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_or_4_nl
      = ((~((mantissa[56]) | (~((mantissa[55:54]!=2'b01))))) & (~(((mantissa[52])
      | (~((mantissa[51:50]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[48]) | (~((mantissa[47:46]!=2'b01)))))
      & (~(((mantissa[44]) | (~((mantissa[43:42]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[40]) | (~((mantissa[39:38]!=2'b01))))) & (~(((mantissa[36])
      | (~((mantissa[35:34]!=2'b01)))) & c_h_1_9)) & (~((~((~((mantissa[32]) | (~((mantissa[31:30]!=2'b01)))))
      & (~(((mantissa[28]) | (~((mantissa[27:26]!=2'b01)))) & c_h_1_12)))) & c_h_1_13))))
      & c_h_1_14)) & (~((~((~((mantissa[24]) | (~((mantissa[23:22]!=2'b01))))) &
      (~(((mantissa[20]) | (~((mantissa[19:18]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[16])
      | (~((mantissa[15:14]!=2'b01))))) & (~(((mantissa[12]) | (~((mantissa[11:10]!=2'b01))))
      & c_h_1_20)))) & c_h_1_21)) & (~(((mantissa[8]) | (~((mantissa[7:6]!=2'b01)))
      | (((mantissa[4]) | (~((mantissa[3:2]!=2'b01)))) & c_h_1_24) | c_h_1_25) &
      c_h_1_26)))) & c_h_1_27))) | return_add_generic_AC_RND_CONV_false_ls_all_sign_wrs_c_168_6_sdt_6;
  assign rtn = {c_h_1_27 , return_add_generic_AC_RND_CONV_false_ls_all_sign_and_221_nl
      , return_add_generic_AC_RND_CONV_false_ls_all_sign_and_219_nl , return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_nl
      , return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_and_1_nl
      , return_add_generic_AC_RND_CONV_false_ls_all_sign_return_add_generic_AC_RND_CONV_false_ls_all_sign_or_4_nl};
endmodule




//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/mgc_shift_r_beh_v5.v 
module mgc_shift_r_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

endmodule

//------> ../td_ccore_solutions/leading_sign_53_0_db1eac3e3536deac7d8d0fc62647951ea87c_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Mon May 27 10:59:48 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_53_0
// ------------------------------------------------------------------


module leading_sign_53_0 (
  mantissa, rtn
);
  input [52:0] mantissa;
  output [5:0] rtn;


  // Interconnect Declarations
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_18_3_sdt_3;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_42_4_sdt_4;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_62_3_sdt_3;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_90_5_sdt_5;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_110_3_sdt_3;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_134_4_sdt_4;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_2;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_14_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_34_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_58_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_78_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_106_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_126_2_sdt_1;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_23;
  wire c_h_1_24;
  wire c_h_1_25;

  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_205_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_216_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_3_nl;

  // Interconnect Declarations for Component Instantiations 
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_2
      = ~((mantissa[50:49]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_1
      = ~((mantissa[52:51]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_14_2_sdt_1
      = ~((mantissa[48:47]!=2'b00));
  assign c_h_1_2 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_2;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_18_3_sdt_3
      = (mantissa[46:45]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_14_2_sdt_1;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_2
      = ~((mantissa[42:41]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_1
      = ~((mantissa[44:43]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_34_2_sdt_1
      = ~((mantissa[40:39]!=2'b00));
  assign c_h_1_5 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_18_3_sdt_3;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_42_4_sdt_4
      = (mantissa[38:37]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_34_2_sdt_1
      & c_h_1_5;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_2
      = ~((mantissa[34:33]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_1
      = ~((mantissa[36:35]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_58_2_sdt_1
      = ~((mantissa[32:31]!=2'b00));
  assign c_h_1_9 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_2;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_62_3_sdt_3
      = (mantissa[30:29]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_58_2_sdt_1;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_2
      = ~((mantissa[26:25]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_1
      = ~((mantissa[28:27]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_78_2_sdt_1
      = ~((mantissa[24:23]!=2'b00));
  assign c_h_1_12 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_42_4_sdt_4;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_90_5_sdt_5
      = (mantissa[22:21]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_78_2_sdt_1
      & c_h_1_12 & c_h_1_13;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_2
      = ~((mantissa[18:17]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_1
      = ~((mantissa[20:19]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_106_2_sdt_1
      = ~((mantissa[16:15]!=2'b00));
  assign c_h_1_17 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_2;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_110_3_sdt_3
      = (mantissa[14:13]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_106_2_sdt_1;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_2
      = ~((mantissa[10:9]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_1
      = ~((mantissa[12:11]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_126_2_sdt_1
      = ~((mantissa[8:7]!=2'b00));
  assign c_h_1_20 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_110_3_sdt_3;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_134_4_sdt_4
      = (mantissa[6:5]==2'b00) & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_126_2_sdt_1
      & c_h_1_20;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_2
      = ~((mantissa[2:1]!=2'b00));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_1
      = ~((mantissa[4:3]!=2'b00));
  assign c_h_1_23 = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_1
      & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_2;
  assign c_h_1_24 = c_h_1_21 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_25 = c_h_1_14 & return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_90_5_sdt_5;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_205_nl
      = c_h_1_14 & (c_h_1_24 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_90_5_sdt_5));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_nl
      = c_h_1_6 & (c_h_1_13 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_42_4_sdt_4))
      & (~((~(c_h_1_21 & (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_134_4_sdt_4)))
      & c_h_1_25));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_216_nl
      = c_h_1_2 & (c_h_1_5 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_18_3_sdt_3))
      & (~((~(c_h_1_9 & (c_h_1_12 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~((~(c_h_1_17 & (c_h_1_20 | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_110_3_sdt_3))
      & (c_h_1_23 | (~ c_h_1_24)))) & c_h_1_25));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_1_nl
      = return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_14_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_34_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_58_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_50_2_sdt_2))
      & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_78_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_106_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_98_2_sdt_2))
      & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_1
      & (return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_126_2_sdt_1
      | (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_118_2_sdt_2))))
      & c_h_1_21)) & (~((~(return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_1
      & (~ return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_wrs_c_142_2_sdt_2)))
      & c_h_1_24)))) & c_h_1_25));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_3_nl
      = ((~((mantissa[52]) | (~((mantissa[51:50]!=2'b01))))) & (~(((mantissa[48])
      | (~((mantissa[47:46]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[44]) | (~((mantissa[43:42]!=2'b01)))))
      & (~(((mantissa[40]) | (~((mantissa[39:38]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[36]) | (~((mantissa[35:34]!=2'b01))))) & (~(((mantissa[32])
      | (~((mantissa[31:30]!=2'b01)))) & c_h_1_9)) & (~((~((~((mantissa[28]) | (~((mantissa[27:26]!=2'b01)))))
      & (~(((mantissa[24]) | (~((mantissa[23:22]!=2'b01)))) & c_h_1_12)))) & c_h_1_13))))
      & c_h_1_14)) & (~((~((~((mantissa[20]) | (~((mantissa[19:18]!=2'b01))))) &
      (~(((mantissa[16]) | (~((mantissa[15:14]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[12])
      | (~((mantissa[11:10]!=2'b01))))) & (~(((mantissa[8]) | (~((mantissa[7:6]!=2'b01))))
      & c_h_1_20)))) & c_h_1_21)) & (~(((mantissa[4]) | (~((mantissa[3:2]!=2'b01)))
      | c_h_1_23) & c_h_1_24)))) & c_h_1_25))) | ((~ (mantissa[0])) & c_h_1_23 &
      c_h_1_24 & c_h_1_25);
  assign rtn = {c_h_1_25 , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_205_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_216_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_1_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_3_nl};
endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   u110020015@ws41
//  Generated date: Mon May 27 12:39:13 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_7_16_10_1024_1024_16_5_gen
// ------------------------------------------------------------------


module stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_7_16_10_1024_1024_16_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [15:0] q;
  output we;
  output [15:0] d;
  output [9:0] adr;
  input [9:0] adr_d;
  input [15:0] d_d;
  input en_d;
  input we_d;
  output [15:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_6_64_10_1024_1024_64_5_gen
// ------------------------------------------------------------------


module stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_6_64_10_1024_1024_64_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [9:0] adr;
  input [9:0] adr_d;
  input [63:0] d_d;
  input en_d;
  input we_d;
  output [63:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_5_16_10_1024_1024_16_5_gen
// ------------------------------------------------------------------


module stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_5_16_10_1024_1024_16_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [15:0] q;
  output we;
  output [15:0] d;
  output [9:0] adr;
  input [9:0] adr_d;
  input [15:0] d_d;
  input en_d;
  input we_d;
  output [15:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_4_64_10_1024_1024_64_5_gen
// ------------------------------------------------------------------


module stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_4_64_10_1024_1024_64_5_gen
    (
  en, q, we, d, adr, adr_d, d_d, en_d, we_d, q_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  output en;
  input [63:0] q;
  output we;
  output [63:0] d;
  output [9:0] adr;
  input [9:0] adr_d;
  input [63:0] d_d;
  input en_d;
  input we_d;
  output [63:0] q_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign q_d = q;
  assign we = (port_0_rw_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module stage_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output, for_C_0_tr0, BUTTERFLY_C_24_tr0, BUTTERFLY_C_24_tr1,
      BUTTERFLY_1_C_24_tr0, BUTTERFLY_1_C_24_tr1, for_1_C_2_tr0
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [56:0] fsm_output;
  reg [56:0] fsm_output;
  input for_C_0_tr0;
  input BUTTERFLY_C_24_tr0;
  input BUTTERFLY_C_24_tr1;
  input BUTTERFLY_1_C_24_tr0;
  input BUTTERFLY_1_C_24_tr1;
  input for_1_C_2_tr0;


  // FSM State Type Declaration for stage_run_run_fsm_1
  parameter
    run_rlp_C_0 = 6'd0,
    main_C_0 = 6'd1,
    for_C_0 = 6'd2,
    BUTTERFLY_C_0 = 6'd3,
    BUTTERFLY_C_1 = 6'd4,
    BUTTERFLY_C_2 = 6'd5,
    BUTTERFLY_C_3 = 6'd6,
    BUTTERFLY_C_4 = 6'd7,
    BUTTERFLY_C_5 = 6'd8,
    BUTTERFLY_C_6 = 6'd9,
    BUTTERFLY_C_7 = 6'd10,
    BUTTERFLY_C_8 = 6'd11,
    BUTTERFLY_C_9 = 6'd12,
    BUTTERFLY_C_10 = 6'd13,
    BUTTERFLY_C_11 = 6'd14,
    BUTTERFLY_C_12 = 6'd15,
    BUTTERFLY_C_13 = 6'd16,
    BUTTERFLY_C_14 = 6'd17,
    BUTTERFLY_C_15 = 6'd18,
    BUTTERFLY_C_16 = 6'd19,
    BUTTERFLY_C_17 = 6'd20,
    BUTTERFLY_C_18 = 6'd21,
    BUTTERFLY_C_19 = 6'd22,
    BUTTERFLY_C_20 = 6'd23,
    BUTTERFLY_C_21 = 6'd24,
    BUTTERFLY_C_22 = 6'd25,
    BUTTERFLY_C_23 = 6'd26,
    BUTTERFLY_C_24 = 6'd27,
    BUTTERFLY_1_C_0 = 6'd28,
    BUTTERFLY_1_C_1 = 6'd29,
    BUTTERFLY_1_C_2 = 6'd30,
    BUTTERFLY_1_C_3 = 6'd31,
    BUTTERFLY_1_C_4 = 6'd32,
    BUTTERFLY_1_C_5 = 6'd33,
    BUTTERFLY_1_C_6 = 6'd34,
    BUTTERFLY_1_C_7 = 6'd35,
    BUTTERFLY_1_C_8 = 6'd36,
    BUTTERFLY_1_C_9 = 6'd37,
    BUTTERFLY_1_C_10 = 6'd38,
    BUTTERFLY_1_C_11 = 6'd39,
    BUTTERFLY_1_C_12 = 6'd40,
    BUTTERFLY_1_C_13 = 6'd41,
    BUTTERFLY_1_C_14 = 6'd42,
    BUTTERFLY_1_C_15 = 6'd43,
    BUTTERFLY_1_C_16 = 6'd44,
    BUTTERFLY_1_C_17 = 6'd45,
    BUTTERFLY_1_C_18 = 6'd46,
    BUTTERFLY_1_C_19 = 6'd47,
    BUTTERFLY_1_C_20 = 6'd48,
    BUTTERFLY_1_C_21 = 6'd49,
    BUTTERFLY_1_C_22 = 6'd50,
    BUTTERFLY_1_C_23 = 6'd51,
    BUTTERFLY_1_C_24 = 6'd52,
    for_1_C_0 = 6'd53,
    for_1_C_1 = 6'd54,
    for_1_C_2 = 6'd55,
    main_C_1 = 6'd56;

  reg [5:0] state_var;
  reg [5:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : stage_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000000000010;
        state_var_NS = for_C_0;
      end
      for_C_0 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000000000100;
        if ( for_C_0_tr0 ) begin
          state_var_NS = BUTTERFLY_C_0;
        end
        else begin
          state_var_NS = BUTTERFLY_1_C_0;
        end
      end
      BUTTERFLY_C_0 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000000001000;
        state_var_NS = BUTTERFLY_C_1;
      end
      BUTTERFLY_C_1 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000000010000;
        state_var_NS = BUTTERFLY_C_2;
      end
      BUTTERFLY_C_2 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000000100000;
        state_var_NS = BUTTERFLY_C_3;
      end
      BUTTERFLY_C_3 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000001000000;
        state_var_NS = BUTTERFLY_C_4;
      end
      BUTTERFLY_C_4 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000010000000;
        state_var_NS = BUTTERFLY_C_5;
      end
      BUTTERFLY_C_5 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000100000000;
        state_var_NS = BUTTERFLY_C_6;
      end
      BUTTERFLY_C_6 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000001000000000;
        state_var_NS = BUTTERFLY_C_7;
      end
      BUTTERFLY_C_7 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000010000000000;
        state_var_NS = BUTTERFLY_C_8;
      end
      BUTTERFLY_C_8 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000100000000000;
        state_var_NS = BUTTERFLY_C_9;
      end
      BUTTERFLY_C_9 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000001000000000000;
        state_var_NS = BUTTERFLY_C_10;
      end
      BUTTERFLY_C_10 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000010000000000000;
        state_var_NS = BUTTERFLY_C_11;
      end
      BUTTERFLY_C_11 : begin
        fsm_output = 57'b000000000000000000000000000000000000000000100000000000000;
        state_var_NS = BUTTERFLY_C_12;
      end
      BUTTERFLY_C_12 : begin
        fsm_output = 57'b000000000000000000000000000000000000000001000000000000000;
        state_var_NS = BUTTERFLY_C_13;
      end
      BUTTERFLY_C_13 : begin
        fsm_output = 57'b000000000000000000000000000000000000000010000000000000000;
        state_var_NS = BUTTERFLY_C_14;
      end
      BUTTERFLY_C_14 : begin
        fsm_output = 57'b000000000000000000000000000000000000000100000000000000000;
        state_var_NS = BUTTERFLY_C_15;
      end
      BUTTERFLY_C_15 : begin
        fsm_output = 57'b000000000000000000000000000000000000001000000000000000000;
        state_var_NS = BUTTERFLY_C_16;
      end
      BUTTERFLY_C_16 : begin
        fsm_output = 57'b000000000000000000000000000000000000010000000000000000000;
        state_var_NS = BUTTERFLY_C_17;
      end
      BUTTERFLY_C_17 : begin
        fsm_output = 57'b000000000000000000000000000000000000100000000000000000000;
        state_var_NS = BUTTERFLY_C_18;
      end
      BUTTERFLY_C_18 : begin
        fsm_output = 57'b000000000000000000000000000000000001000000000000000000000;
        state_var_NS = BUTTERFLY_C_19;
      end
      BUTTERFLY_C_19 : begin
        fsm_output = 57'b000000000000000000000000000000000010000000000000000000000;
        state_var_NS = BUTTERFLY_C_20;
      end
      BUTTERFLY_C_20 : begin
        fsm_output = 57'b000000000000000000000000000000000100000000000000000000000;
        state_var_NS = BUTTERFLY_C_21;
      end
      BUTTERFLY_C_21 : begin
        fsm_output = 57'b000000000000000000000000000000001000000000000000000000000;
        state_var_NS = BUTTERFLY_C_22;
      end
      BUTTERFLY_C_22 : begin
        fsm_output = 57'b000000000000000000000000000000010000000000000000000000000;
        state_var_NS = BUTTERFLY_C_23;
      end
      BUTTERFLY_C_23 : begin
        fsm_output = 57'b000000000000000000000000000000100000000000000000000000000;
        state_var_NS = BUTTERFLY_C_24;
      end
      BUTTERFLY_C_24 : begin
        fsm_output = 57'b000000000000000000000000000001000000000000000000000000000;
        if ( BUTTERFLY_C_24_tr0 ) begin
          state_var_NS = for_1_C_0;
        end
        else if ( BUTTERFLY_C_24_tr1 ) begin
          state_var_NS = BUTTERFLY_C_0;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      BUTTERFLY_1_C_0 : begin
        fsm_output = 57'b000000000000000000000000000010000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_1;
      end
      BUTTERFLY_1_C_1 : begin
        fsm_output = 57'b000000000000000000000000000100000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_2;
      end
      BUTTERFLY_1_C_2 : begin
        fsm_output = 57'b000000000000000000000000001000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_3;
      end
      BUTTERFLY_1_C_3 : begin
        fsm_output = 57'b000000000000000000000000010000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_4;
      end
      BUTTERFLY_1_C_4 : begin
        fsm_output = 57'b000000000000000000000000100000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_5;
      end
      BUTTERFLY_1_C_5 : begin
        fsm_output = 57'b000000000000000000000001000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_6;
      end
      BUTTERFLY_1_C_6 : begin
        fsm_output = 57'b000000000000000000000010000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_7;
      end
      BUTTERFLY_1_C_7 : begin
        fsm_output = 57'b000000000000000000000100000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_8;
      end
      BUTTERFLY_1_C_8 : begin
        fsm_output = 57'b000000000000000000001000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_9;
      end
      BUTTERFLY_1_C_9 : begin
        fsm_output = 57'b000000000000000000010000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_10;
      end
      BUTTERFLY_1_C_10 : begin
        fsm_output = 57'b000000000000000000100000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_11;
      end
      BUTTERFLY_1_C_11 : begin
        fsm_output = 57'b000000000000000001000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_12;
      end
      BUTTERFLY_1_C_12 : begin
        fsm_output = 57'b000000000000000010000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_13;
      end
      BUTTERFLY_1_C_13 : begin
        fsm_output = 57'b000000000000000100000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_14;
      end
      BUTTERFLY_1_C_14 : begin
        fsm_output = 57'b000000000000001000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_15;
      end
      BUTTERFLY_1_C_15 : begin
        fsm_output = 57'b000000000000010000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_16;
      end
      BUTTERFLY_1_C_16 : begin
        fsm_output = 57'b000000000000100000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_17;
      end
      BUTTERFLY_1_C_17 : begin
        fsm_output = 57'b000000000001000000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_18;
      end
      BUTTERFLY_1_C_18 : begin
        fsm_output = 57'b000000000010000000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_19;
      end
      BUTTERFLY_1_C_19 : begin
        fsm_output = 57'b000000000100000000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_20;
      end
      BUTTERFLY_1_C_20 : begin
        fsm_output = 57'b000000001000000000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_21;
      end
      BUTTERFLY_1_C_21 : begin
        fsm_output = 57'b000000010000000000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_22;
      end
      BUTTERFLY_1_C_22 : begin
        fsm_output = 57'b000000100000000000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_23;
      end
      BUTTERFLY_1_C_23 : begin
        fsm_output = 57'b000001000000000000000000000000000000000000000000000000000;
        state_var_NS = BUTTERFLY_1_C_24;
      end
      BUTTERFLY_1_C_24 : begin
        fsm_output = 57'b000010000000000000000000000000000000000000000000000000000;
        if ( BUTTERFLY_1_C_24_tr0 ) begin
          state_var_NS = for_1_C_0;
        end
        else if ( BUTTERFLY_1_C_24_tr1 ) begin
          state_var_NS = BUTTERFLY_1_C_0;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      for_1_C_0 : begin
        fsm_output = 57'b000100000000000000000000000000000000000000000000000000000;
        state_var_NS = for_1_C_1;
      end
      for_1_C_1 : begin
        fsm_output = 57'b001000000000000000000000000000000000000000000000000000000;
        state_var_NS = for_1_C_2;
      end
      for_1_C_2 : begin
        fsm_output = 57'b010000000000000000000000000000000000000000000000000000000;
        if ( for_1_C_2_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_1_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 57'b100000000000000000000000000000000000000000000000000000000;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 57'b000000000000000000000000000000000000000000000000000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_staller
// ------------------------------------------------------------------


module stage_run_staller (
  clk, rst, arst_n, run_wen, run_wten, ap_start_rsci_wen_comp, ap_done_rsci_wen_comp,
      out1_rsci_wen_comp
);
  input clk;
  input rst;
  input arst_n;
  output run_wen;
  output run_wten;
  reg run_wten;
  input ap_start_rsci_wen_comp;
  input ap_done_rsci_wen_comp;
  input out1_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = ap_start_rsci_wen_comp & ap_done_rsci_wen_comp & out1_rsci_wen_comp;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten <= 1'b0;
    end
    else if ( rst ) begin
      run_wten <= 1'b0;
    end
    else begin
      run_wten <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_out_u_triosy_obj_out_u_triosy_wait_ctrl
// ------------------------------------------------------------------


module stage_run_out_u_triosy_obj_out_u_triosy_wait_ctrl (
  run_wten, out_u_triosy_obj_iswt0, out_u_triosy_obj_biwt
);
  input run_wten;
  input out_u_triosy_obj_iswt0;
  output out_u_triosy_obj_biwt;



  // Interconnect Declarations for Component Instantiations 
  assign out_u_triosy_obj_biwt = (~ run_wten) & out_u_triosy_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_out_f_d_triosy_obj_out_f_d_triosy_wait_ctrl
// ------------------------------------------------------------------


module stage_run_out_f_d_triosy_obj_out_f_d_triosy_wait_ctrl (
  run_wten, out_f_d_triosy_obj_iswt0, out_f_d_triosy_obj_biwt
);
  input run_wten;
  input out_f_d_triosy_obj_iswt0;
  output out_f_d_triosy_obj_biwt;



  // Interconnect Declarations for Component Instantiations 
  assign out_f_d_triosy_obj_biwt = (~ run_wten) & out_f_d_triosy_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_in_u_triosy_obj_in_u_triosy_wait_ctrl
// ------------------------------------------------------------------


module stage_run_in_u_triosy_obj_in_u_triosy_wait_ctrl (
  run_wten, in_u_triosy_obj_iswt0, in_u_triosy_obj_biwt
);
  input run_wten;
  input in_u_triosy_obj_iswt0;
  output in_u_triosy_obj_biwt;



  // Interconnect Declarations for Component Instantiations 
  assign in_u_triosy_obj_biwt = (~ run_wten) & in_u_triosy_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_in_f_d_triosy_obj_in_f_d_triosy_wait_ctrl
// ------------------------------------------------------------------


module stage_run_in_f_d_triosy_obj_in_f_d_triosy_wait_ctrl (
  run_wten, in_f_d_triosy_obj_iswt0, in_f_d_triosy_obj_biwt
);
  input run_wten;
  input in_f_d_triosy_obj_iswt0;
  output in_f_d_triosy_obj_biwt;



  // Interconnect Declarations for Component Instantiations 
  assign in_f_d_triosy_obj_biwt = (~ run_wten) & in_f_d_triosy_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_mode1_triosy_obj_mode1_triosy_wait_ctrl
// ------------------------------------------------------------------


module stage_run_mode1_triosy_obj_mode1_triosy_wait_ctrl (
  run_wten, mode1_triosy_obj_iswt0, mode1_triosy_obj_biwt
);
  input run_wten;
  input mode1_triosy_obj_iswt0;
  output mode1_triosy_obj_biwt;



  // Interconnect Declarations for Component Instantiations 
  assign mode1_triosy_obj_biwt = (~ run_wten) & mode1_triosy_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_out1_rsci_out1_wait_ctrl
// ------------------------------------------------------------------


module stage_run_out1_rsci_out1_wait_ctrl (
  out1_rsci_iswt0, out1_rsci_biwt, out1_rsci_irdy
);
  input out1_rsci_iswt0;
  output out1_rsci_biwt;
  input out1_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign out1_rsci_biwt = out1_rsci_iswt0 & out1_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_wait_dp
// ------------------------------------------------------------------


module stage_run_wait_dp (
  in_f_d_rsci_en_d, in_u_rsci_en_d, out_f_d_rsci_en_d, out_u_rsci_en_d, run_wen,
      in_f_d_rsci_cgo, in_f_d_rsci_cgo_ir_unreg, in_u_rsci_cgo, in_u_rsci_cgo_ir_unreg,
      out_f_d_rsci_cgo, out_f_d_rsci_cgo_ir_unreg, out_u_rsci_cgo, out_u_rsci_cgo_ir_unreg
);
  output in_f_d_rsci_en_d;
  output in_u_rsci_en_d;
  output out_f_d_rsci_en_d;
  output out_u_rsci_en_d;
  input run_wen;
  input in_f_d_rsci_cgo;
  input in_f_d_rsci_cgo_ir_unreg;
  input in_u_rsci_cgo;
  input in_u_rsci_cgo_ir_unreg;
  input out_f_d_rsci_cgo;
  input out_f_d_rsci_cgo_ir_unreg;
  input out_u_rsci_cgo;
  input out_u_rsci_cgo_ir_unreg;



  // Interconnect Declarations for Component Instantiations 
  assign in_f_d_rsci_en_d = run_wen & (in_f_d_rsci_cgo | in_f_d_rsci_cgo_ir_unreg);
  assign in_u_rsci_en_d = run_wen & (in_u_rsci_cgo | in_u_rsci_cgo_ir_unreg);
  assign out_f_d_rsci_en_d = run_wen & (out_f_d_rsci_cgo | out_f_d_rsci_cgo_ir_unreg);
  assign out_u_rsci_en_d = run_wen & (out_u_rsci_cgo | out_u_rsci_cgo_ir_unreg);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_ap_done_rsci_ap_done_wait_ctrl
// ------------------------------------------------------------------


module stage_run_ap_done_rsci_ap_done_wait_ctrl (
  ap_done_rsci_iswt0, ap_done_rsci_biwt, ap_done_rsci_irdy
);
  input ap_done_rsci_iswt0;
  output ap_done_rsci_biwt;
  input ap_done_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign ap_done_rsci_biwt = ap_done_rsci_iswt0 & ap_done_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_ap_start_rsci_ap_start_wait_ctrl
// ------------------------------------------------------------------


module stage_run_ap_start_rsci_ap_start_wait_ctrl (
  ap_start_rsci_iswt0, ap_start_rsci_biwt, ap_start_rsci_ivld
);
  input ap_start_rsci_iswt0;
  output ap_start_rsci_biwt;
  input ap_start_rsci_ivld;



  // Interconnect Declarations for Component Instantiations 
  assign ap_start_rsci_biwt = ap_start_rsci_iswt0 & ap_start_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_out_u_triosy_obj
// ------------------------------------------------------------------


module stage_run_out_u_triosy_obj (
  out_u_triosy_lz, run_wten, out_u_triosy_obj_iswt0
);
  output out_u_triosy_lz;
  input run_wten;
  input out_u_triosy_obj_iswt0;


  // Interconnect Declarations
  wire out_u_triosy_obj_biwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) out_u_triosy_obj (
      .ld(out_u_triosy_obj_biwt),
      .lz(out_u_triosy_lz)
    );
  stage_run_out_u_triosy_obj_out_u_triosy_wait_ctrl stage_run_out_u_triosy_obj_out_u_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .out_u_triosy_obj_iswt0(out_u_triosy_obj_iswt0),
      .out_u_triosy_obj_biwt(out_u_triosy_obj_biwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_out_f_d_triosy_obj
// ------------------------------------------------------------------


module stage_run_out_f_d_triosy_obj (
  out_f_d_triosy_lz, run_wten, out_f_d_triosy_obj_iswt0
);
  output out_f_d_triosy_lz;
  input run_wten;
  input out_f_d_triosy_obj_iswt0;


  // Interconnect Declarations
  wire out_f_d_triosy_obj_biwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) out_f_d_triosy_obj (
      .ld(out_f_d_triosy_obj_biwt),
      .lz(out_f_d_triosy_lz)
    );
  stage_run_out_f_d_triosy_obj_out_f_d_triosy_wait_ctrl stage_run_out_f_d_triosy_obj_out_f_d_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .out_f_d_triosy_obj_iswt0(out_f_d_triosy_obj_iswt0),
      .out_f_d_triosy_obj_biwt(out_f_d_triosy_obj_biwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_in_u_triosy_obj
// ------------------------------------------------------------------


module stage_run_in_u_triosy_obj (
  in_u_triosy_lz, run_wten, in_u_triosy_obj_iswt0
);
  output in_u_triosy_lz;
  input run_wten;
  input in_u_triosy_obj_iswt0;


  // Interconnect Declarations
  wire in_u_triosy_obj_biwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) in_u_triosy_obj (
      .ld(in_u_triosy_obj_biwt),
      .lz(in_u_triosy_lz)
    );
  stage_run_in_u_triosy_obj_in_u_triosy_wait_ctrl stage_run_in_u_triosy_obj_in_u_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .in_u_triosy_obj_iswt0(in_u_triosy_obj_iswt0),
      .in_u_triosy_obj_biwt(in_u_triosy_obj_biwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_in_f_d_triosy_obj
// ------------------------------------------------------------------


module stage_run_in_f_d_triosy_obj (
  in_f_d_triosy_lz, run_wten, in_f_d_triosy_obj_iswt0
);
  output in_f_d_triosy_lz;
  input run_wten;
  input in_f_d_triosy_obj_iswt0;


  // Interconnect Declarations
  wire in_f_d_triosy_obj_biwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) in_f_d_triosy_obj (
      .ld(in_f_d_triosy_obj_biwt),
      .lz(in_f_d_triosy_lz)
    );
  stage_run_in_f_d_triosy_obj_in_f_d_triosy_wait_ctrl stage_run_in_f_d_triosy_obj_in_f_d_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .in_f_d_triosy_obj_iswt0(in_f_d_triosy_obj_iswt0),
      .in_f_d_triosy_obj_biwt(in_f_d_triosy_obj_biwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_mode1_triosy_obj
// ------------------------------------------------------------------


module stage_run_mode1_triosy_obj (
  mode1_triosy_lz, run_wten, mode1_triosy_obj_iswt0
);
  output mode1_triosy_lz;
  input run_wten;
  input mode1_triosy_obj_iswt0;


  // Interconnect Declarations
  wire mode1_triosy_obj_biwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) mode1_triosy_obj (
      .ld(mode1_triosy_obj_biwt),
      .lz(mode1_triosy_lz)
    );
  stage_run_mode1_triosy_obj_mode1_triosy_wait_ctrl stage_run_mode1_triosy_obj_mode1_triosy_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .mode1_triosy_obj_iswt0(mode1_triosy_obj_iswt0),
      .mode1_triosy_obj_biwt(mode1_triosy_obj_biwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_out1_rsci
// ------------------------------------------------------------------


module stage_run_out1_rsci (
  out1_rsc_dat, out1_rsc_vld, out1_rsc_rdy, out1_rsci_oswt, out1_rsci_wen_comp, out1_rsci_idat
);
  output [79:0] out1_rsc_dat;
  output out1_rsc_vld;
  input out1_rsc_rdy;
  input out1_rsci_oswt;
  output out1_rsci_wen_comp;
  input [79:0] out1_rsci_idat;


  // Interconnect Declarations
  wire out1_rsci_biwt;
  wire out1_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd8),
  .width(32'sd80)) out1_rsci (
      .irdy(out1_rsci_irdy),
      .ivld(out1_rsci_oswt),
      .idat(out1_rsci_idat),
      .rdy(out1_rsc_rdy),
      .vld(out1_rsc_vld),
      .dat(out1_rsc_dat)
    );
  stage_run_out1_rsci_out1_wait_ctrl stage_run_out1_rsci_out1_wait_ctrl_inst (
      .out1_rsci_iswt0(out1_rsci_oswt),
      .out1_rsci_biwt(out1_rsci_biwt),
      .out1_rsci_irdy(out1_rsci_irdy)
    );
  assign out1_rsci_wen_comp = (~ out1_rsci_oswt) | out1_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_ap_done_rsci
// ------------------------------------------------------------------


module stage_run_ap_done_rsci (
  ap_done_rsc_dat, ap_done_rsc_vld, ap_done_rsc_rdy, ap_done_rsci_oswt, ap_done_rsci_wen_comp
);
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input ap_done_rsci_oswt;
  output ap_done_rsci_wen_comp;


  // Interconnect Declarations
  wire ap_done_rsci_biwt;
  wire ap_done_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd1)) ap_done_rsci (
      .irdy(ap_done_rsci_irdy),
      .ivld(ap_done_rsci_oswt),
      .idat(1'b1),
      .rdy(ap_done_rsc_rdy),
      .vld(ap_done_rsc_vld),
      .dat(ap_done_rsc_dat)
    );
  stage_run_ap_done_rsci_ap_done_wait_ctrl stage_run_ap_done_rsci_ap_done_wait_ctrl_inst
      (
      .ap_done_rsci_iswt0(ap_done_rsci_oswt),
      .ap_done_rsci_biwt(ap_done_rsci_biwt),
      .ap_done_rsci_irdy(ap_done_rsci_irdy)
    );
  assign ap_done_rsci_wen_comp = (~ ap_done_rsci_oswt) | ap_done_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run_ap_start_rsci
// ------------------------------------------------------------------


module stage_run_ap_start_rsci (
  ap_start_rsc_dat, ap_start_rsc_vld, ap_start_rsc_rdy, ap_start_rsci_oswt, ap_start_rsci_wen_comp
);
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  input ap_start_rsci_oswt;
  output ap_start_rsci_wen_comp;


  // Interconnect Declarations
  wire ap_start_rsci_biwt;
  wire ap_start_rsci_ivld;
  wire ap_start_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd1)) ap_start_rsci (
      .rdy(ap_start_rsc_rdy),
      .vld(ap_start_rsc_vld),
      .dat(ap_start_rsc_dat),
      .irdy(ap_start_rsci_oswt),
      .ivld(ap_start_rsci_ivld),
      .idat(ap_start_rsci_idat)
    );
  stage_run_ap_start_rsci_ap_start_wait_ctrl stage_run_ap_start_rsci_ap_start_wait_ctrl_inst
      (
      .ap_start_rsci_iswt0(ap_start_rsci_oswt),
      .ap_start_rsci_biwt(ap_start_rsci_biwt),
      .ap_start_rsci_ivld(ap_start_rsci_ivld)
    );
  assign ap_start_rsci_wen_comp = (~ ap_start_rsci_oswt) | ap_start_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_run
// ------------------------------------------------------------------


module stage_run (
  clk, rst, arst_n, ap_start_rsc_dat, ap_start_rsc_vld, ap_start_rsc_rdy, ap_done_rsc_dat,
      ap_done_rsc_vld, ap_done_rsc_rdy, mode1_rsc_dat, mode1_triosy_lz, in_f_d_triosy_lz,
      in_u_triosy_lz, out_f_d_triosy_lz, out_u_triosy_lz, out1_rsc_dat, out1_rsc_vld,
      out1_rsc_rdy, in_f_d_rsci_adr_d, in_f_d_rsci_d_d, in_f_d_rsci_en_d, in_f_d_rsci_q_d,
      in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, in_u_rsci_adr_d, in_u_rsci_d_d,
      in_u_rsci_en_d, in_u_rsci_q_d, in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      out_f_d_rsci_adr_d, out_f_d_rsci_d_d, out_f_d_rsci_en_d, out_f_d_rsci_q_d,
      out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, out_u_rsci_adr_d, out_u_rsci_d_d,
      out_u_rsci_en_d, out_u_rsci_q_d, out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      in_f_d_rsci_we_d_pff, in_u_rsci_we_d_pff, out_f_d_rsci_we_d_pff, out_u_rsci_we_d_pff
);
  input clk;
  input rst;
  input arst_n;
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input [15:0] mode1_rsc_dat;
  output mode1_triosy_lz;
  output in_f_d_triosy_lz;
  output in_u_triosy_lz;
  output out_f_d_triosy_lz;
  output out_u_triosy_lz;
  output [79:0] out1_rsc_dat;
  output out1_rsc_vld;
  input out1_rsc_rdy;
  output [9:0] in_f_d_rsci_adr_d;
  output [63:0] in_f_d_rsci_d_d;
  output in_f_d_rsci_en_d;
  input [63:0] in_f_d_rsci_q_d;
  output in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [9:0] in_u_rsci_adr_d;
  output [15:0] in_u_rsci_d_d;
  output in_u_rsci_en_d;
  input [15:0] in_u_rsci_q_d;
  output in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [9:0] out_f_d_rsci_adr_d;
  output [63:0] out_f_d_rsci_d_d;
  output out_f_d_rsci_en_d;
  input [63:0] out_f_d_rsci_q_d;
  output out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [9:0] out_u_rsci_adr_d;
  output [15:0] out_u_rsci_d_d;
  output out_u_rsci_en_d;
  input [15:0] out_u_rsci_q_d;
  output out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output in_f_d_rsci_we_d_pff;
  output in_u_rsci_we_d_pff;
  output out_f_d_rsci_we_d_pff;
  output out_u_rsci_we_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire ap_start_rsci_wen_comp;
  wire ap_done_rsci_wen_comp;
  wire [15:0] mode1_rsci_idat;
  wire out1_rsci_wen_comp;
  reg [15:0] out1_rsci_idat_79_64;
  wire [56:0] fsm_output;
  wire return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_9_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_8_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_7_e1_eq_e2_equal_tmp;
  wire return_mult_generic_AC_RND_CONV_false_2_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_2_exp_ovf_oif_aelse_and_tmp;
  wire return_extract_19_return_extract_19_nor_tmp;
  wire return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp;
  wire operator_11_true_19_operator_11_true_19_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_tmp;
  wire return_mult_generic_AC_RND_CONV_false_1_exp_ovf_return_mult_generic_AC_RND_CONV_false_1_exp_ovf_or_tmp;
  wire return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_1_return_add_generic_AC_RND_CONV_false_6_op2_normal_return_extract_13_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_6_e1_eq_e2_equal_tmp;
  wire return_extract_13_m_zero_return_extract_13_m_zero_nor_tmp;
  wire operator_11_true_13_operator_11_true_13_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_tmp;
  wire return_mult_generic_AC_RND_CONV_false_exp_ovf_return_mult_generic_AC_RND_CONV_false_exp_ovf_or_tmp;
  wire return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp;
  wire return_extract_12_m_zero_return_extract_12_m_zero_nor_tmp;
  wire operator_11_true_12_operator_11_true_12_and_tmp;
  wire return_extract_2_and_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_1_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp;
  wire return_add_generic_AC_RND_CONV_false_e1_eq_e2_equal_tmp;
  wire operator_11_true_24_operator_11_true_24_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_if_1_return_add_generic_AC_RND_CONV_false_4_op2_normal_return_extract_9_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_or_tmp;
  wire [10:0] return_add_generic_AC_RND_CONV_false_4_e_dif_acc_tmp;
  wire [11:0] nl_return_add_generic_AC_RND_CONV_false_4_e_dif_acc_tmp;
  wire return_add_generic_AC_RND_CONV_false_4_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_23_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_22_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp;
  wire return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp;
  wire return_mult_generic_AC_RND_CONV_false_5_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_5_exp_ovf_oif_aelse_and_tmp;
  wire return_extract_51_return_extract_51_nor_tmp;
  wire return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp;
  wire operator_11_true_51_operator_11_true_51_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp;
  wire return_mult_generic_AC_RND_CONV_false_4_exp_ovf_return_mult_generic_AC_RND_CONV_false_4_exp_ovf_or_tmp;
  wire return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_tmp;
  wire return_add_generic_AC_RND_CONV_false_19_e1_eq_e2_equal_tmp;
  wire return_extract_45_m_zero_return_extract_45_m_zero_nor_tmp;
  wire operator_11_true_45_operator_11_true_45_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp;
  wire return_mult_generic_AC_RND_CONV_false_3_exp_ovf_return_mult_generic_AC_RND_CONV_false_3_exp_ovf_or_tmp;
  wire return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp;
  wire return_extract_44_m_zero_return_extract_44_m_zero_nor_tmp;
  wire operator_11_true_44_operator_11_true_44_and_tmp;
  wire return_add_generic_AC_RND_CONV_false_14_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_15_aif_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp;
  wire return_add_generic_AC_RND_CONV_false_13_return_add_generic_AC_RND_CONV_false_13_or_1_tmp;
  wire operator_11_true_33_operator_11_true_33_and_tmp;
  wire BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_tmp;
  wire stage_PE_1_and_1_tmp;
  wire operator_16_false_operator_16_false_nor_tmp;
  wire or_dcpl_11;
  wire and_dcpl_1;
  wire or_dcpl_48;
  wire and_dcpl_28;
  wire or_dcpl_49;
  wire and_dcpl_32;
  wire and_dcpl_36;
  wire and_dcpl_63;
  wire and_dcpl_128;
  wire and_dcpl_129;
  wire and_dcpl_135;
  wire and_dcpl_138;
  wire or_dcpl_75;
  wire or_dcpl_79;
  wire or_dcpl_87;
  wire and_dcpl_140;
  wire and_dcpl_146;
  wire or_dcpl_92;
  wire or_dcpl_95;
  wire or_dcpl_99;
  wire or_dcpl_101;
  wire or_dcpl_102;
  wire or_dcpl_105;
  wire or_dcpl_106;
  wire or_dcpl_108;
  wire and_dcpl_151;
  wire and_dcpl_152;
  wire or_dcpl_115;
  wire or_dcpl_118;
  wire or_dcpl_125;
  wire or_dcpl_126;
  wire or_dcpl_128;
  wire or_dcpl_132;
  wire or_dcpl_133;
  wire or_dcpl_135;
  wire or_dcpl_136;
  wire and_dcpl_165;
  wire or_dcpl_148;
  wire or_dcpl_159;
  wire or_dcpl_163;
  wire or_dcpl_166;
  wire and_dcpl_166;
  wire or_dcpl_185;
  wire or_dcpl_187;
  wire and_dcpl_168;
  wire or_dcpl_199;
  wire or_dcpl_201;
  wire or_dcpl_203;
  wire or_dcpl_207;
  wire or_dcpl_211;
  wire or_dcpl_214;
  wire or_dcpl_216;
  wire or_dcpl_219;
  wire or_dcpl_224;
  wire or_dcpl_225;
  wire or_dcpl_228;
  wire or_dcpl_231;
  wire or_dcpl_234;
  wire or_dcpl_235;
  wire or_dcpl_237;
  wire or_dcpl_240;
  wire or_dcpl_242;
  wire or_dcpl_244;
  wire or_dcpl_249;
  wire or_dcpl_252;
  wire or_dcpl_261;
  wire or_dcpl_275;
  wire or_dcpl_278;
  wire or_dcpl_282;
  wire or_dcpl_287;
  wire or_dcpl_289;
  wire or_dcpl_296;
  wire or_dcpl_302;
  wire or_dcpl_395;
  wire and_dcpl_210;
  wire and_dcpl_211;
  wire and_dcpl_213;
  wire and_dcpl_214;
  wire and_dcpl_217;
  wire or_dcpl_397;
  wire and_dcpl_233;
  wire and_dcpl_236;
  wire or_dcpl_401;
  wire or_dcpl_404;
  wire or_dcpl_406;
  wire or_dcpl_407;
  wire or_dcpl_415;
  wire or_dcpl_417;
  wire or_dcpl_418;
  wire or_dcpl_420;
  wire or_dcpl_421;
  wire or_dcpl_422;
  wire or_dcpl_423;
  wire or_dcpl_424;
  wire or_dcpl_425;
  wire and_dcpl_241;
  wire or_dcpl_431;
  wire or_dcpl_438;
  wire or_dcpl_440;
  wire or_dcpl_444;
  wire or_dcpl_445;
  wire or_dcpl_447;
  wire or_dcpl_449;
  wire or_dcpl_461;
  wire or_dcpl_462;
  wire or_dcpl_464;
  wire or_dcpl_465;
  wire or_dcpl_466;
  wire and_dcpl_257;
  wire and_dcpl_258;
  wire and_dcpl_259;
  wire and_dcpl_260;
  wire and_dcpl_261;
  wire and_dcpl_262;
  wire and_dcpl_263;
  wire and_dcpl_264;
  wire and_dcpl_265;
  wire and_dcpl_266;
  wire or_dcpl_488;
  wire and_dcpl_267;
  wire and_dcpl_268;
  wire or_dcpl_493;
  wire or_dcpl_495;
  wire or_dcpl_500;
  wire or_dcpl_501;
  wire or_dcpl_502;
  wire or_dcpl_503;
  wire or_dcpl_511;
  wire or_dcpl_512;
  wire or_dcpl_513;
  wire or_dcpl_514;
  wire or_dcpl_517;
  wire or_dcpl_518;
  wire or_dcpl_519;
  wire and_dcpl_284;
  wire and_dcpl_286;
  wire or_dcpl_531;
  wire or_dcpl_534;
  wire or_dcpl_542;
  wire and_dcpl_326;
  wire or_dcpl_548;
  wire or_dcpl_549;
  wire or_dcpl_550;
  wire or_dcpl_551;
  wire or_dcpl_552;
  wire or_dcpl_553;
  wire or_dcpl_556;
  wire or_dcpl_557;
  wire or_dcpl_558;
  wire or_dcpl_560;
  wire or_dcpl_561;
  wire or_dcpl_566;
  wire or_dcpl_568;
  wire or_dcpl_570;
  wire or_dcpl_571;
  wire or_dcpl_573;
  wire or_dcpl_574;
  wire or_dcpl_575;
  wire or_dcpl_576;
  wire or_dcpl_579;
  wire or_dcpl_580;
  wire or_dcpl_586;
  wire or_dcpl_587;
  wire or_dcpl_597;
  wire or_dcpl_607;
  wire or_dcpl_610;
  wire or_dcpl_618;
  wire or_dcpl_628;
  wire or_dcpl_631;
  wire or_dcpl_660;
  wire or_dcpl_661;
  wire or_dcpl_662;
  wire or_dcpl_666;
  wire or_dcpl_682;
  wire or_dcpl_693;
  wire or_dcpl_694;
  wire or_dcpl_697;
  wire or_dcpl_704;
  wire or_dcpl_705;
  wire or_dcpl_707;
  wire or_dcpl_712;
  wire or_dcpl_713;
  wire or_dcpl_716;
  wire or_dcpl_719;
  wire or_dcpl_722;
  wire or_dcpl_736;
  wire or_dcpl_749;
  wire or_dcpl_750;
  wire or_dcpl_751;
  wire or_dcpl_769;
  wire or_dcpl_776;
  wire or_dcpl_780;
  wire or_dcpl_788;
  wire or_dcpl_789;
  wire or_dcpl_790;
  wire or_dcpl_793;
  wire or_dcpl_799;
  wire or_dcpl_803;
  wire or_dcpl_840;
  wire and_dcpl_348;
  wire and_dcpl_349;
  wire or_dcpl_863;
  wire or_dcpl_870;
  wire or_dcpl_876;
  wire or_dcpl_882;
  wire or_dcpl_906;
  wire or_dcpl_911;
  wire or_dcpl_912;
  wire or_dcpl_913;
  wire or_dcpl_914;
  wire or_dcpl_919;
  wire or_dcpl_928;
  wire or_dcpl_929;
  wire or_dcpl_937;
  wire or_dcpl_940;
  wire or_dcpl_949;
  wire or_dcpl_953;
  wire or_dcpl_961;
  wire or_dcpl_976;
  wire or_dcpl_985;
  wire or_dcpl_999;
  wire or_dcpl_1001;
  wire or_dcpl_1015;
  wire or_dcpl_1069;
  wire and_dcpl_385;
  wire not_tmp_302;
  wire and_dcpl_399;
  wire and_dcpl_408;
  wire and_dcpl_413;
  wire or_tmp_61;
  wire or_tmp_82;
  wire or_tmp_83;
  wire or_tmp_112;
  wire or_tmp_113;
  wire or_tmp_208;
  wire or_tmp_234;
  wire or_tmp_261;
  wire or_tmp_348;
  wire or_tmp_403;
  wire or_tmp_440;
  wire or_tmp_561;
  wire or_tmp_564;
  wire or_tmp_570;
  wire or_tmp_771;
  wire or_tmp_823;
  wire or_tmp_852;
  wire or_tmp_857;
  wire and_592_cse;
  wire and_571_cse;
  wire and_666_cse;
  wire and_1013_cse;
  wire and_1608_cse;
  wire and_1598_cse;
  wire and_1163_cse;
  wire and_2281_cse;
  reg for_i_0_sva;
  wire return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_6_lor_lpi_2_dfm_1;
  wire return_extract_3_m_zero_sva_mx1w0;
  wire return_mult_generic_AC_RND_CONV_false_6_op1_nan_sva_1;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3;
  wire return_mult_generic_AC_RND_CONV_false_6_e_incr_lpi_2_dfm_2;
  wire return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_or_2;
  wire return_add_generic_AC_RND_CONV_false_12_exception_sva_1;
  reg operator_11_true_return_24_sva;
  reg return_add_generic_AC_RND_CONV_false_10_op1_inf_sva;
  reg return_add_generic_AC_RND_CONV_false_10_op2_inf_sva;
  reg return_add_generic_AC_RND_CONV_false_10_op1_nan_sva;
  reg return_add_generic_AC_RND_CONV_false_10_op2_nan_sva;
  wire return_add_generic_AC_RND_CONV_false_12_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_12_else_4_unequal_tmp;
  reg return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  wire return_add_generic_AC_RND_CONV_false_11_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva;
  reg return_add_generic_AC_RND_CONV_false_23_op1_inf_sva;
  reg return_add_generic_AC_RND_CONV_false_14_op2_inf_sva;
  reg return_add_generic_AC_RND_CONV_false_23_op1_nan_sva;
  reg return_add_generic_AC_RND_CONV_false_14_op2_nan_sva;
  wire return_add_generic_AC_RND_CONV_false_11_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_10_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  wire return_add_generic_AC_RND_CONV_false_10_op2_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_10_op2_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_10_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_10_else_4_unequal_tmp;
  reg operator_11_true_return_15_sva;
  reg return_extract_17_m_zero_sva;
  wire return_add_generic_AC_RND_CONV_false_9_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_9_op2_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_9_op2_nan_sva_mx7w0;
  wire return_add_generic_AC_RND_CONV_false_9_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_9_else_4_unequal_tmp;
  reg operator_11_true_return_1_sva;
  reg return_extract_15_m_zero_sva;
  wire return_add_generic_AC_RND_CONV_false_8_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1;
  reg operator_11_true_return_26_sva;
  reg return_extract_26_m_zero_sva;
  wire return_add_generic_AC_RND_CONV_false_8_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_8_op1_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_8_op1_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_8_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_8_else_4_unequal_tmp;
  reg operator_11_true_return_17_sva;
  reg return_extract_1_m_zero_sva;
  wire [11:0] return_add_generic_AC_RND_CONV_false_9_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1;
  reg return_extract_24_m_zero_sva;
  wire return_add_generic_AC_RND_CONV_false_7_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_7_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva_mx1;
  wire return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1;
  reg return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm;
  reg return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm;
  reg [49:0] return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm;
  wire return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_8_e_dif_qr_lpi_3_dfm_mx0;
  reg return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm;
  reg return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm;
  wire return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_2_m_r_51_lpi_3_dfm_mx1;
  wire [50:0] return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_2_zero_m_return_mult_generic_AC_RND_CONV_false_2_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_2_r_zero_return_mult_generic_AC_RND_CONV_false_2_r_zero_nor_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_2_lor_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_2_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_2_r_nan_sva_1;
  reg return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_or_2;
  wire return_add_generic_AC_RND_CONV_false_6_exception_sva_1;
  reg return_add_generic_AC_RND_CONV_false_22_op1_inf_sva;
  wire return_add_generic_AC_RND_CONV_false_6_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp;
  wire drf_qr_lval_14_smx_0_lpi_3_dfm_mx1;
  wire [50:0] return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_1_zero_m_return_mult_generic_AC_RND_CONV_false_1_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_1_r_zero_return_mult_generic_AC_RND_CONV_false_1_r_zero_nor_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_1_lor_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_6_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_1_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_1_r_nan_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_1_op2_zero_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_1_e_incr_lpi_3_dfm_2;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_or_2;
  wire return_add_generic_AC_RND_CONV_false_6_op2_nan_sva_1;
  reg return_extract_17_return_extract_17_nor_cse_sva;
  reg return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm;
  wire return_add_generic_AC_RND_CONV_false_6_op2_mu_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_50_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_49_0_mx0;
  wire return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_6_e_dif_qr_lpi_3_dfm_mx0;
  reg return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm;
  wire stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0;
  wire return_add_generic_AC_RND_CONV_false_3_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_3_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_11_mux_2_itm_mx3;
  wire [50:0] return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_zero_m_return_mult_generic_AC_RND_CONV_false_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_r_zero_return_mult_generic_AC_RND_CONV_false_r_zero_nor_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_lor_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_6_op1_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_r_nan_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_op2_zero_sva_1;
  wire [11:0] return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_e_incr_lpi_3_dfm_2;
  wire return_mult_generic_AC_RND_CONV_false_if_1_aelse_return_mult_generic_AC_RND_CONV_false_if_1_aelse_or_2;
  wire return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1;
  wire return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_1;
  reg return_extract_15_return_extract_15_nor_cse_sva;
  wire return_add_generic_AC_RND_CONV_false_2_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_2_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_2_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_1_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_9_op1_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_1_op1_nan_sva_mx3w0;
  wire return_add_generic_AC_RND_CONV_false_9_op1_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_1_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_1_else_4_unequal_tmp;
  wire [10:0] drf_qr_lval_1_smx_lpi_3_dfm_mx1;
  wire [11:0] return_add_generic_AC_RND_CONV_false_1_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_else_4_unequal_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_4_m_r_51_lpi_3_dfm_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1;
  reg inverse_lpi_1_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_17_do_sub_sva_1;
  wire return_add_generic_AC_RND_CONV_false_25_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_25_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_25_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_24_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_24_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_24_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_23_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_23_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_23_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_22_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_22_op2_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_22_op2_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_22_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_22_else_4_unequal_tmp;
  wire [11:0] return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_21_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1;
  reg return_add_generic_AC_RND_CONV_false_11_mux_itm;
  wire return_add_generic_AC_RND_CONV_false_21_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_21_op1_inf_sva_1;
  wire return_add_generic_AC_RND_CONV_false_21_op1_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_21_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_21_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_20_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_20_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_20_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva_mx2;
  wire return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2;
  reg drf_qr_lval_13_smx_0_lpi_3_dfm;
  wire return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_mx1;
  wire [50:0] return_mult_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_5_zero_m_return_mult_generic_AC_RND_CONV_false_5_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_5_r_zero_return_mult_generic_AC_RND_CONV_false_5_r_zero_nor_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_5_lor_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_5_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_5_r_nan_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_or_2;
  wire return_add_generic_AC_RND_CONV_false_19_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_19_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_11_mux_2_itm_mx9;
  wire [50:0] return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_4_zero_m_return_mult_generic_AC_RND_CONV_false_4_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_4_r_zero_return_mult_generic_AC_RND_CONV_false_4_r_zero_nor_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_4_lor_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_4_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_4_r_nan_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_4_op1_zero_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_4_op2_zero_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_4_e_incr_lpi_3_dfm_2;
  wire return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_or_2;
  wire return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_19_op2_mu_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0_mx0;
  wire return_add_generic_AC_RND_CONV_false_19_op2_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_16_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_16_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_16_else_4_unequal_tmp;
  wire drf_qr_lval_14_smx_0_lpi_3_dfm_mx3;
  wire [50:0] return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_3_zero_m_return_mult_generic_AC_RND_CONV_false_3_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_3_r_zero_return_mult_generic_AC_RND_CONV_false_3_r_zero_nor_mdf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_3_lor_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_3_op2_inf_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_3_r_nan_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_3_op1_zero_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_3_e_incr_lpi_3_dfm_2;
  wire return_mult_generic_AC_RND_CONV_false_3_if_1_aelse_return_mult_generic_AC_RND_CONV_false_3_if_1_aelse_or_2;
  wire return_add_generic_AC_RND_CONV_false_19_op1_nan_sva_1;
  wire return_add_generic_AC_RND_CONV_false_15_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_15_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_15_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_14_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_14_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_14_else_4_unequal_tmp;
  wire [10:0] drf_qr_lval_11_smx_lpi_3_dfm_mx2;
  wire return_add_generic_AC_RND_CONV_false_13_exception_sva_1;
  wire return_add_generic_AC_RND_CONV_false_13_r_inf_lpi_3_dfm_2;
  reg return_add_generic_AC_RND_CONV_false_13_else_4_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm_1;
  wire operator_16_false_1_operator_16_false_1_and_mdf_sva_1;
  reg operator_16_false_operator_16_false_nor_cse_sva;
  reg t_in_10_0_lpi_1_dfm_1_10;
  reg t_in_10_0_lpi_1_dfm_1_9;
  reg mode_lpi_1_dfm;
  reg [9:0] BUTTERFLY_1_n_9_0_sva_1;
  reg BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm;
  reg [15:0] operator_16_false_io_read_mode1_rsc_cse_sva;
  reg [12:0] operator_33_true_12_acc_psp_sva;
  reg return_add_generic_AC_RND_CONV_false_10_do_sub_sva;
  reg return_add_generic_AC_RND_CONV_false_16_do_sub_sva;
  reg return_add_generic_AC_RND_CONV_false_11_do_sub_sva;
  reg return_add_generic_AC_RND_CONV_false_12_do_sub_sva;
  reg return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva;
  wire return_add_generic_AC_RND_CONV_false_mux_28;
  wire [9:0] return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1;
  reg [63:0] stage_PE_1_x_im_d_sva;
  reg [63:0] stage_PE_1_x_re_d_sva;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1;
  reg return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva;
  wire stage_d_mul_return_d_4_63_sva_1;
  wire stage_d_mul_return_d_2_63_sva_1;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w3;
  wire stage_d_mul_return_d_63_sva_1;
  reg return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1;
  reg return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva;
  wire [9:0] return_add_generic_AC_RND_CONV_false_4_e_r_qelse_qr_10_1_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1;
  reg return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva;
  wire stage_d_mul_return_d_5_63_sva_1;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_4_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w2;
  reg return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva;
  wire [10:0] return_mult_generic_AC_RND_CONV_false_3_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w6;
  reg return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva;
  wire [9:0] return_add_generic_AC_RND_CONV_false_5_e_r_qelse_qr_10_1_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_17_e_r_qelse_qr_10_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_if_5_or_3;
  reg reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd;
  wire for_1_if_and_ssc;
  reg out1_rsci_idat_63;
  reg [10:0] out1_rsci_idat_62_52;
  reg out1_rsci_idat_51;
  reg [50:0] out1_rsci_idat_50_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_11_e_dif_qr_lpi_3_dfm_mx0_10_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_3_e_dif_qr_lpi_3_dfm_mx0_10_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_2_e_dif_qr_lpi_3_dfm_mx0_10_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt;
  wire [11:0] nl_return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt;
  wire [9:0] return_add_generic_AC_RND_CONV_false_4_e_dif_qif_acc_pmx_lpi_3_dfm_mx0_9_0;
  wire [10:0] return_add_generic_AC_RND_CONV_false_25_e_dif_qr_lpi_3_dfm_mx0_10_0;
  wire stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0;
  wire stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0;
  wire or_1670_ssc;
  wire or_1673_ssc;
  wire or_1678_ssc;
  reg reg_out_u_triosy_obj_iswt0_cse;
  reg reg_out1_rsci_iswt0_cse;
  reg reg_out_u_rsci_cgo_ir_cse;
  reg reg_out_f_d_rsci_cgo_ir_cse;
  reg reg_in_u_rsci_cgo_ir_cse;
  reg reg_in_f_d_rsci_cgo_ir_cse;
  reg reg_ap_start_rsci_iswt0_cse;
  wire operator_16_false_and_cse;
  wire t_in_and_cse;
  wire mode_and_cse;
  wire stage_PE_1_and_2_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_cse;
  wire BUTTERFLY_1_n_and_cse;
  wire return_extract_17_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_9_op1_smaller_return_add_generic_AC_RND_CONV_false_9_op1_smaller_or_cse;
  wire return_add_generic_AC_RND_CONV_false_10_r_zero_and_cse;
  wire return_add_generic_AC_RND_CONV_false_22_op1_mu_and_cse;
  wire return_add_generic_AC_RND_CONV_false_23_op1_nan_and_cse;
  wire return_add_generic_AC_RND_CONV_false_22_op1_smaller_return_add_generic_AC_RND_CONV_false_22_op1_smaller_or_cse;
  wire return_add_generic_AC_RND_CONV_false_10_op2_nan_and_cse;
  wire return_add_generic_AC_RND_CONV_false_12_op_bigger_and_2_cse;
  wire return_add_generic_AC_RND_CONV_false_12_op_smaller_and_1_cse;
  wire [50:0] stage_PE_1_gm_re_d_mux_cse;
  wire stage_PE_1_gm_im_d_mux_cse;
  wire [50:0] stage_PE_1_gm_im_d_mux_2_cse;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_6_cse;
  wire or_590_cse;
  wire xor_cse;
  wire return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse;
  wire xor_2_cse;
  wire xor_3_cse;
  wire xor_4_cse;
  wire return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse;
  wire and_2333_cse;
  wire or_1144_cse;
  wire return_add_generic_AC_RND_CONV_false_3_r_nan_mux1h_cse;
  wire or_918_cse;
  wire and_2331_cse;
  wire return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse;
  wire [50:0] return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse;
  wire return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse;
  wire return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse;
  wire and_2332_cse;
  wire return_add_generic_AC_RND_CONV_false_16_r_nan_mux1h_cse;
  wire or_920_cse;
  wire return_add_generic_AC_RND_CONV_false_25_op1_smaller_return_add_generic_AC_RND_CONV_false_25_op1_smaller_or_cse;
  wire stage_PE_1_and_cse;
  wire and_83_cse;
  wire nor_3_cse;
  wire or_46_cse;
  wire nor_24_cse;
  wire and_416_cse;
  wire return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_and_cse;
  wire return_add_generic_AC_RND_CONV_false_9_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_9_op1_smaller_oelse_and_cse;
  wire return_add_generic_AC_RND_CONV_false_20_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_20_op1_smaller_oelse_and_cse;
  wire return_add_generic_AC_RND_CONV_false_22_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_22_op1_smaller_oelse_and_cse;
  wire return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_and_cse;
  wire return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_and_cse;
  wire and_522_cse;
  wire or_38_cse;
  wire return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_and_cse;
  wire and_470_cse;
  wire and_468_cse;
  reg drf_qr_lval_14_smx_0_lpi_3_dfm;
  reg return_add_generic_AC_RND_CONV_false_11_mux_2_itm;
  wire [50:0] stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0;
  wire [50:0] stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0;
  reg [50:0] return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm;
  wire return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_10_op2_mu_1_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_10_op2_mu_1_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1;
  reg return_add_generic_AC_RND_CONV_false_22_op1_mu_52_lpi_3_dfm;
  reg [50:0] return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm;
  wire return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_op2_mu_52_lpi_3_dfm_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx1;
  wire return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_17_op1_mu_52_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_17_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_17_op2_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_20_op2_mu_1_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_20_op2_mu_1_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_20_op2_mu_1_0_lpi_3_dfm_1;
  wire or_1205_ssc;
  wire or_1206_ssc;
  wire and_654_ssc;
  wire or_1208_ssc;
  wire or_1209_ssc;
  wire or_1231_ssc;
  wire or_1232_ssc;
  wire or_1233_ssc;
  wire or_1234_ssc;
  wire and_720_ssc;
  wire and_494_m1c;
  wire return_add_generic_AC_RND_CONV_false_12_res_mant_and_ssc;
  reg [6:0] return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_56_50;
  reg [49:0] return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_49_0;
  wire stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0;
  wire stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0;
  wire BUTTERFLY_1_else_3_else_and_ssc;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  wire and_2334_cse;
  wire return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_and_1_cse;
  wire return_add_generic_AC_RND_CONV_false_8_op1_smaller_return_add_generic_AC_RND_CONV_false_8_op1_smaller_or_cse;
  wire return_add_generic_AC_RND_CONV_false_7_op1_smaller_return_add_generic_AC_RND_CONV_false_7_op1_smaller_or_cse;
  wire return_add_generic_AC_RND_CONV_false_20_op1_smaller_return_add_generic_AC_RND_CONV_false_20_op1_smaller_or_cse;
  wire return_add_generic_AC_RND_CONV_false_13_op1_mu_52_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_4_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire BUTTERFLY_1_fiy_mux1h_2_cse;
  wire BUTTERFLY_1_fiy_mux1h_6_cse;
  wire or_200_cse;
  wire return_add_generic_AC_RND_CONV_false_10_exp_mux1h_8_cse;
  wire return_add_generic_AC_RND_CONV_false_10_exp_mux1h_11_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_21_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_27_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_6_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_12_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_31_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_34_cse;
  wire return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_2_cse;
  wire return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_3_cse;
  wire return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_cse;
  wire return_add_generic_AC_RND_CONV_false_5_op_smaller_mux_cse;
  wire return_add_generic_AC_RND_CONV_false_22_op1_mu_mux_cse;
  wire return_add_generic_AC_RND_CONV_false_22_op1_mu_mux_1_cse;
  wire return_add_generic_AC_RND_CONV_false_10_exp_mux_5_cse;
  wire return_add_generic_AC_RND_CONV_false_5_op_smaller_mux_1_cse;
  wire return_add_generic_AC_RND_CONV_false_1_op_bigger_mux_4_cse;
  wire return_add_generic_AC_RND_CONV_false_13_mux_25_cse;
  wire return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_2_cse;
  wire return_add_generic_AC_RND_CONV_false_1_op_bigger_mux_5_cse;
  wire nor_158_cse;
  wire return_extract_26_exception_or_3_cse;
  wire stage_PE_1_tmp_re_d_and_ssc;
  reg [6:0] stage_PE_1_tmp_re_d_1_sva_1_63_57;
  wire [5:0] stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_5;
  wire [3:0] stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_4_1;
  wire [5:0] stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_5;
  wire [3:0] stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_4_1;
  wire or_219_cse;
  wire stage_PE_1_tmp_re_d_1_sva_1_mx0c0;
  wire or_1181_rmff;
  wire or_1180_rmff;
  wire or_1179_rmff;
  wire or_1178_rmff;
  reg return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva;
  reg return_add_generic_AC_RND_CONV_false_12_mux_itm;
  reg return_add_generic_AC_RND_CONV_false_17_mux_6_itm;
  wire [9:0] return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_11;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
  wire return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx1w0;
  reg return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs;
  wire return_add_generic_AC_RND_CONV_false_1_mux_32;
  wire return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs_mx1w0;
  reg return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs;
  wire return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_9;
  reg return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_10_unequal_tmp;
  wire return_add_generic_AC_RND_CONV_false_13_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_22_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_23_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_24_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_25_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_14_or_1_svs_1;
  reg [9:0] BUTTERFLY_1_i_9_0_sva;
  reg [9:0] BUTTERFLY_1_fry_9_0_sva;
  reg BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm;
  reg return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs;
  wire return_add_generic_AC_RND_CONV_false_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_9_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_10_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_11_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_12_or_1_svs_1;
  wire return_add_generic_AC_RND_CONV_false_1_or_1_svs_1;
  reg [1:0] BUTTERFLY_1_else_3_else_acc_4_itm_15_14;
  wire [14:0] stage_monty_mul_acc_2_psp_sva_1;
  wire [15:0] nl_stage_monty_mul_acc_2_psp_sva_1;
  wire or_tmp;
  wire or_tmp_916;
  wire or_tmp_917;
  wire or_tmp_919;
  wire or_tmp_920;
  wire or_tmp_921;
  wire or_tmp_922;
  wire or_tmp_924;
  wire [9:0] return_add_generic_AC_RND_CONV_false_e_r_return_add_generic_AC_RND_CONV_false_e_r_or_cse;
  wire [9:0] return_add_generic_AC_RND_CONV_false_1_e_r_return_add_generic_AC_RND_CONV_false_1_e_r_or_cse;
  wire [9:0] drf_qr_lval_4_smx_9_0_lpi_3_dfm_mx0;
  wire [9:0] stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w3_10_1;
  wire [9:0] stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w9_10_1;
  reg [5:0] return_add_generic_AC_RND_CONV_false_12_ls_sva;
  reg [9:0] drf_qr_lval_13_smx_10_1_lpi_3_dfm;
  reg [5:0] return_add_generic_AC_RND_CONV_false_10_ls_sva;
  reg [9:0] drf_qr_lval_14_smx_10_1_lpi_3_dfm;
  reg [5:0] return_add_generic_AC_RND_CONV_false_11_ls_sva;
  wire nor_160_m1c;
  wire nor_161_m1c;
  wire nor_162_m1c;
  wire nor_163_m1c;
  wire BUTTERFLY_if_1_if_and_9_cse;
  wire BUTTERFLY_if_1_if_and_5_cse;
  wire BUTTERFLY_if_1_if_and_11_cse;
  wire BUTTERFLY_if_1_if_and_8_cse;
  wire BUTTERFLY_if_1_if_and_10_cse;
  wire BUTTERFLY_if_1_if_and_6_cse;
  wire BUTTERFLY_if_1_and_7_cse;
  wire BUTTERFLY_if_1_and_11_cse;
  wire BUTTERFLY_if_1_and_13_cse;
  wire BUTTERFLY_if_1_and_10_cse;
  wire BUTTERFLY_if_1_and_12_cse;
  wire BUTTERFLY_if_1_and_8_cse;
  wire BUTTERFLY_if_1_if_or_1_cse;
  wire BUTTERFLY_if_1_or_1_cse;
  wire [50:0] return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_itm;
  wire [50:0] return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_1_itm;
  wire [50:0] return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_2_itm;
  wire [50:0] return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_7_itm;
  wire [50:0] return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_8_itm;
  wire [13:0] BUTTERFLY_1_else_3_else_mux1h_itm;
  wire or_1540_itm;
  wire return_add_generic_AC_RND_CONV_false_13_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_13_op1_smaller_oelse_and_1_itm;
  wire [5:0] return_add_generic_AC_RND_CONV_false_4_mux_10_itm;
  wire [5:0] return_add_generic_AC_RND_CONV_false_17_mux_10_itm;
  wire or_tmp_927;
  wire or_tmp_929;
  wire or_tmp_930;
  wire [11:0] z_out_1;
  wire or_tmp_940;
  wire [9:0] z_out_2;
  wire [10:0] nl_z_out_2;
  wire [17:0] z_out_3;
  wire [18:0] nl_z_out_3;
  wire [15:0] z_out_5;
  wire [16:0] nl_z_out_5;
  wire [53:0] z_out_6;
  wire [54:0] nl_z_out_6;
  wire or_tmp_979;
  wire [9:0] z_out_7;
  wire [10:0] nl_z_out_7;
  wire or_tmp_983;
  wire [12:0] z_out_8;
  wire [13:0] nl_z_out_8;
  wire [63:0] O_1_out;
  wire [61:0] O_1_out_1;
  wire [9:0] z_out_9;
  wire [9:0] z_out_10;
  wire [50:0] z_out_11;
  wire [56:0] z_out_15;
  wire [54:0] z_out_16;
  wire [54:0] z_out_17;
  wire [105:0] z_out_18;
  wire all_same_out;
  wire [5:0] rtn_out;
  wire [10:0] z_out_19;
  wire [11:0] nl_z_out_19;
  wire [9:0] z_out_20;
  wire [10:0] nl_z_out_20;
  wire [105:0] z_out_21;
  wire signed [107:0] nl_z_out_21;
  wire [11:0] z_out_23;
  wire [11:0] z_out_24;
  wire [11:0] z_out_25;
  wire [11:0] z_out_26;
  wire [12:0] z_out_27;
  wire [10:0] z_out_28;
  wire [12:0] z_out_29;
  wire [56:0] z_out_30;
  wire [11:0] z_out_36;
  wire [12:0] nl_z_out_36;
  wire [17:0] z_out_37;
  wire [15:0] z_out_38;
  wire [16:0] nl_z_out_38;
  wire [11:0] z_out_39;
  wire [16:0] z_out_40;
  wire [53:0] z_out_42;
  wire or_tmp_1248;
  wire or_tmp_1249;
  wire or_tmp_1250;
  wire or_tmp_1251;
  wire [56:0] z_out_43;
  wire [5:0] rtn_out_1;
  wire [11:0] z_out_44;
  wire [17:0] z_out_45;
  wire [18:0] nl_z_out_45;
  reg return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm;
  reg return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm;
  reg return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_52_lpi_3_dfm;
  reg return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_51_lpi_3_dfm;
  reg return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm;
  reg drf_qr_lval_15_smx_0_lpi_3_dfm;
  reg [5:0] return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva;
  reg stage_PE_1_index_const_15_lpi_2_dfm;
  reg stage_PE_1_index_const_10_lpi_2_dfm;
  reg stage_PE_1_index_const_0_lpi_2_dfm;
  reg stage_PE_1_qr_0_lpi_2_dfm;
  reg stage_PE_1_qr_1_0_lpi_2_dfm;
  reg [61:0] stage_PE_1_gm_im_d_61_0_lpi_3_dfm;
  reg [5:0] return_add_generic_AC_RND_CONV_false_15_e_dif_sat_sva;
  reg return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_18_e_r_qr_0_lpi_3_dfm;
  reg [50:0] return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm;
  reg return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs;
  reg return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm;
  reg return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_itm;
  reg return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm;
  reg return_add_generic_AC_RND_CONV_false_18_mux_itm;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_8;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_7;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_8;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_8;
  reg [51:0] return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0;
  wire out1_rsci_idat_63_0_mx0c1;
  wire out1_rsci_idat_63_0_mx0c2;
  wire out1_rsci_idat_79_64_mx0c1;
  wire mode_lpi_1_dfm_mx0w0;
  wire [8:0] BUTTERFLY_i_div_psp_sva_1;
  wire return_extract_15_return_extract_15_nor_cse_sva_mx1;
  wire return_add_generic_AC_RND_CONV_false_15_r_nan_or_mx2w0;
  wire return_extract_15_return_extract_15_nor_cse_sva_mx2;
  wire return_add_generic_AC_RND_CONV_false_4_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_4_e_r_qelse_or_svs_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_4_e_dif_sat_sva_1;
  wire [9:0] BUTTERFLY_i_9_0_sva_1;
  wire [10:0] nl_BUTTERFLY_i_9_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx1;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx5;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx6;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx1;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx2;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx6;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx7;
  wire return_extract_9_return_extract_9_or_1_cse_sva_1;
  wire return_add_generic_AC_RND_CONV_false_9_if_2_return_add_generic_AC_RND_CONV_false_9_if_2_and_1_mx2w0;
  wire return_add_generic_AC_RND_CONV_false_12_if_2_return_add_generic_AC_RND_CONV_false_12_if_2_nor_mx4w0;
  wire return_add_generic_AC_RND_CONV_false_7_if_2_return_add_generic_AC_RND_CONV_false_7_if_2_and_1_mx1w0;
  wire return_add_generic_AC_RND_CONV_false_8_if_2_return_add_generic_AC_RND_CONV_false_8_if_2_and_1_mx2w0;
  wire [5:0] return_add_generic_AC_RND_CONV_false_2_e_dif_sat_sva_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx6c1;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx6c2;
  wire operator_11_true_return_17_sva_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_5_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_svs_1;
  wire return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm_mx1;
  wire return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm_mx4;
  wire return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm_mx0w4;
  wire stage_PE_1_tmp_im_d_1_sva_1_mx0c3;
  wire return_add_generic_AC_RND_CONV_false_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_2_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_11_if_2_return_add_generic_AC_RND_CONV_false_11_if_2_nor_mx2w0;
  wire return_add_generic_AC_RND_CONV_false_10_if_2_return_add_generic_AC_RND_CONV_false_10_if_2_and_1_mx5w0;
  wire return_add_generic_AC_RND_CONV_false_6_do_sub_sva_1;
  wire return_add_generic_AC_RND_CONV_false_2_r_nan_and_2;
  wire stage_PE_1_tmp_re_d_1_sva_1_mx0c4;
  wire [50:0] return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_1_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_3_res_mant_3_0_sva_1;
  wire [50:0] stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0w0;
  wire [50:0] stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0;
  wire [9:0] return_add_generic_AC_RND_CONV_false_2_e_r_qelse_qr_10_1_lpi_3_dfm_1;
  wire [52:0] return_mult_generic_AC_RND_CONV_false_res_bef_rnd_3_53_1_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_if_1_and_1_tmp_1;
  wire return_extract_12_return_extract_12_or_1_cse_sva_1;
  wire [50:0] stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx0w3;
  wire [50:0] stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1;
  wire [50:0] stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0w0;
  wire [9:0] return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_50_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0;
  wire return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_6_res_mant_3_0_sva_1;
  wire [52:0] return_mult_generic_AC_RND_CONV_false_1_res_bef_rnd_3_53_1_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_tmp_1;
  wire return_extract_13_return_extract_13_or_1_cse_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_6_e_dif_sat_sva_1;
  wire return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_52_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_51_lpi_3_dfm_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_mult_generic_AC_RND_CONV_false_2_e_incr_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_7_res_mant_3_0_sva_1;
  wire [52:0] return_mult_generic_AC_RND_CONV_false_2_res_bef_rnd_3_53_1_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_2_if_1_and_1_tmp_1;
  wire return_extract_19_return_extract_19_or_sva_1;
  wire return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_51_lpi_3_dfm_mx3;
  wire return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_52_lpi_3_dfm_mx3;
  wire [5:0] return_add_generic_AC_RND_CONV_false_9_e_dif_sat_sva_1;
  wire [49:0] return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_8_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_9_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_11_res_mant_3_0_sva_1;
  wire [49:0] return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_10_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_12_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_17_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_17_e_r_qelse_or_svs_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_13_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_15_res_mant_3_0_sva_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_14_res_mant_3_0_sva_1;
  wire return_add_generic_AC_RND_CONV_false_16_res_mant_3_0_sva_1;
  wire [52:0] return_mult_generic_AC_RND_CONV_false_3_res_bef_rnd_3_53_1_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_3_if_1_and_1_tmp_1;
  wire return_extract_44_return_extract_44_or_1_cse_sva_1;
  wire [50:0] stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0w0;
  wire return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_50_mx0;
  wire [49:0] return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0;
  wire return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_0_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_19_res_mant_3_0_sva_1;
  wire [52:0] return_mult_generic_AC_RND_CONV_false_4_res_bef_rnd_3_53_1_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_4_if_1_and_1_tmp_1;
  wire return_extract_45_return_extract_45_or_1_cse_sva_1;
  wire [49:0] return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_mult_generic_AC_RND_CONV_false_5_e_incr_lpi_3_dfm_2;
  wire return_add_generic_AC_RND_CONV_false_20_res_mant_3_0_sva_1;
  wire [52:0] return_mult_generic_AC_RND_CONV_false_5_res_bef_rnd_3_53_1_lpi_3_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_5_if_1_and_1_tmp_1;
  wire return_extract_51_return_extract_51_or_sva_1;
  wire return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0;
  wire [50:0] return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1;
  wire [9:0] return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1;
  wire return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1;
  wire [49:0] return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_22_res_mant_3_0_sva_1;
  wire [49:0] return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0;
  wire return_add_generic_AC_RND_CONV_false_23_res_mant_3_0_sva_1;
  wire [5:0] return_add_generic_AC_RND_CONV_false_23_e_dif_sat_sva_1;
  wire return_add_generic_AC_RND_CONV_false_25_res_mant_3_0_sva_1;
  wire return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1;
  wire [52:0] return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1;
  wire return_mult_generic_AC_RND_CONV_false_6_if_1_and_1_tmp_1;
  wire [14:0] operator_32_false_2_acc_psp_1_sva_1;
  wire [15:0] nl_operator_32_false_2_acc_psp_1_sva_1;
  wire return_add_generic_AC_RND_CONV_false_5_sticky_bit_and_54;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_54;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_56;
  wire return_add_generic_AC_RND_CONV_false_6_mux_35;
  wire return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_nor_2;
  wire return_add_generic_AC_RND_CONV_false_12_sticky_bit_and_54;
  wire return_add_generic_AC_RND_CONV_false_12_sticky_bit_and_56;
  wire return_add_generic_AC_RND_CONV_false_12_sticky_bit_and_58;
  wire stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w3_0;
  wire stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w9_0;
  wire stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx1_50;
  wire stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx2_50;
  wire stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50;
  wire [9:0] stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1;
  wire stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50;
  wire [9:0] stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_0;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_0;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_0;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_0;
  wire [13:0] U_ROM_1i10_1o14_out_2;
  wire [13:0] U_ROM_1i10_1o14_out_3;
  wire [55:0] return_add_generic_AC_RND_CONV_false_res_mant_conc_2_itm_56_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_conc_6_itm_54_4;
  wire [49:0] return_add_generic_AC_RND_CONV_false_23_conc_6_itm_53_4;
  wire [55:0] return_add_generic_AC_RND_CONV_false_1_res_mant_conc_2_itm_56_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_1_conc_6_itm_54_4;
  wire [49:0] return_add_generic_AC_RND_CONV_false_6_conc_6_itm_53_4;
  wire [55:0] return_add_generic_AC_RND_CONV_false_8_res_mant_conc_7_itm_56_1;
  wire [49:0] return_add_generic_AC_RND_CONV_false_10_conc_6_itm_53_4;
  wire [55:0] return_add_generic_AC_RND_CONV_false_14_res_mant_conc_2_itm_56_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_14_conc_6_itm_54_4;
  wire [49:0] return_add_generic_AC_RND_CONV_false_19_conc_6_itm_53_4;
  wire [55:0] return_add_generic_AC_RND_CONV_false_13_res_mant_conc_2_itm_56_1;
  wire [50:0] return_add_generic_AC_RND_CONV_false_13_conc_6_itm_54_4;
  wire [51:0] return_mult_generic_AC_RND_CONV_false_6_if_conc_itm_51_0;
  wire operator_6_false_or_ssc;
  wire operator_6_false_or_1_ssc;
  wire return_add_generic_AC_RND_CONV_false_4_or_ssc;
  reg [4:0] BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0;
  reg [1:0] BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1;
  reg [8:0] BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2;
  wire BUTTERFLY_1_else_1_if_and_ssc;
  reg return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_0;
  reg [49:0] return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1;
  wire return_add_generic_AC_RND_CONV_false_15_op_bigger_and_ssc;
  reg return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_0;
  reg [49:0] return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1;
  wire return_add_generic_AC_RND_CONV_false_17_m_r_and_ssc;
  reg [5:0] BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_0;
  reg BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_1;
  reg [2:0] BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_0;
  reg BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1;
  wire BUTTERFLY_1_else_3_else_and_1_ssc;
  reg [6:0] stage_PE_1_tmp_im_d_1_sva_1_rsp_0;
  reg [56:0] stage_PE_1_tmp_im_d_1_sva_1_rsp_1;
  wire stage_PE_1_tmp_im_d_and_ssc;
  reg [5:0] stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_0;
  reg [50:0] stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_1;
  wire [5:0] stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5;
  wire [3:0] stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1;
  wire [5:0] stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5;
  wire [3:0] stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1;
  wire [5:0] drf_qr_lval_smx_lpi_3_dfm_mx0_10_5;
  wire [4:0] drf_qr_lval_smx_lpi_3_dfm_mx0_4_0;
  wire [5:0] drf_qr_lval_16_smx_lpi_3_dfm_mx0_10_5;
  wire [4:0] drf_qr_lval_16_smx_lpi_3_dfm_mx0_4_0;
  wire operator_6_false_1_or_1_ssc;
  wire operator_6_false_or_3_ssc;
  wire return_add_generic_AC_RND_CONV_false_4_or_20_ssc;
  wire return_add_generic_AC_RND_CONV_false_4_or_18_ssc;
  wire [4:0] return_add_generic_AC_RND_CONV_false_mux_26_itm_4_0;
  wire [4:0] return_add_generic_AC_RND_CONV_false_13_mux_28_itm_4_0;
  wire return_add_generic_AC_RND_CONV_false_e_dif1_or_1_ssc;
  wire return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_nor_cse;
  wire return_extract_15_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_9_e_dif_qelse_return_add_generic_AC_RND_CONV_false_9_e_dif_qelse_and_cse;
  wire [51:0] return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
  wire return_add_generic_AC_RND_CONV_false_4_if_5_return_add_generic_AC_RND_CONV_false_4_if_5_nor_cse;
  wire [11:0] return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_or_2_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_149_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_141_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_133_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_125_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_117_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_109_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_101_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_93_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_85_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_77_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_69_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_61_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_155_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_147_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_139_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_131_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_123_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_115_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_107_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_99_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_91_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_83_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_75_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_67_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_59_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_153_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_145_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_137_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_129_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_121_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_113_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_105_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_97_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_89_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_81_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_73_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_65_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_57_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_151_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_143_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_135_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_127_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_119_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_111_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_103_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_95_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_87_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_79_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_71_cse;
  wire return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_63_cse;
  wire return_add_generic_AC_RND_CONV_false_4_sticky_bit_and_cse;
  wire return_add_generic_AC_RND_CONV_false_4_sticky_bit_and_52_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_2_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_6_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_7_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_8_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_9_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_10_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_11_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_12_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_13_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_14_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_15_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_16_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_17_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_18_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_19_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_20_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_21_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_22_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_23_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_24_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_25_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_26_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_27_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_28_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_29_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_30_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_31_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_32_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_33_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_34_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_35_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_36_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_37_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_38_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_39_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_40_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_41_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_42_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_43_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_44_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_45_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_46_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_47_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_48_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_49_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_50_cse;
  wire return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_51_cse;
  wire return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse;
  wire [55:0] return_add_generic_AC_RND_CONV_false_5_mux_19_cse;
  wire [55:0] return_add_generic_AC_RND_CONV_false_5_mux_18_cse;
  wire [55:0] return_add_generic_AC_RND_CONV_false_6_mux_33_cse;
  wire [55:0] return_add_generic_AC_RND_CONV_false_12_mux_19_cse;
  wire [55:0] return_add_generic_AC_RND_CONV_false_12_mux_21_cse;
  wire [55:0] return_add_generic_AC_RND_CONV_false_5_mux_20_cse;
  wire [55:0] return_add_generic_AC_RND_CONV_false_4_mux_24_cse;
  wire [1:0] BUTTERFLY_else_1_BUTTERFLY_else_1_and_cse;
  wire return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_or_cse;
  wire operator_6_false_8_nor_1_cse;
  wire and_1153_rgt;
  wire return_add_generic_AC_RND_CONV_false_10_or_cse;
  wire [5:0] return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_cse;
  wire [5:0] return_add_generic_AC_RND_CONV_false_21_e_dif_sat_or_cse;
  wire return_mult_generic_AC_RND_CONV_false_exp_ovf_oif_aelse_nor_cse;
  wire return_mult_generic_AC_RND_CONV_false_if_or_3_cse;
  wire [3:0] return_mult_generic_AC_RND_CONV_false_if_nand_1_cse;
  wire return_mult_generic_AC_RND_CONV_false_if_or_cse;
  wire [5:0] return_add_generic_AC_RND_CONV_false_8_e_dif_sat_or_cse;
  wire [5:0] return_add_generic_AC_RND_CONV_false_e_dif_sat_or_cse;
  wire nand_12_cse;
  wire return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse;
  wire operator_6_false_1_or_8_cse;
  wire operator_6_false_1_or_4_cse;
  wire operator_6_false_1_or_6_cse;
  wire operator_6_false_or_15_cse;
  wire operator_6_false_or_6_cse;
  wire operator_6_false_or_12_cse;
  wire BUTTERFLY_i_nor_2_cse_1;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_or_6_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_35_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_33_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_43_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_47_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_27_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_31_cse;
  wire return_add_generic_AC_RND_CONV_false_12_res_mant_or_cse;
  wire operator_6_false_or_20_cse;
  wire return_add_generic_AC_RND_CONV_false_20_ma1_lt_ma2_mux_1_cse;
  wire [50:0] return_add_generic_AC_RND_CONV_false_20_ma1_lt_ma2_mux_4_cse;
  wire BUTTERFLY_1_else_1_if_BUTTERFLY_1_else_1_if_mux_2_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_86_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_87_cse;
  wire return_extract_15_m_zero_mux1h_cse;
  wire return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse;
  wire return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse;
  wire return_extract_1_exception_or_cse;
  wire return_add_generic_AC_RND_CONV_false_4_res_rounded_or_1_cse;
  wire return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_or_1_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_99_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_105_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_97_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_95_cse;
  wire BUTTERFLY_i_or_4_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_13_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_52_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_7_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_15_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_54_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_9_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_17_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_56_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_11_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_19_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_67_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_71_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_77_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_73_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_70_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_69_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_75_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_73_cse;
  wire and_1615_cse;
  wire and_1583_cse;
  wire and_1584_cse;
  wire and_1626_cse;
  wire return_extract_26_m_zero_sva_2;
  wire or_1375_cse;
  wire return_add_generic_AC_RND_CONV_false_8_exp_and_ssc;
  reg drf_qr_lval_11_smx_lpi_3_dfm_10;
  reg drf_qr_lval_11_smx_lpi_3_dfm_9;
  reg m_in_15_1_lpi_1_dfm_1_1;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_1;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_1;
  reg reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd;
  reg [3:0] reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1;
  reg [3:0] reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2;
  reg reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3;
  wire return_add_generic_AC_RND_CONV_false_17_and_2_m1c;
  wire return_add_generic_AC_RND_CONV_false_17_and_4_m1c;
  wire return_add_generic_AC_RND_CONV_false_17_and_6_m1c;
  wire return_extract_32_or_1_tmp;
  wire and_453_tmp;
  wire return_add_generic_AC_RND_CONV_false_11_and_24_m1c;
  wire return_add_generic_AC_RND_CONV_false_11_and_28_m1c;
  wire and_491_tmp;
  wire and_497_tmp;
  wire return_extract_26_exception_and_5_m1c;
  wire return_extract_26_exception_and_7_m1c;
  wire return_extract_26_exception_and_10_m1c;
  wire return_extract_26_exception_and_12_m1c;
  wire return_add_generic_AC_RND_CONV_false_12_and_2_m1c;
  wire return_add_generic_AC_RND_CONV_false_12_and_6_m1c;
  reg [4:0] reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd;
  reg [4:0] reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_1;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_1;
  reg m_in_15_1_lpi_1_dfm_1_2;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_2;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_2;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_6_cse;
  wire BUTTERFLY_1_fiy_or_1_cse;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_or_3_rgt;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_or_8_rgt;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_or_9_rgt;
  wire [4:0] return_add_generic_AC_RND_CONV_false_1_mux_25_itm_4_0;
  reg [3:0] drf_qr_lval_11_smx_lpi_3_dfm_8_5;
  reg [4:0] drf_qr_lval_11_smx_lpi_3_dfm_4_0;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_2;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_2;
  reg m_in_15_1_lpi_1_dfm_1_3;
  wire [4:0] return_add_generic_AC_RND_CONV_false_3_mux_16_mx0_4_0;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_3;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_3;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_7_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_11_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_7_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_16_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_12_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_13_cse;
  wire return_add_generic_AC_RND_CONV_false_17_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_17_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_23_cse;
  wire return_extract_26_exception_and_6_cse;
  wire return_extract_26_exception_and_11_cse;
  wire return_add_generic_AC_RND_CONV_false_11_exp_and_2_cse;
  wire return_add_generic_AC_RND_CONV_false_11_exp_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_10_exp_and_2_cse;
  wire return_add_generic_AC_RND_CONV_false_10_exp_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_14_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_and_15_cse;
  wire return_add_generic_AC_RND_CONV_false_10_exp_and_6_cse;
  wire return_add_generic_AC_RND_CONV_false_10_exp_and_7_cse;
  wire return_add_generic_AC_RND_CONV_false_10_exp_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_12_op_bigger_and_8_cse;
  wire return_add_generic_AC_RND_CONV_false_12_op_bigger_and_9_cse;
  wire return_add_generic_AC_RND_CONV_false_10_exp_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse;
  wire return_add_generic_AC_RND_CONV_false_17_e_r_and_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_34_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse;
  wire BUTTERFLY_1_else_2_or_cse;
  wire BUTTERFLY_1_else_2_and_27_cse;
  wire BUTTERFLY_1_else_3_else_and_11_cse;
  wire BUTTERFLY_1_else_3_else_or_rgt;
  wire stage_PE_1_tmp_re_d_or_4_rgt;
  wire stage_PE_1_tmp_re_d_and_5_rgt;
  wire stage_PE_1_tmp_re_d_and_7_rgt;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_3;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_3;
  reg m_in_15_1_lpi_1_dfm_1_4;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_4;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_4;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_13_cse;
  wire return_add_generic_AC_RND_CONV_false_17_and_9_cse;
  wire return_add_generic_AC_RND_CONV_false_17_and_10_cse;
  wire return_add_generic_AC_RND_CONV_false_17_and_11_cse;
  wire return_add_generic_AC_RND_CONV_false_17_and_12_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_31_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_32_cse;
  wire return_extract_26_exception_and_17_cse;
  wire return_extract_26_exception_and_18_cse;
  wire return_extract_26_exception_and_21_cse;
  wire return_extract_26_exception_and_22_cse;
  wire BUTTERFLY_1_else_1_if_and_3_cse;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_4;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_4;
  reg m_in_15_1_lpi_1_dfm_1_5;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_5;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_5;
  wire BUTTERFLY_1_else_2_and_46_cse;
  wire BUTTERFLY_1_else_3_else_and_26_cse;
  wire BUTTERFLY_1_else_3_else_and_27_cse;
  wire BUTTERFLY_1_else_3_else_and_28_cse;
  wire BUTTERFLY_1_else_3_else_and_30_cse;
  wire BUTTERFLY_1_else_3_else_and_24_cse;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_6;
  reg stage_PE_1_index_const_9_1_lpi_2_dfm_5;
  reg stage_PE_1_qr_10_1_lpi_2_dfm_5;
  reg m_in_15_1_lpi_1_dfm_1_6;
  reg t_in_10_0_lpi_1_dfm_1_8;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_7;
  reg stage_PE_1_qr_1_10_1_lpi_2_dfm_6;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_6;
  reg m_in_15_1_lpi_1_dfm_1_7;
  reg reg_stage_PE_1_qr_10_1_lpi_2_dfm_7_0_ftd;
  reg reg_stage_PE_1_qr_10_1_lpi_2_dfm_7_0_ftd_1;
  reg t_in_10_0_lpi_1_dfm_1_7;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_7;
  reg m_in_15_1_lpi_1_dfm_1_8;
  reg t_in_10_0_lpi_1_dfm_1_6;
  wire stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_8;
  reg m_in_15_1_lpi_1_dfm_1_9;
  reg t_in_10_0_lpi_1_dfm_1_5;
  reg m_in_15_1_lpi_1_dfm_1_10;
  reg t_in_10_0_lpi_1_dfm_1_4;
  reg m_in_15_1_lpi_1_dfm_1_11;
  reg stage_PE_1_index_const_14_11_lpi_2_dfm_0;
  reg t_in_10_0_lpi_1_dfm_1_3;
  reg m_in_15_1_lpi_1_dfm_1_12;
  reg stage_PE_1_index_const_14_11_lpi_2_dfm_1;
  reg t_in_10_0_lpi_1_dfm_1_2;
  reg m_in_15_1_lpi_1_dfm_1_14;
  reg m_in_15_1_lpi_1_dfm_1_13;
  reg stage_PE_1_index_const_14_11_lpi_2_dfm_3;
  reg stage_PE_1_index_const_14_11_lpi_2_dfm_2;
  reg t_in_10_0_lpi_1_dfm_1_1;
  reg t_in_10_0_lpi_1_dfm_1_0;
  wire or_dcpl_1189;
  wire or_dcpl_1191;
  wire BUTTERFLY_1_i_or_cse;
  wire BUTTERFLY_else_1_or_cse;
  wire [50:0] return_extract_32_mux_4_cse;
  wire return_add_generic_AC_RND_CONV_false_e_dif_qif_or_cse;
  wire return_add_generic_AC_RND_CONV_false_e_dif_qif_and_1_cse;
  wire nor_204_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_51_itm;
  wire return_add_generic_AC_RND_CONV_false_4_or_53_itm;
  wire return_add_generic_AC_RND_CONV_false_4_or_55_itm;
  wire return_add_generic_AC_RND_CONV_false_4_or_57_itm;
  wire return_mult_generic_AC_RND_CONV_false_exp_or_4_itm;
  wire [5:0] operator_6_false_8_acc_itm;
  wire [6:0] nl_operator_6_false_8_acc_itm;
  wire return_mult_generic_AC_RND_CONV_false_2_if_acc_1_itm_12_1;
  wire return_mult_generic_AC_RND_CONV_false_if_acc_1_itm_12_1;
  wire return_mult_generic_AC_RND_CONV_false_1_if_acc_1_itm_12_1;
  wire return_mult_generic_AC_RND_CONV_false_5_if_acc_1_itm_12_1;
  wire return_mult_generic_AC_RND_CONV_false_3_if_acc_1_itm_12_1;
  wire return_mult_generic_AC_RND_CONV_false_4_if_acc_1_itm_12_1;
  wire return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1;
  wire return_add_generic_AC_RND_CONV_false_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_1_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_9_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_10_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_12_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_13_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_14_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_22_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10_1;
  wire return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1;
  wire return_add_generic_AC_RND_CONV_false_20_acc_3_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_19_acc_3_itm_11_1;
  wire return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1;
  wire [3:0] return_add_generic_AC_RND_CONV_false_5_conc_itm_3_0;
  wire [3:0] return_add_generic_AC_RND_CONV_false_2_conc_68_itm_3_0;
  wire [3:0] return_add_generic_AC_RND_CONV_false_2_conc_69_itm_3_0;
  wire [3:0] return_add_generic_AC_RND_CONV_false_2_conc_70_itm_3_0;
  wire [1:0] BUTTERFLY_i_conc_3_itm_10_9;
  wire [8:0] BUTTERFLY_i_conc_3_itm_8_0;
  wire [5:0] exs_26_itm_5_0;
  wire [6:0] nl_exs_26_itm_5_0;
  wire [5:0] exs_27_itm_5_0;
  wire [6:0] nl_exs_27_itm_5_0;
  wire return_add_generic_AC_RND_CONV_false_2_or_2_seb;
  wire BUTTERFLY_1_nor_1_seb;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_24_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_23_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_30_cse;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_29_cse;
  wire BUTTERFLY_1_else_1_if_and_1_cse;
  wire stage_PE_1_tmp_re_d_or_6_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_3_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_4_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_5_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_6_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_15_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_16_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_13_cse;
  wire return_add_generic_AC_RND_CONV_false_11_and_14_cse;
  wire and_1589_cse;
  wire return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_and_cse;
  wire return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_mux_2_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_112_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_113_cse;
  wire return_add_generic_AC_RND_CONV_false_4_or_116_cse;
  wire return_add_generic_AC_RND_CONV_false_4_and_132_cse;
  wire [15:0] z_out_4_31_16;
  wire return_mult_generic_AC_RND_CONV_false_if_mux_6_ssc;
  wire z_out_31_52;
  wire z_out_32_52;
  wire z_out_33_52;
  wire z_out_34_52;
  wire z_out_35_52;
  wire return_mult_generic_AC_RND_CONV_false_1_if_mux_6_tmp;

  wire[10:0] return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_or_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_6_else_2_else_return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_6_else_2_else_mux_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_acc_nl;
  wire[11:0] nl_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_acc_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl;
  wire BUTTERFLY_if_1_and_nl;
  wire BUTTERFLY_if_1_and_1_nl;
  wire[50:0] return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_oelse_3_not_1_nl;
  wire stage_PE_qif_qelse_or_nl;
  wire stage_PE_qif_qelse_mux_nl;
  wire stage_PE_qif_qelse_mux_1_nl;
  wire stage_PE_qif_qelse_mux_14_nl;
  wire stage_PE_qif_qelse_mux_13_nl;
  wire stage_PE_qif_qelse_mux_12_nl;
  wire stage_PE_qif_qelse_mux_11_nl;
  wire[9:0] BUTTERFLY_fry_BUTTERFLY_fry_mux_nl;
  wire not_709_nl;
  wire return_extract_15_return_extract_15_nor_nl;
  wire return_extract_47_return_extract_47_nor_nl;
  wire return_extract_20_m_zero_return_extract_20_m_zero_nor_nl;
  wire return_extract_25_m_zero_return_extract_25_m_zero_nor_nl;
  wire return_extract_54_m_zero_return_extract_54_m_zero_nor_nl;
  wire operator_11_true_15_operator_11_true_15_and_nl;
  wire operator_11_true_21_operator_11_true_21_and_nl;
  wire operator_11_true_27_operator_11_true_27_and_nl;
  wire operator_11_true_53_operator_11_true_53_and_nl;
  wire operator_11_true_59_operator_11_true_59_and_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_6_nl;
  wire return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_3_nl;
  wire return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_3_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_5_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_8_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_or_10_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_or_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_or_5_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_or_6_nl;
  wire return_extract_15_return_extract_15_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_2_nl;
  wire return_extract_47_return_extract_47_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_17_e_r_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_17_if_2_return_add_generic_AC_RND_CONV_false_17_if_2_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_17_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_17_and_7_nl;
  wire return_add_generic_AC_RND_CONV_false_17_and_8_nl;
  wire return_add_generic_AC_RND_CONV_false_18_if_2_return_add_generic_AC_RND_CONV_false_18_if_2_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_18_r_sign_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_5_do_sub_return_add_generic_AC_RND_CONV_false_5_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_10_do_sub_return_add_generic_AC_RND_CONV_false_10_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_23_do_sub_return_add_generic_AC_RND_CONV_false_23_do_sub_xor_nl;
  wire return_extract_18_and_nl;
  wire return_add_generic_AC_RND_CONV_false_21_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_8_e_dif_sat_or_1_nl;
  wire[5:0] return_add_generic_AC_RND_CONV_false_11_e_dif_sat_or_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_or_10_nl;
  wire reg_return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_rgt_nl;
  wire return_add_generic_AC_RND_CONV_false_1_op_bigger_return_add_generic_AC_RND_CONV_false_13_op2_mu_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_13_op2_mu_or_nl;
  wire return_add_generic_AC_RND_CONV_false_14_op_bigger_return_add_generic_AC_RND_CONV_false_13_op2_mu_nor_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_5_ma1_lt_ma2_acc_2_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_5_ma1_lt_ma2_acc_2_nl;
  wire and_933_nl;
  wire return_extract_22_m_zero_return_extract_22_m_zero_nor_nl;
  wire return_extract_53_m_zero_return_extract_53_m_zero_nor_nl;
  wire return_extract_59_m_zero_return_extract_59_m_zero_nor_nl;
  wire operator_11_true_20_operator_11_true_20_and_nl;
  wire operator_11_true_25_operator_11_true_25_and_nl;
  wire return_add_generic_AC_RND_CONV_false_12_r_nan_and_nl;
  wire operator_11_true_52_operator_11_true_52_and_nl;
  wire operator_11_true_57_operator_11_true_57_and_nl;
  wire return_add_generic_AC_RND_CONV_false_25_r_nan_and_nl;
  wire return_extract_21_m_zero_return_extract_21_m_zero_nor_nl;
  wire return_extract_27_m_zero_return_extract_27_m_zero_nor_nl;
  wire return_extract_17_m_zero_or_2_nl;
  wire return_extract_17_m_zero_mux_nl;
  wire operator_11_true_22_operator_11_true_22_and_nl;
  wire operator_11_true_47_operator_11_true_47_and_nl;
  wire operator_11_true_54_operator_11_true_54_and_nl;
  wire return_extract_17_return_extract_17_or_1_nl;
  wire or_1586_nl;
  wire or_1606_nl;
  wire return_extract_52_m_zero_return_extract_52_m_zero_nor_nl;
  wire return_extract_57_m_zero_return_extract_57_m_zero_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_7_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_8_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_9_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_10_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_11_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_12_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_17_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_18_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_19_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_20_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_21_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_22_nl;
  wire return_add_generic_AC_RND_CONV_false_13_or_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl;
  wire[52:0] return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl;
  wire[53:0] nl_return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl;
  wire return_add_generic_AC_RND_CONV_false_2_if_2_return_add_generic_AC_RND_CONV_false_2_if_2_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_15_if_2_return_add_generic_AC_RND_CONV_false_15_if_2_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_11_or_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_27_nl;
  wire return_add_generic_AC_RND_CONV_false_11_and_35_nl;
  wire return_add_generic_AC_RND_CONV_false_2_do_sub_return_add_generic_AC_RND_CONV_false_2_do_sub_return_add_generic_AC_RND_CONV_false_2_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_15_do_sub_return_add_generic_AC_RND_CONV_false_15_do_sub_return_add_generic_AC_RND_CONV_false_15_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_22_do_sub_return_add_generic_AC_RND_CONV_false_22_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_10_or_3_nl;
  wire return_add_generic_AC_RND_CONV_false_if_2_return_add_generic_AC_RND_CONV_false_if_2_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_1_if_2_return_add_generic_AC_RND_CONV_false_1_if_2_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_13_if_2_return_add_generic_AC_RND_CONV_false_13_if_2_and_2_nl;
  wire return_add_generic_AC_RND_CONV_false_14_if_2_return_add_generic_AC_RND_CONV_false_14_if_2_and_2_nl;
  wire return_extract_26_exception_or_nl;
  wire return_extract_26_exception_or_4_nl;
  wire return_extract_26_exception_and_4_nl;
  wire return_extract_26_exception_or_5_nl;
  wire return_extract_26_exception_and_8_nl;
  wire and_493_nl;
  wire return_extract_26_exception_or_6_nl;
  wire return_extract_26_exception_and_9_nl;
  wire return_add_generic_AC_RND_CONV_false_10_or_4_nl;
  wire and_498_nl;
  wire return_add_generic_AC_RND_CONV_false_10_and_4_nl;
  wire return_add_generic_AC_RND_CONV_false_3_r_nan_and_nl;
  wire return_add_generic_AC_RND_CONV_false_16_r_nan_and_nl;
  wire return_add_generic_AC_RND_CONV_false_24_r_nan_and_nl;
  wire return_extract_58_and_2_nl;
  wire return_extract_58_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_9_do_sub_return_add_generic_AC_RND_CONV_false_9_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_8_do_sub_return_add_generic_AC_RND_CONV_false_8_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_21_do_sub_return_add_generic_AC_RND_CONV_false_21_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_3_if_2_return_add_generic_AC_RND_CONV_false_3_if_2_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_16_if_2_return_add_generic_AC_RND_CONV_false_16_if_2_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_12_or_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_10_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_5_nl;
  wire return_add_generic_AC_RND_CONV_false_12_and_14_nl;
  wire return_add_generic_AC_RND_CONV_false_3_do_sub_return_add_generic_AC_RND_CONV_false_3_do_sub_return_add_generic_AC_RND_CONV_false_3_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_7_do_sub_return_add_generic_AC_RND_CONV_false_7_do_sub_xor_nl;
  wire return_add_generic_AC_RND_CONV_false_16_do_sub_return_add_generic_AC_RND_CONV_false_16_do_sub_return_add_generic_AC_RND_CONV_false_16_do_sub_xnor_nl;
  wire return_add_generic_AC_RND_CONV_false_20_do_sub_return_add_generic_AC_RND_CONV_false_20_do_sub_xor_nl;
  wire return_extract_26_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_2_not_4_nl;
  wire return_extract_26_and_2_nl;
  wire return_extract_56_and_2_nl;
  wire return_extract_56_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_12_op_bigger_or_4_nl;
  wire return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_6_nl;
  wire return_add_generic_AC_RND_CONV_false_12_res_mant_return_add_generic_AC_RND_CONV_false_12_res_mant_return_add_generic_AC_RND_CONV_false_12_res_mant_or_nl;
  wire return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_33_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_and_35_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_1_nl;
  wire[5:0] return_add_generic_AC_RND_CONV_false_25_e_dif_sat_or_nl;
  wire return_add_generic_AC_RND_CONV_false_25_e_dif_sat_or_1_nl;
  wire[12:0] return_mult_generic_AC_RND_CONV_false_2_if_acc_1_nl;
  wire[13:0] nl_return_mult_generic_AC_RND_CONV_false_2_if_acc_1_nl;
  wire[12:0] return_mult_generic_AC_RND_CONV_false_if_acc_1_nl;
  wire[13:0] nl_return_mult_generic_AC_RND_CONV_false_if_acc_1_nl;
  wire[12:0] return_mult_generic_AC_RND_CONV_false_1_if_acc_1_nl;
  wire[13:0] nl_return_mult_generic_AC_RND_CONV_false_1_if_acc_1_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux_29_nl;
  wire[12:0] return_mult_generic_AC_RND_CONV_false_5_if_acc_1_nl;
  wire[13:0] nl_return_mult_generic_AC_RND_CONV_false_5_if_acc_1_nl;
  wire[12:0] return_mult_generic_AC_RND_CONV_false_3_if_acc_1_nl;
  wire[13:0] nl_return_mult_generic_AC_RND_CONV_false_3_if_acc_1_nl;
  wire[12:0] return_mult_generic_AC_RND_CONV_false_4_if_acc_1_nl;
  wire[13:0] nl_return_mult_generic_AC_RND_CONV_false_4_if_acc_1_nl;
  wire[11:0] return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl;
  wire[12:0] nl_return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_4_mux_18_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_1_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux_19_nl;
  wire return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_2_nl;
  wire return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_2_r_nan_or_1_nl;
  wire and_358_nl;
  wire and_366_nl;
  wire return_add_generic_AC_RND_CONV_false_6_mux_6_nl;
  wire return_add_generic_AC_RND_CONV_false_6_r_sign_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_and_nl;
  wire and_367_nl;
  wire and_374_nl;
  wire return_add_generic_AC_RND_CONV_false_19_mux_6_nl;
  wire return_add_generic_AC_RND_CONV_false_19_r_sign_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_and_nl;
  wire return_add_generic_AC_RND_CONV_false_4_if_7_not_5_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_4_acc_2_nl;
  wire[11:0] nl_return_add_generic_AC_RND_CONV_false_4_acc_2_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux_15_nl;
  wire return_add_generic_AC_RND_CONV_false_4_if_5_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_4_e_dif_sat_or_2_nl;
  wire and_411_nl;
  wire and_415_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_17_mux_18_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nand_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nand_1_nl;
  wire return_add_generic_AC_RND_CONV_false_17_mux_19_nl;
  wire return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nand_2_nl;
  wire return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_7_r_sign_mux_1_nl;
  wire nand_108_nl;
  wire return_add_generic_AC_RND_CONV_false_20_r_sign_mux_1_nl;
  wire nand_109_nl;
  wire return_add_generic_AC_RND_CONV_false_2_e_dif_sat_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_oelse_3_return_mult_generic_AC_RND_CONV_false_1_if_3_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_oelse_3_return_mult_generic_AC_RND_CONV_false_3_if_3_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_oelse_3_return_mult_generic_AC_RND_CONV_false_if_3_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_oelse_3_return_mult_generic_AC_RND_CONV_false_4_if_3_nor_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_5_mux_25_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_5_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_7_nl;
  wire return_add_generic_AC_RND_CONV_false_5_mux_23_nl;
  wire return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_3_nl;
  wire return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_5_mux_27_nl;
  wire return_add_generic_AC_RND_CONV_false_5_if_5_or_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_1_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_1_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_9_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_9_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_10_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_10_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_11_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_11_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_12_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_12_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_13_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_13_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_14_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_14_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_22_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_22_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_23_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_23_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_24_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_24_acc_2_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_25_acc_2_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_25_acc_2_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif_sat_or_1_nl;
  wire and_460_nl;
  wire and_464_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_nl;
  wire or_265_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_2_nl;
  wire or_340_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_1_else_2_else_return_mult_generic_AC_RND_CONV_false_1_else_2_else_and_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_1_else_2_else_else_mux_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_3_else_2_else_return_mult_generic_AC_RND_CONV_false_3_else_2_else_and_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_3_else_2_else_else_mux_nl;
  wire[11:0] operator_33_true_1_acc_nl;
  wire[12:0] nl_operator_33_true_1_acc_nl;
  wire return_add_generic_AC_RND_CONV_false_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_1_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_1_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_2_if_7_return_add_generic_AC_RND_CONV_false_2_if_7_nor_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_else_2_else_return_mult_generic_AC_RND_CONV_false_else_2_else_and_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_else_2_else_else_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_2_e_r_qelse_not_5_nl;
  wire return_add_generic_AC_RND_CONV_false_2_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_2_if_5_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_if_not_nl;
  wire return_mult_generic_AC_RND_CONV_false_return_mult_generic_AC_RND_CONV_false_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_not_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_4_else_2_else_return_mult_generic_AC_RND_CONV_false_4_else_2_else_and_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_4_else_2_else_else_mux_nl;
  wire return_add_generic_AC_RND_CONV_false_8_r_sign_mux_1_nl;
  wire nand_114_nl;
  wire return_add_generic_AC_RND_CONV_false_21_r_sign_mux_1_nl;
  wire nand_115_nl;
  wire return_add_generic_AC_RND_CONV_false_15_if_7_return_add_generic_AC_RND_CONV_false_15_if_7_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_3_if_7_return_add_generic_AC_RND_CONV_false_3_if_7_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_3_e_r_return_add_generic_AC_RND_CONV_false_3_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_2_nl;
  wire or_278_nl;
  wire return_add_generic_AC_RND_CONV_false_3_r_nan_or_1_nl;
  wire and_502_nl;
  wire and_510_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_not_7_nl;
  wire return_add_generic_AC_RND_CONV_false_3_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_3_if_5_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_return_mult_generic_AC_RND_CONV_false_1_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_dif_sat_or_1_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_2_else_2_else_return_mult_generic_AC_RND_CONV_false_2_else_2_else_and_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_2_else_2_else_else_mux_nl;
  wire and_514_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_oelse_3_return_mult_generic_AC_RND_CONV_false_2_if_3_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_return_mult_generic_AC_RND_CONV_false_2_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_6_r_nan_or_1_nl;
  wire and_521_nl;
  wire return_add_generic_AC_RND_CONV_false_6_if_7_return_add_generic_AC_RND_CONV_false_6_if_7_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_5_nl;
  wire or_290_nl;
  wire return_add_generic_AC_RND_CONV_false_6_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_6_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_7_nl;
  wire or_299_nl;
  wire return_add_generic_AC_RND_CONV_false_7_r_nan_or_1_nl;
  wire and_529_nl;
  wire return_add_generic_AC_RND_CONV_false_7_if_7_return_add_generic_AC_RND_CONV_false_7_if_7_nor_nl;
  wire return_extract_25_return_extract_25_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_7_mux_18_nl;
  wire return_add_generic_AC_RND_CONV_false_7_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_9_nl;
  wire or_308_nl;
  wire return_add_generic_AC_RND_CONV_false_8_r_nan_or_1_nl;
  wire and_534_nl;
  wire return_add_generic_AC_RND_CONV_false_8_if_7_return_add_generic_AC_RND_CONV_false_8_if_7_nor_nl;
  wire return_extract_27_return_extract_27_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_8_mux_14_nl;
  wire return_add_generic_AC_RND_CONV_false_8_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_9_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_9_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_10_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_10_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_11_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_11_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_12_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_12_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_12_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_13_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_14_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_15_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_18_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_19_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_20_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_21_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_22_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_23_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_24_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_25_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_26_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_27_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_28_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_29_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_30_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_31_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_32_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_33_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_34_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_35_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_36_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_37_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_38_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_39_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_40_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_41_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_42_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_43_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_44_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_45_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_46_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_47_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_48_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_49_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_50_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_51_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_52_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_53_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_54_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_55_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_56_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_57_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_58_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_59_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_60_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_61_nl;
  wire return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_62_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_17_acc_2_nl;
  wire[11:0] nl_return_add_generic_AC_RND_CONV_false_17_acc_2_nl;
  wire return_add_generic_AC_RND_CONV_false_17_mux_15_nl;
  wire return_add_generic_AC_RND_CONV_false_17_if_5_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_13_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_13_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_14_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_14_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_15_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_15_if_5_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_return_mult_generic_AC_RND_CONV_false_3_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_mux_1_nl;
  wire return_add_generic_AC_RND_CONV_false_16_if_7_return_add_generic_AC_RND_CONV_false_16_if_7_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_16_e_r_return_add_generic_AC_RND_CONV_false_16_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_13_nl;
  wire or_351_nl;
  wire return_add_generic_AC_RND_CONV_false_16_r_nan_or_1_nl;
  wire and_535_nl;
  wire and_542_nl;
  wire return_add_generic_AC_RND_CONV_false_16_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_16_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_smaller_mux_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_return_mult_generic_AC_RND_CONV_false_4_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_mux_1_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_5_else_2_else_return_mult_generic_AC_RND_CONV_false_5_else_2_else_and_nl;
  wire[10:0] return_mult_generic_AC_RND_CONV_false_5_else_2_else_else_mux_nl;
  wire and_546_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_oelse_3_return_mult_generic_AC_RND_CONV_false_5_if_3_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_return_mult_generic_AC_RND_CONV_false_5_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_mux_1_nl;
  wire and_551_nl;
  wire return_add_generic_AC_RND_CONV_false_19_if_7_return_add_generic_AC_RND_CONV_false_19_if_7_nor_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_15_nl;
  wire or_358_nl;
  wire return_add_generic_AC_RND_CONV_false_19_mux_16_nl;
  wire return_add_generic_AC_RND_CONV_false_19_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_17_nl;
  wire or_364_nl;
  wire return_add_generic_AC_RND_CONV_false_20_r_nan_or_1_nl;
  wire and_554_nl;
  wire return_add_generic_AC_RND_CONV_false_20_if_7_return_add_generic_AC_RND_CONV_false_20_if_7_nor_nl;
  wire return_extract_57_return_extract_57_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_20_mux_18_nl;
  wire return_add_generic_AC_RND_CONV_false_20_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_19_nl;
  wire or_368_nl;
  wire return_add_generic_AC_RND_CONV_false_21_r_nan_or_1_nl;
  wire and_557_nl;
  wire return_add_generic_AC_RND_CONV_false_21_if_7_return_add_generic_AC_RND_CONV_false_21_if_7_nor_nl;
  wire return_extract_59_return_extract_59_or_2_nl;
  wire return_add_generic_AC_RND_CONV_false_23_e_dif_sat_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_21_mux_14_nl;
  wire return_add_generic_AC_RND_CONV_false_21_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_22_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_22_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_23_mux_17_nl;
  wire return_add_generic_AC_RND_CONV_false_23_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_24_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_24_if_5_or_nl;
  wire return_add_generic_AC_RND_CONV_false_25_mux_10_nl;
  wire return_add_generic_AC_RND_CONV_false_25_if_5_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_if_if_not_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_mux_1_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_18_acc_3_nl;
  wire[11:0] nl_return_add_generic_AC_RND_CONV_false_18_acc_3_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_20_acc_3_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_20_acc_3_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_8_acc_3_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_8_acc_3_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_19_acc_3_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_19_acc_3_nl;
  wire[11:0] return_add_generic_AC_RND_CONV_false_15_acc_3_nl;
  wire[12:0] nl_return_add_generic_AC_RND_CONV_false_15_acc_3_nl;
  wire BUTTERFLY_1_i_mux1h_1_nl;
  wire[8:0] mux1h_6_nl;
  wire or_2472_nl;
  wire or_2473_nl;
  wire BUTTERFLY_if_1_if_mux1h_nl;
  wire BUTTERFLY_if_1_if_or_nl;
  wire[9:0] or_2035_nl;
  wire[9:0] and_2431_nl;
  wire[9:0] mux1h_nl;
  wire and_2423_nl;
  wire and_2424_nl;
  wire and_2425_nl;
  wire and_2426_nl;
  wire or_2461_nl;
  wire not_760_nl;
  wire BUTTERFLY_if_1_if_mux1h_2_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_return_add_generic_AC_RND_CONV_false_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_nl;
  wire or_245_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_r_return_add_generic_AC_RND_CONV_false_1_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_14_e_r_qelse_mux_nl;
  wire or_257_nl;
  wire return_add_generic_AC_RND_CONV_false_9_e_r_return_add_generic_AC_RND_CONV_false_9_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_nl;
  wire or_375_nl;
  wire return_add_generic_AC_RND_CONV_false_10_e_r_return_add_generic_AC_RND_CONV_false_10_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_21_nl;
  wire or_386_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_return_add_generic_AC_RND_CONV_false_11_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_5_nl;
  wire or_397_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_r_return_add_generic_AC_RND_CONV_false_12_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_3_nl;
  wire or_407_nl;
  wire BUTTERFLY_if_1_if_mux1h_3_nl;
  wire return_add_generic_AC_RND_CONV_false_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_9_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_10_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_11_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_12_r_nan_or_nl;
  wire BUTTERFLY_if_1_if_or_2_nl;
  wire BUTTERFLY_if_1_if_and_7_nl;
  wire[50:0] nor_182_nl;
  wire[50:0] nor_183_nl;
  wire[50:0] mux1h_1_nl;
  wire and_2433_nl;
  wire and_2434_nl;
  wire and_2435_nl;
  wire and_2432_nl;
  wire or_1217_nl;
  wire or_1218_nl;
  wire[1:0] mux1h_7_nl;
  wire[2:0] mux1h_8_nl;
  wire mux1h_12_nl;
  wire[4:0] mux1h_13_nl;
  wire[4:0] mux1h_14_nl;
  wire BUTTERFLY_if_1_mux1h_2_nl;
  wire[8:0] mux1h_9_nl;
  wire or_2474_nl;
  wire or_2475_nl;
  wire BUTTERFLY_if_1_mux1h_1_nl;
  wire BUTTERFLY_if_1_or_nl;
  wire[9:0] or_2036_nl;
  wire[9:0] and_2449_nl;
  wire[9:0] mux1h_2_nl;
  wire and_2441_nl;
  wire and_2442_nl;
  wire and_2443_nl;
  wire and_2444_nl;
  wire or_2460_nl;
  wire not_763_nl;
  wire BUTTERFLY_if_1_mux1h_6_nl;
  wire return_add_generic_AC_RND_CONV_false_13_e_r_return_add_generic_AC_RND_CONV_false_13_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_11_nl;
  wire or_320_nl;
  wire return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_14_e_r_qelse_mux_3_nl;
  wire or_332_nl;
  wire return_add_generic_AC_RND_CONV_false_22_e_r_return_add_generic_AC_RND_CONV_false_22_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_7_nl;
  wire or_417_nl;
  wire return_add_generic_AC_RND_CONV_false_23_e_r_return_add_generic_AC_RND_CONV_false_23_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_23_nl;
  wire or_429_nl;
  wire return_add_generic_AC_RND_CONV_false_24_e_r_return_add_generic_AC_RND_CONV_false_24_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_5_nl;
  wire or_439_nl;
  wire return_add_generic_AC_RND_CONV_false_25_e_r_return_add_generic_AC_RND_CONV_false_25_e_r_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_9_nl;
  wire or_449_nl;
  wire BUTTERFLY_if_1_mux1h_7_nl;
  wire return_add_generic_AC_RND_CONV_false_13_r_nan_or_1_nl;
  wire return_add_generic_AC_RND_CONV_false_22_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_23_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_24_r_nan_or_nl;
  wire return_add_generic_AC_RND_CONV_false_25_r_nan_or_nl;
  wire BUTTERFLY_if_1_or_2_nl;
  wire BUTTERFLY_if_1_and_9_nl;
  wire[50:0] nor_186_nl;
  wire[50:0] nor_187_nl;
  wire[50:0] mux1h_3_nl;
  wire and_2451_nl;
  wire and_2452_nl;
  wire and_2453_nl;
  wire and_2450_nl;
  wire or_1191_nl;
  wire or_1192_nl;
  wire[1:0] mux1h_10_nl;
  wire[2:0] mux1h_11_nl;
  wire mux1h_15_nl;
  wire[4:0] mux1h_16_nl;
  wire[4:0] mux1h_17_nl;
  wire return_add_generic_AC_RND_CONV_false_e_r_qelse_not_5_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_r_qelse_not_3_nl;
  wire[8:0] BUTTERFLY_n_and_nl;
  wire[8:0] BUTTERFLY_n_mux1h_1_nl;
  wire BUTTERFLY_1_fiy_nand_nl;
  wire or_1355_nl;
  wire or_1996_nl;
  wire or_1998_nl;
  wire or_2005_nl;
  wire or_2010_nl;
  wire stage_PE_1_tmp_im_d_or_1_nl;
  wire stage_PE_1_tmp_re_d_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_op1_normal_not_5_nl;
  wire[12:0] acc_1_nl;
  wire[13:0] nl_acc_1_nl;
  wire operator_6_false_1_mux1h_9_nl;
  wire operator_6_false_1_mux1h_10_nl;
  wire[2:0] operator_6_false_1_mux1h_11_nl;
  wire operator_6_false_1_mux1h_12_nl;
  wire[2:0] operator_6_false_1_mux1h_13_nl;
  wire operator_6_false_1_mux1h_14_nl;
  wire operator_6_false_1_mux1h_15_nl;
  wire operator_6_false_1_or_16_nl;
  wire operator_6_false_1_or_17_nl;
  wire operator_6_false_1_or_18_nl;
  wire[5:0] operator_6_false_1_mux1h_16_nl;
  wire operator_6_false_1_or_19_nl;
  wire operator_6_false_1_or_20_nl;
  wire operator_6_false_1_or_21_nl;
  wire BUTTERFLY_fry_mux_10_nl;
  wire BUTTERFLY_fry_mux_11_nl;
  wire BUTTERFLY_fry_mux_12_nl;
  wire BUTTERFLY_fry_mux_13_nl;
  wire BUTTERFLY_fry_mux_14_nl;
  wire BUTTERFLY_fry_mux_15_nl;
  wire BUTTERFLY_fry_mux_16_nl;
  wire BUTTERFLY_fry_mux_17_nl;
  wire BUTTERFLY_fry_mux_18_nl;
  wire BUTTERFLY_fry_mux_19_nl;
  wire[31:0] operator_32_false_acc_nl;
  wire[34:0] nl_operator_32_false_acc_nl;
  wire return_add_generic_AC_RND_CONV_false_4_res_rounded_return_add_generic_AC_RND_CONV_false_4_res_rounded_and_1_nl;
  wire[51:0] return_add_generic_AC_RND_CONV_false_4_res_rounded_mux1h_2_nl;
  wire return_add_generic_AC_RND_CONV_false_4_res_rounded_mux1h_3_nl;
  wire return_add_generic_AC_RND_CONV_false_4_res_rounded_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_mux_14_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_1_or_4_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_mux_14_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_1_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_mux_14_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_if_1_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_mux_14_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_if_1_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_mux_14_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_if_1_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_mux_14_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_if_1_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_and_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_mux_12_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_if_1_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_or_1_nl;
  wire BUTTERFLY_if_mux_14_nl;
  wire stage_PE_stage_PE_stage_PE_mux_3_nl;
  wire BUTTERFLY_if_mux_15_nl;
  wire BUTTERFLY_if_mux_16_nl;
  wire BUTTERFLY_if_mux_17_nl;
  wire BUTTERFLY_if_mux_18_nl;
  wire BUTTERFLY_if_mux_19_nl;
  wire BUTTERFLY_if_mux_20_nl;
  wire BUTTERFLY_if_mux_21_nl;
  wire BUTTERFLY_if_mux_22_nl;
  wire BUTTERFLY_if_mux_23_nl;
  wire operator_6_false_mux1h_9_nl;
  wire operator_6_false_mux1h_10_nl;
  wire[2:0] operator_6_false_mux1h_11_nl;
  wire operator_6_false_mux1h_12_nl;
  wire[2:0] operator_6_false_mux1h_13_nl;
  wire operator_6_false_mux1h_14_nl;
  wire operator_6_false_mux1h_15_nl;
  wire operator_6_false_or_23_nl;
  wire[5:0] operator_6_false_mux1h_16_nl;
  wire[5:0] operator_6_false_acc_1_nl;
  wire[6:0] nl_operator_6_false_acc_1_nl;
  wire[5:0] operator_6_false_2_acc_1_nl;
  wire[6:0] nl_operator_6_false_2_acc_1_nl;
  wire[5:0] operator_6_false_4_acc_3_nl;
  wire[6:0] nl_operator_6_false_4_acc_3_nl;
  wire[5:0] operator_6_false_23_acc_3_nl;
  wire[6:0] nl_operator_6_false_23_acc_3_nl;
  wire[5:0] operator_6_false_17_acc_3_nl;
  wire[6:0] nl_operator_6_false_17_acc_3_nl;
  wire[5:0] operator_6_false_21_acc_3_nl;
  wire[6:0] nl_operator_6_false_21_acc_3_nl;
  wire[5:0] operator_6_false_29_acc_1_nl;
  wire[6:0] nl_operator_6_false_29_acc_1_nl;
  wire[5:0] operator_6_false_31_acc_1_nl;
  wire[6:0] nl_operator_6_false_31_acc_1_nl;
  wire operator_6_false_mux1h_17_nl;
  wire operator_6_false_or_24_nl;
  wire BUTTERFLY_1_and_2_nl;
  wire BUTTERFLY_1_mux_1_nl;
  wire[4:0] BUTTERFLY_1_and_3_nl;
  wire[4:0] BUTTERFLY_1_mux1h_5_nl;
  wire[3:0] BUTTERFLY_1_mux1h_6_nl;
  wire[1:0] BUTTERFLY_1_BUTTERFLY_1_and_2_nl;
  wire BUTTERFLY_1_nor_2_nl;
  wire BUTTERFLY_i_and_14_nl;
  wire BUTTERFLY_i_mux1h_24_nl;
  wire BUTTERFLY_i_and_15_nl;
  wire BUTTERFLY_i_mux1h_25_nl;
  wire[36:0] BUTTERFLY_i_and_16_nl;
  wire[36:0] BUTTERFLY_i_mux1h_26_nl;
  wire[2:0] BUTTERFLY_i_and_17_nl;
  wire[2:0] BUTTERFLY_i_mux1h_27_nl;
  wire not_815_nl;
  wire BUTTERFLY_i_and_18_nl;
  wire BUTTERFLY_i_mux1h_28_nl;
  wire[4:0] BUTTERFLY_i_mux1h_29_nl;
  wire[4:0] BUTTERFLY_i_mux1h_30_nl;
  wire BUTTERFLY_i_BUTTERFLY_i_and_1_nl;
  wire BUTTERFLY_i_and_19_nl;
  wire BUTTERFLY_i_mux1h_31_nl;
  wire BUTTERFLY_i_and_20_nl;
  wire BUTTERFLY_i_mux1h_32_nl;
  wire BUTTERFLY_i_and_21_nl;
  wire BUTTERFLY_i_mux1h_33_nl;
  wire[32:0] BUTTERFLY_i_and_22_nl;
  wire[32:0] BUTTERFLY_i_mux1h_34_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_not_10_nl;
  wire BUTTERFLY_i_and_23_nl;
  wire BUTTERFLY_i_mux1h_35_nl;
  wire[4:0] BUTTERFLY_i_and_24_nl;
  wire[4:0] BUTTERFLY_i_mux1h_36_nl;
  wire BUTTERFLY_i_and_25_nl;
  wire BUTTERFLY_i_and_26_nl;
  wire return_add_generic_AC_RND_CONV_false_11_op_bigger_not_12_nl;
  wire BUTTERFLY_i_and_27_nl;
  wire BUTTERFLY_i_mux1h_37_nl;
  wire BUTTERFLY_i_mux1h_38_nl;
  wire BUTTERFLY_i_mux1h_39_nl;
  wire BUTTERFLY_i_mux1h_40_nl;
  wire BUTTERFLY_i_mux1h_41_nl;
  wire BUTTERFLY_i_mux1h_42_nl;
  wire BUTTERFLY_i_mux1h_43_nl;
  wire BUTTERFLY_i_mux1h_44_nl;
  wire BUTTERFLY_i_mux1h_45_nl;
  wire BUTTERFLY_i_mux1h_46_nl;
  wire BUTTERFLY_i_mux1h_47_nl;
  wire[12:0] acc_12_nl;
  wire[13:0] nl_acc_12_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif_qif_and_7_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_10_nl;
  wire[4:0] return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_11_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_12_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_13_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif_qif_nor_1_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_14_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif_qif_return_add_generic_AC_RND_CONV_false_e_dif_qif_nor_2_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_15_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_e_dif_qif_return_add_generic_AC_RND_CONV_false_e_dif_qif_nor_3_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_16_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_17_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_18_nl;
  wire[12:0] acc_13_nl;
  wire[13:0] nl_acc_13_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_10_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_11_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_12_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_13_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_14_nl;
  wire[1:0] return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_15_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_16_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_17_nl;
  wire return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_18_nl;
  wire[12:0] acc_14_nl;
  wire[13:0] nl_acc_14_nl;
  wire[1:0] return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_10_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_11_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_12_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_13_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_return_add_generic_AC_RND_CONV_false_1_e_dif1_nand_2_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_14_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_nor_3_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_15_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_1_e_dif1_nor_4_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_16_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_1_e_dif1_nor_5_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_17_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_return_add_generic_AC_RND_CONV_false_1_e_dif1_nand_3_nl;
  wire return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_18_nl;
  wire[12:0] acc_15_nl;
  wire[13:0] nl_acc_15_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_8_e_dif1_mux_4_nl;
  wire[13:0] acc_16_nl;
  wire[14:0] nl_acc_16_nl;
  wire return_mult_generic_AC_RND_CONV_false_exp_return_mult_generic_AC_RND_CONV_false_exp_and_1_nl;
  wire[5:0] return_mult_generic_AC_RND_CONV_false_exp_mux1h_12_nl;
  wire[3:0] return_mult_generic_AC_RND_CONV_false_exp_mux1h_13_nl;
  wire return_mult_generic_AC_RND_CONV_false_exp_mux1h_14_nl;
  wire return_mult_generic_AC_RND_CONV_false_exp_or_12_nl;
  wire return_mult_generic_AC_RND_CONV_false_exp_mux1h_15_nl;
  wire[1:0] return_mult_generic_AC_RND_CONV_false_exp_return_mult_generic_AC_RND_CONV_false_exp_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_exp_or_13_nl;
  wire[8:0] return_mult_generic_AC_RND_CONV_false_exp_mux1h_16_nl;
  wire return_mult_generic_AC_RND_CONV_false_exp_mux1h_17_nl;
  wire[11:0] acc_17_nl;
  wire[12:0] nl_acc_17_nl;
  wire operator_6_false_9_mux_4_nl;
  wire[3:0] operator_6_false_9_mux_5_nl;
  wire[3:0] operator_6_false_9_mux_6_nl;
  wire operator_6_false_9_mux_7_nl;
  wire[13:0] acc_18_nl;
  wire[14:0] nl_acc_18_nl;
  wire operator_6_false_14_operator_6_false_14_mux_2_nl;
  wire[57:0] acc_19_nl;
  wire[58:0] nl_acc_19_nl;
  wire[44:0] return_add_generic_AC_RND_CONV_false_4_mux1h_25_nl;
  wire[10:0] return_add_generic_AC_RND_CONV_false_4_mux1h_26_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux1h_27_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_137_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_138_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_139_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_140_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_117_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_141_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_142_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_143_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_144_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_145_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_146_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_147_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_148_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_149_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_150_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_151_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_152_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_153_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_154_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_155_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_156_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_157_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux1h_28_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_158_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux1h_29_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_121_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_122_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_123_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_159_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux1h_30_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_124_nl;
  wire[29:0] return_add_generic_AC_RND_CONV_false_4_and_160_nl;
  wire[29:0] return_add_generic_AC_RND_CONV_false_4_mux1h_31_nl;
  wire return_add_generic_AC_RND_CONV_false_4_not_59_nl;
  wire[9:0] return_add_generic_AC_RND_CONV_false_4_mux1h_32_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_4_and_161_nl;
  wire[3:0] return_add_generic_AC_RND_CONV_false_4_mux1h_33_nl;
  wire return_add_generic_AC_RND_CONV_false_4_not_60_nl;
  wire[5:0] return_add_generic_AC_RND_CONV_false_4_mux1h_34_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux1h_35_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_125_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_126_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_127_nl;
  wire[2:0] return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_8_nl;
  wire return_add_generic_AC_RND_CONV_false_4_nor_1_nl;
  wire[53:0] acc_20_nl;
  wire[54:0] nl_acc_20_nl;
  wire[53:0] acc_21_nl;
  wire[54:0] nl_acc_21_nl;
  wire return_add_generic_AC_RND_CONV_false_6_ma1_lt_ma2_mux_5_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_6_ma1_lt_ma2_mux_6_nl;
  wire[53:0] acc_22_nl;
  wire[54:0] nl_acc_22_nl;
  wire return_add_generic_AC_RND_CONV_false_9_ma1_lt_ma2_mux_4_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_9_ma1_lt_ma2_mux_5_nl;
  wire[53:0] acc_23_nl;
  wire[54:0] nl_acc_23_nl;
  wire return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_mux1h_4_nl;
  wire[50:0] return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_mux1h_5_nl;
  wire[53:0] acc_24_nl;
  wire[54:0] nl_acc_24_nl;
  wire[18:0] acc_26_nl;
  wire[19:0] nl_acc_26_nl;
  wire[5:0] operator_6_false_8_mux1h_12_nl;
  wire operator_6_false_8_mux1h_13_nl;
  wire operator_6_false_8_mux1h_14_nl;
  wire[3:0] operator_6_false_8_mux1h_15_nl;
  wire[3:0] operator_6_false_8_mux1h_16_nl;
  wire operator_6_false_8_mux1h_17_nl;
  wire operator_6_false_8_or_3_nl;
  wire operator_6_false_8_or_4_nl;
  wire[4:0] operator_6_false_8_and_2_nl;
  wire[4:0] operator_6_false_8_mux1h_18_nl;
  wire operator_6_false_8_and_3_nl;
  wire operator_6_false_8_mux1h_19_nl;
  wire operator_6_false_8_mux1h_20_nl;
  wire[3:0] operator_6_false_8_mux1h_21_nl;
  wire[3:0] operator_6_false_8_mux1h_22_nl;
  wire operator_6_false_8_mux1h_23_nl;
  wire[15:0] BUTTERFLY_1_else_1_if_BUTTERFLY_1_else_1_if_mux_4_nl;
  wire[12:0] acc_28_nl;
  wire[13:0] nl_acc_28_nl;
  wire[9:0] return_mult_generic_AC_RND_CONV_false_exp_return_mult_generic_AC_RND_CONV_false_exp_mux_4_nl;
  wire return_mult_generic_AC_RND_CONV_false_exp_return_mult_generic_AC_RND_CONV_false_exp_mux_5_nl;
  wire return_mult_generic_AC_RND_CONV_false_exp_mux1h_18_nl;
  wire[17:0] acc_29_nl;
  wire[18:0] nl_acc_29_nl;
  wire[15:0] stage_u_add_mux1h_8_nl;
  wire stage_u_add_or_4_nl;
  wire stage_u_add_or_5_nl;
  wire[1:0] stage_u_add_mux1h_9_nl;
  wire[2:0] stage_u_add_mux1h_10_nl;
  wire stage_u_add_mux1h_11_nl;
  wire stage_u_add_mux1h_12_nl;
  wire[3:0] stage_u_add_mux1h_13_nl;
  wire[4:0] stage_u_add_mux1h_14_nl;
  wire[12:0] acc_31_nl;
  wire[13:0] nl_acc_31_nl;
  wire[9:0] return_mult_generic_AC_RND_CONV_false_2_exp_mux_3_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_exp_mux_4_nl;
  wire[5:0] BUTTERFLY_else_2_mux_14_nl;
  wire BUTTERFLY_else_2_mux_15_nl;
  wire BUTTERFLY_else_2_mux_16_nl;
  wire[3:0] BUTTERFLY_else_2_mux_17_nl;
  wire[3:0] BUTTERFLY_else_2_mux_18_nl;
  wire BUTTERFLY_else_2_mux_19_nl;
  wire[2:0] BUTTERFLY_else_2_BUTTERFLY_else_2_and_6_nl;
  wire[1:0] BUTTERFLY_else_2_mux_20_nl;
  wire BUTTERFLY_else_2_BUTTERFLY_else_2_and_7_nl;
  wire BUTTERFLY_else_2_BUTTERFLY_else_2_and_8_nl;
  wire BUTTERFLY_else_2_BUTTERFLY_else_2_and_9_nl;
  wire[3:0] BUTTERFLY_else_2_BUTTERFLY_else_2_and_10_nl;
  wire[3:0] BUTTERFLY_else_2_BUTTERFLY_else_2_and_11_nl;
  wire BUTTERFLY_else_2_mux_21_nl;
  wire return_add_generic_AC_RND_CONV_false_mux_36_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[5:0] return_add_generic_AC_RND_CONV_false_4_mux1h_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux1h_15_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_4_mux1h_8_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_a;
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_nl = MUX1HOT_v_6_4_2((z_out_30[56:51]),
      (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[56:51]), stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_0,
      (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_56_50[6:1]), {return_add_generic_AC_RND_CONV_false_4_or_20_ssc
      , return_add_generic_AC_RND_CONV_false_4_or_18_ssc , return_add_generic_AC_RND_CONV_false_4_or_ssc
      , or_dcpl_397});
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_15_nl = MUX1HOT_s_1_4_2((z_out_30[50]),
      (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[50]), (stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_1[50]),
      (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_56_50[0]), {return_add_generic_AC_RND_CONV_false_4_or_20_ssc
      , return_add_generic_AC_RND_CONV_false_4_or_18_ssc , return_add_generic_AC_RND_CONV_false_4_or_ssc
      , or_dcpl_397});
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_8_nl = MUX1HOT_v_50_4_2((z_out_30[49:0]),
      (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[49:0]), (stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_1[49:0]),
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_49_0, {return_add_generic_AC_RND_CONV_false_4_or_20_ssc
      , return_add_generic_AC_RND_CONV_false_4_or_18_ssc , return_add_generic_AC_RND_CONV_false_4_or_ssc
      , or_dcpl_397});
  assign nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_a = {return_add_generic_AC_RND_CONV_false_4_mux1h_nl
      , return_add_generic_AC_RND_CONV_false_4_mux1h_15_nl , return_add_generic_AC_RND_CONV_false_4_mux1h_8_nl};
  wire return_add_generic_AC_RND_CONV_false_4_mux1h_1_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_123_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_114_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_125_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_115_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_129_nl;
  wire return_add_generic_AC_RND_CONV_false_4_and_135_nl;
  wire[2:0] return_add_generic_AC_RND_CONV_false_4_mux1h_23_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux1h_24_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux1h_9_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_110_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_58_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_60_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_62_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_64_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_s;
  assign return_add_generic_AC_RND_CONV_false_4_and_123_nl = (~ return_add_generic_AC_RND_CONV_false_acc_2_itm_11_1)
      & (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_4_or_114_nl = (return_add_generic_AC_RND_CONV_false_acc_2_itm_11_1
      & (fsm_output[5])) | (return_add_generic_AC_RND_CONV_false_13_acc_2_itm_11_1
      & (fsm_output[30]));
  assign return_add_generic_AC_RND_CONV_false_4_and_125_nl = (~ return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva)
      & return_extract_26_exception_or_3_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_115_nl = (return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva
      & return_extract_26_exception_or_3_cse) | (return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1
      & or_tmp_983) | return_add_generic_AC_RND_CONV_false_4_and_132_cse | return_add_generic_AC_RND_CONV_false_4_or_54_cse;
  assign return_add_generic_AC_RND_CONV_false_4_and_129_nl = (~ return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1)
      & or_tmp_983;
  assign return_add_generic_AC_RND_CONV_false_4_and_135_nl = (~ return_add_generic_AC_RND_CONV_false_13_acc_2_itm_11_1)
      & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_1_nl = MUX1HOT_s_1_16_2((return_add_generic_AC_RND_CONV_false_4_mux_10_itm[5]),
      (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1[0]), (rtn_out[5]), (drf_qr_lval_smx_lpi_3_dfm_mx0_10_5[0]),
      (rtn_out[5]), (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[0]), (return_add_generic_AC_RND_CONV_false_10_ls_sva[5]),
      (return_add_generic_AC_RND_CONV_false_11_ls_sva[5]), (drf_qr_lval_11_smx_lpi_3_dfm_8_5[0]),
      (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2[3]), (return_add_generic_AC_RND_CONV_false_12_ls_sva[5]),
      (drf_qr_lval_13_smx_10_1_lpi_3_dfm[4]), (drf_qr_lval_14_smx_10_1_lpi_3_dfm[4]),
      (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[4]), (return_add_generic_AC_RND_CONV_false_17_mux_10_itm[5]),
      (drf_qr_lval_16_smx_lpi_3_dfm_mx0_10_5[0]), {(fsm_output[3]) , return_add_generic_AC_RND_CONV_false_4_or_112_cse
      , return_add_generic_AC_RND_CONV_false_4_or_113_cse , return_add_generic_AC_RND_CONV_false_4_and_123_nl
      , return_add_generic_AC_RND_CONV_false_4_or_114_nl , return_add_generic_AC_RND_CONV_false_4_and_125_nl
      , return_add_generic_AC_RND_CONV_false_4_or_115_nl , return_add_generic_AC_RND_CONV_false_4_or_116_cse
      , return_add_generic_AC_RND_CONV_false_4_and_129_nl , return_add_generic_AC_RND_CONV_false_4_or_51_itm
      , return_add_generic_AC_RND_CONV_false_4_or_52_cse , return_add_generic_AC_RND_CONV_false_4_or_53_itm
      , return_add_generic_AC_RND_CONV_false_4_or_55_itm , return_add_generic_AC_RND_CONV_false_4_or_57_itm
      , (fsm_output[28]) , return_add_generic_AC_RND_CONV_false_4_and_135_nl});
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_23_nl = MUX1HOT_v_3_17_2((return_add_generic_AC_RND_CONV_false_4_mux_10_itm[4:2]),
      (return_add_generic_AC_RND_CONV_false_5_conc_itm_3_0[3:1]), (return_add_generic_AC_RND_CONV_false_mux_26_itm_4_0[4:2]),
      (return_add_generic_AC_RND_CONV_false_1_mux_25_itm_4_0[4:2]), (return_add_generic_AC_RND_CONV_false_2_conc_68_itm_3_0[3:1]),
      (return_add_generic_AC_RND_CONV_false_3_mux_16_mx0_4_0[4:2]), (return_add_generic_AC_RND_CONV_false_2_conc_69_itm_3_0[3:1]),
      (return_add_generic_AC_RND_CONV_false_2_conc_70_itm_3_0[3:1]), (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2[2:0]),
      (return_add_generic_AC_RND_CONV_false_12_ls_sva[4:2]), (drf_qr_lval_13_smx_10_1_lpi_3_dfm[3:1]),
      (return_add_generic_AC_RND_CONV_false_10_ls_sva[4:2]), (drf_qr_lval_14_smx_10_1_lpi_3_dfm[3:1]),
      (return_add_generic_AC_RND_CONV_false_11_ls_sva[4:2]), (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[3:1]),
      (return_add_generic_AC_RND_CONV_false_17_mux_10_itm[4:2]), (return_add_generic_AC_RND_CONV_false_13_mux_28_itm_4_0[4:2]),
      {(fsm_output[3]) , or_38_cse , (fsm_output[5]) , return_extract_26_exception_or_3_cse
      , or_dcpl_780 , or_tmp_983 , or_dcpl_423 , return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
      , return_add_generic_AC_RND_CONV_false_4_or_51_itm , return_add_generic_AC_RND_CONV_false_4_or_52_cse
      , return_add_generic_AC_RND_CONV_false_4_or_53_itm , return_add_generic_AC_RND_CONV_false_4_or_54_cse
      , return_add_generic_AC_RND_CONV_false_4_or_55_itm , return_add_generic_AC_RND_CONV_false_4_or_56_cse
      , return_add_generic_AC_RND_CONV_false_4_or_57_itm , (fsm_output[28]) , (fsm_output[30])});
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_24_nl = MUX1HOT_s_1_17_2((return_add_generic_AC_RND_CONV_false_4_mux_10_itm[1]),
      (return_add_generic_AC_RND_CONV_false_5_conc_itm_3_0[0]), (return_add_generic_AC_RND_CONV_false_mux_26_itm_4_0[1]),
      (return_add_generic_AC_RND_CONV_false_1_mux_25_itm_4_0[1]), (return_add_generic_AC_RND_CONV_false_2_conc_68_itm_3_0[0]),
      (return_add_generic_AC_RND_CONV_false_3_mux_16_mx0_4_0[1]), (return_add_generic_AC_RND_CONV_false_2_conc_69_itm_3_0[0]),
      (return_add_generic_AC_RND_CONV_false_2_conc_70_itm_3_0[0]), reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3,
      (return_add_generic_AC_RND_CONV_false_12_ls_sva[1]), (drf_qr_lval_13_smx_10_1_lpi_3_dfm[0]),
      (return_add_generic_AC_RND_CONV_false_10_ls_sva[1]), (drf_qr_lval_14_smx_10_1_lpi_3_dfm[0]),
      (return_add_generic_AC_RND_CONV_false_11_ls_sva[1]), (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[0]),
      (return_add_generic_AC_RND_CONV_false_17_mux_10_itm[1]), (return_add_generic_AC_RND_CONV_false_13_mux_28_itm_4_0[1]),
      {(fsm_output[3]) , or_38_cse , (fsm_output[5]) , return_extract_26_exception_or_3_cse
      , or_dcpl_780 , or_tmp_983 , or_dcpl_423 , return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
      , return_add_generic_AC_RND_CONV_false_4_or_51_itm , return_add_generic_AC_RND_CONV_false_4_or_52_cse
      , return_add_generic_AC_RND_CONV_false_4_or_53_itm , return_add_generic_AC_RND_CONV_false_4_or_54_cse
      , return_add_generic_AC_RND_CONV_false_4_or_55_itm , return_add_generic_AC_RND_CONV_false_4_or_56_cse
      , return_add_generic_AC_RND_CONV_false_4_or_57_itm , (fsm_output[28]) , (fsm_output[30])});
  assign return_add_generic_AC_RND_CONV_false_4_or_110_nl = return_add_generic_AC_RND_CONV_false_4_and_132_cse
      | return_add_generic_AC_RND_CONV_false_4_or_54_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_58_nl = return_add_generic_AC_RND_CONV_false_4_and_5_cse
      | return_add_generic_AC_RND_CONV_false_4_and_13_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_60_nl = return_add_generic_AC_RND_CONV_false_4_and_7_cse
      | return_add_generic_AC_RND_CONV_false_4_and_15_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_62_nl = return_add_generic_AC_RND_CONV_false_4_and_9_cse
      | return_add_generic_AC_RND_CONV_false_4_and_17_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_64_nl = return_add_generic_AC_RND_CONV_false_4_and_11_cse
      | return_add_generic_AC_RND_CONV_false_4_and_19_cse;
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_9_nl = MUX1HOT_s_1_15_2((return_add_generic_AC_RND_CONV_false_4_mux_10_itm[0]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3, (rtn_out[0]), (return_add_generic_AC_RND_CONV_false_mux_26_itm_4_0[0]),
      (return_add_generic_AC_RND_CONV_false_1_mux_25_itm_4_0[0]), (return_add_generic_AC_RND_CONV_false_11_ls_sva[0]),
      (return_add_generic_AC_RND_CONV_false_3_mux_16_mx0_4_0[0]), (return_add_generic_AC_RND_CONV_false_10_ls_sva[0]),
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm, (return_add_generic_AC_RND_CONV_false_12_ls_sva[0]),
      drf_qr_lval_13_smx_0_lpi_3_dfm, drf_qr_lval_14_smx_0_lpi_3_dfm, drf_qr_lval_15_smx_0_lpi_3_dfm,
      (return_add_generic_AC_RND_CONV_false_17_mux_10_itm[0]), (return_add_generic_AC_RND_CONV_false_13_mux_28_itm_4_0[0]),
      {(fsm_output[3]) , return_add_generic_AC_RND_CONV_false_4_or_112_cse , return_add_generic_AC_RND_CONV_false_4_or_113_cse
      , (fsm_output[5]) , return_extract_26_exception_or_3_cse , return_add_generic_AC_RND_CONV_false_4_or_116_cse
      , or_tmp_983 , return_add_generic_AC_RND_CONV_false_4_or_110_nl , return_add_generic_AC_RND_CONV_false_4_or_58_nl
      , return_add_generic_AC_RND_CONV_false_4_or_52_cse , return_add_generic_AC_RND_CONV_false_4_or_60_nl
      , return_add_generic_AC_RND_CONV_false_4_or_62_nl , return_add_generic_AC_RND_CONV_false_4_or_64_nl
      , (fsm_output[28]) , (fsm_output[30])});
  assign nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_s = {return_add_generic_AC_RND_CONV_false_4_mux1h_1_nl
      , return_add_generic_AC_RND_CONV_false_4_mux1h_23_nl , return_add_generic_AC_RND_CONV_false_4_mux1h_24_nl
      , return_add_generic_AC_RND_CONV_false_4_mux1h_9_nl};
  wire return_add_generic_AC_RND_CONV_false_4_or_98_nl;
  wire or_2189_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_10_lshift_rg_s;
  assign return_add_generic_AC_RND_CONV_false_4_or_98_nl = (fsm_output[7]) | (fsm_output[14])
      | (fsm_output[18]) | (fsm_output[32]);
  assign or_2189_nl = (fsm_output[4]) | (fsm_output[29]) | (fsm_output[16]) | (fsm_output[41])
      | (fsm_output[42]) | (fsm_output[17]);
  assign nl_return_add_generic_AC_RND_CONV_false_10_lshift_rg_s = MUX1HOT_v_6_8_2(return_add_generic_AC_RND_CONV_false_4_e_dif_sat_sva_1,
      return_add_generic_AC_RND_CONV_false_e_dif_sat_or_cse, return_add_generic_AC_RND_CONV_false_21_e_dif_sat_or_cse,
      return_add_generic_AC_RND_CONV_false_6_e_dif_sat_sva_1, return_add_generic_AC_RND_CONV_false_8_e_dif_sat_or_cse,
      return_add_generic_AC_RND_CONV_false_23_e_dif_sat_sva_1, return_add_generic_AC_RND_CONV_false_15_e_dif_sat_sva,
      return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva, {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_4_or_97_cse , return_add_generic_AC_RND_CONV_false_4_or_98_nl
      , (fsm_output[12]) , (fsm_output[39]) , (fsm_output[43]) , or_2189_nl , return_add_generic_AC_RND_CONV_false_12_res_mant_or_cse});
  wire return_add_generic_AC_RND_CONV_false_2_or_nl;
  wire [54:0] nl_return_add_generic_AC_RND_CONV_false_15_lshift_rg_a;
  assign return_add_generic_AC_RND_CONV_false_2_or_nl = return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_or_1_cse
      | return_add_generic_AC_RND_CONV_false_2_or_2_seb;
  assign nl_return_add_generic_AC_RND_CONV_false_15_lshift_rg_a = signext_55_54({return_add_generic_AC_RND_CONV_false_2_or_2_seb
      , return_add_generic_AC_RND_CONV_false_2_or_nl , 52'b1111111111111111111111111111111111111111111111111111});
  wire return_add_generic_AC_RND_CONV_false_2_and_nl;
  wire return_add_generic_AC_RND_CONV_false_2_mux1h_2_nl;
  wire return_add_generic_AC_RND_CONV_false_2_and_1_nl;
  wire return_add_generic_AC_RND_CONV_false_2_mux1h_3_nl;
  wire[2:0] return_add_generic_AC_RND_CONV_false_2_mux1h_5_nl;
  wire return_add_generic_AC_RND_CONV_false_2_mux1h_4_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_15_lshift_rg_s;
  assign return_add_generic_AC_RND_CONV_false_2_mux1h_2_nl = MUX1HOT_s_1_4_2((return_add_generic_AC_RND_CONV_false_2_e_dif_sat_sva_1[5]),
      (return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_cse[5]), return_mult_generic_AC_RND_CONV_false_if_or_3_cse,
      (return_add_generic_AC_RND_CONV_false_9_e_dif_sat_sva_1[5]), {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse , return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_or_1_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse});
  assign return_add_generic_AC_RND_CONV_false_2_and_nl = return_add_generic_AC_RND_CONV_false_2_mux1h_2_nl
      & (~ (fsm_output[54]));
  assign return_add_generic_AC_RND_CONV_false_2_mux1h_3_nl = MUX1HOT_s_1_4_2((return_add_generic_AC_RND_CONV_false_2_e_dif_sat_sva_1[4]),
      (return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_cse[4]), (return_mult_generic_AC_RND_CONV_false_if_nand_1_cse[3]),
      (return_add_generic_AC_RND_CONV_false_9_e_dif_sat_sva_1[4]), {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse , return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_or_1_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse});
  assign return_add_generic_AC_RND_CONV_false_2_and_1_nl = return_add_generic_AC_RND_CONV_false_2_mux1h_3_nl
      & (~ (fsm_output[54]));
  assign return_add_generic_AC_RND_CONV_false_2_mux1h_5_nl = MUX1HOT_v_3_5_2((return_add_generic_AC_RND_CONV_false_2_e_dif_sat_sva_1[3:1]),
      (return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_cse[3:1]), (return_mult_generic_AC_RND_CONV_false_if_nand_1_cse[2:0]),
      (return_add_generic_AC_RND_CONV_false_9_e_dif_sat_sva_1[3:1]), (~ (z_out_27[3:1])),
      {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse
      , return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_or_1_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_2_mux1h_4_nl = MUX1HOT_s_1_5_2((return_add_generic_AC_RND_CONV_false_2_e_dif_sat_sva_1[0]),
      (return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_cse[0]), return_mult_generic_AC_RND_CONV_false_if_or_cse,
      (return_add_generic_AC_RND_CONV_false_9_e_dif_sat_sva_1[0]), (~ (z_out_27[0])),
      {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse
      , return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_or_1_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse , (fsm_output[54])});
  assign nl_return_add_generic_AC_RND_CONV_false_15_lshift_rg_s = {return_add_generic_AC_RND_CONV_false_2_and_nl
      , return_add_generic_AC_RND_CONV_false_2_and_1_nl , return_add_generic_AC_RND_CONV_false_2_mux1h_5_nl
      , return_add_generic_AC_RND_CONV_false_2_mux1h_4_nl};
  wire[51:0] return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_mux_3_nl;
  wire[51:0] return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_1_not_1_nl;
  wire [105:0] nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_a;
  assign return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_mux_3_nl
      = MUX_v_52_2_2((z_out_21[103:52]), (out_f_d_rsci_q_d[51:0]), fsm_output[54]);
  assign return_mult_generic_AC_RND_CONV_false_if_1_not_1_nl = ~ (fsm_output[54]);
  assign return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_and_1_nl
      = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000, (z_out_21[51:0]),
      return_mult_generic_AC_RND_CONV_false_if_1_not_1_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_a = {return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_and_cse
      , return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_mux_2_cse
      , return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_mux_3_nl
      , return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_and_1_nl};
  wire return_mult_generic_AC_RND_CONV_false_if_1_or_3_nl;
  wire [5:0] nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_s;
  assign return_mult_generic_AC_RND_CONV_false_if_1_or_3_nl = ((z_out_29[12]) & (fsm_output[10]))
      | ((z_out_29[12]) & (fsm_output[12])) | ((z_out_29[12]) & (fsm_output[14]))
      | ((z_out_29[12]) & (fsm_output[35])) | ((z_out_29[12]) & (fsm_output[37]))
      | ((z_out_29[12]) & (fsm_output[39])) | ((z_out_29[11]) & (fsm_output[54]));
  assign nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_s = MUX_v_6_2_2(rtn_out_1,
      (z_out_27[5:0]), return_mult_generic_AC_RND_CONV_false_if_1_or_3_nl);
  wire[50:0] return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_1_nl;
  wire [53:0] nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_a;
  assign return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_1_nl
      = MUX_v_51_2_2((z_out_21[103:53]), (out_f_d_rsci_q_d[51:1]), fsm_output[54]);
  assign nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_a = {return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_and_cse
      , return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_mux_2_cse
      , return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_1_nl
      , 1'b0};
  wire return_mult_generic_AC_RND_CONV_false_else_1_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_and_nl;
  wire[2:0] return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_nl;
  wire return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_3_nl;
  wire [5:0] nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_s;
  assign return_mult_generic_AC_RND_CONV_false_else_1_and_nl = return_mult_generic_AC_RND_CONV_false_if_or_3_cse
      & (~ (fsm_output[54]));
  assign return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_and_nl
      = (return_mult_generic_AC_RND_CONV_false_if_nand_1_cse[3]) & (~ (fsm_output[54]));
  assign return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_nl
      = MUX_v_3_2_2((return_mult_generic_AC_RND_CONV_false_if_nand_1_cse[2:0]), (~
      (z_out_27[3:1])), fsm_output[54]);
  assign return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_3_nl
      = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_if_or_cse, (~ (z_out_27[0])),
      fsm_output[54]);
  assign nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_s = {return_mult_generic_AC_RND_CONV_false_else_1_and_nl
      , return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_and_nl
      , return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_nl
      , return_mult_generic_AC_RND_CONV_false_else_1_return_mult_generic_AC_RND_CONV_false_else_1_mux_3_nl};
  wire return_add_generic_AC_RND_CONV_false_4_mux1h_6_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_104_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux1h_20_nl;
  wire[49:0] return_add_generic_AC_RND_CONV_false_4_mux1h_21_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_111_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_92_nl;
  wire return_add_generic_AC_RND_CONV_false_4_or_93_nl;
  wire return_add_generic_AC_RND_CONV_false_4_mux1h_22_nl;
  wire [56:0] nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_a;
  assign return_add_generic_AC_RND_CONV_false_4_or_104_nl = return_add_generic_AC_RND_CONV_false_4_or_86_cse
      | ((~ and_dcpl_348) & (fsm_output[37]));
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_6_nl = MUX1HOT_s_1_12_2(return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_6_cse,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx1, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx2,
      return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_10_exp_mux_5_cse,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx6,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx7, return_add_generic_AC_RND_CONV_false_19_op2_mu_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_13_mux_25_cse, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_52_lpi_3_dfm, {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[12]) , (fsm_output[18]) ,
      return_add_generic_AC_RND_CONV_false_4_or_104_nl , (fsm_output[30]) , (fsm_output[32])
      , and_1589_cse , (fsm_output[43]) , or_tmp_1248 , return_add_generic_AC_RND_CONV_false_4_or_87_cse});
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_20_nl = MUX1HOT_s_1_12_2((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[50]),
      (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[50]), (return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_50_mx0,
      return_add_generic_AC_RND_CONV_false_5_op_smaller_mux_1_cse, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm,
      (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[50]),
      return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_50_mx0,
      return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_2_cse, (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[50]),
      return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_51_lpi_3_dfm, {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[12]) , (fsm_output[18]) ,
      return_add_generic_AC_RND_CONV_false_4_or_86_cse , (fsm_output[30]) , (fsm_output[32])
      , (fsm_output[37]) , (fsm_output[43]) , or_tmp_1248 , return_add_generic_AC_RND_CONV_false_4_or_87_cse});
  assign return_add_generic_AC_RND_CONV_false_4_or_111_nl = return_add_generic_AC_RND_CONV_false_10_exp_and_2_cse
      | or_tmp_1248;
  assign return_add_generic_AC_RND_CONV_false_4_or_92_nl = (fsm_output[19]) | or_tmp_1251;
  assign return_add_generic_AC_RND_CONV_false_4_or_93_nl = or_tmp_1249 | or_tmp_1250;
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_21_nl = MUX1HOT_v_50_12_2((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[49:0]),
      (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[49:0]),
      (return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0,
      (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49:0]), return_add_generic_AC_RND_CONV_false_10_op2_mu_1_50_1_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1, (return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      (return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[49:0]),
      return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0,
      return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1,
      {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[12]) , return_add_generic_AC_RND_CONV_false_4_or_111_nl
      , return_add_generic_AC_RND_CONV_false_10_exp_and_3_cse , return_add_generic_AC_RND_CONV_false_4_or_92_nl
      , (fsm_output[30]) , (fsm_output[32]) , (fsm_output[37]) , (fsm_output[43])
      , return_add_generic_AC_RND_CONV_false_4_or_93_nl});
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_22_nl = MUX1HOT_s_1_11_2(return_add_generic_AC_RND_CONV_false_4_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx1, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2,
      return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_0_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_1_op_bigger_mux_4_cse,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx5,
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx6, return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_0_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_1_op_bigger_mux_5_cse, return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm,
      {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[12]) , (fsm_output[18]) , return_add_generic_AC_RND_CONV_false_4_or_95_cse
      , (fsm_output[30]) , (fsm_output[32]) , (fsm_output[37]) , (fsm_output[43])
      , return_add_generic_AC_RND_CONV_false_4_or_87_cse});
  assign nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_a = {1'b0 , return_add_generic_AC_RND_CONV_false_4_mux1h_6_nl
      , return_add_generic_AC_RND_CONV_false_4_mux1h_20_nl , return_add_generic_AC_RND_CONV_false_4_mux1h_21_nl
      , return_add_generic_AC_RND_CONV_false_4_mux1h_22_nl , 3'b000};
  wire return_add_generic_AC_RND_CONV_false_4_or_106_nl;
  wire [5:0] nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_s;
  assign return_add_generic_AC_RND_CONV_false_4_or_106_nl = (fsm_output[7]) | (fsm_output[18])
      | (fsm_output[32]);
  assign nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_s = MUX1HOT_v_6_7_2(return_add_generic_AC_RND_CONV_false_4_e_dif_sat_sva_1,
      return_add_generic_AC_RND_CONV_false_e_dif_sat_or_cse, return_add_generic_AC_RND_CONV_false_21_e_dif_sat_or_cse,
      return_add_generic_AC_RND_CONV_false_6_e_dif_sat_sva_1, return_add_generic_AC_RND_CONV_false_15_e_dif_sat_sva,
      return_add_generic_AC_RND_CONV_false_23_e_dif_sat_sva_1, return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva,
      {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , return_add_generic_AC_RND_CONV_false_4_or_97_cse
      , return_add_generic_AC_RND_CONV_false_4_or_106_nl , (fsm_output[12]) , return_add_generic_AC_RND_CONV_false_4_or_95_cse
      , (fsm_output[43]) , return_add_generic_AC_RND_CONV_false_4_or_87_cse});
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_return_mult_generic_AC_RND_CONV_false_1_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_if_return_mult_generic_AC_RND_CONV_false_2_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_3_if_return_mult_generic_AC_RND_CONV_false_3_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_4_if_return_mult_generic_AC_RND_CONV_false_4_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_5_if_return_mult_generic_AC_RND_CONV_false_5_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_2_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_5_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_6_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_8_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_11_nl;
  wire[50:0] return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_2_nl;
  wire mux_11_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_mux_5_nl;
  wire[49:0] return_mult_generic_AC_RND_CONV_false_if_mux1h_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_nor_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_1_if_and_1_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_12_nl;
  wire return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_13_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_if_and_nl;
  wire return_mult_generic_AC_RND_CONV_false_2_if_and_1_nl;
  wire [52:0] nl_leading_sign_53_0_rg_mantissa;
  assign return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_nl
      = return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm & return_extract_12_return_extract_12_or_1_cse_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_1_if_return_mult_generic_AC_RND_CONV_false_1_if_and_nl
      = return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm & return_extract_13_return_extract_13_or_1_cse_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_2_if_return_mult_generic_AC_RND_CONV_false_2_if_and_nl
      = return_extract_19_return_extract_19_or_sva_1 & BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm;
  assign return_mult_generic_AC_RND_CONV_false_3_if_return_mult_generic_AC_RND_CONV_false_3_if_and_nl
      = return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm & return_extract_44_return_extract_44_or_1_cse_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_4_if_return_mult_generic_AC_RND_CONV_false_4_if_and_nl
      = return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm & return_extract_45_return_extract_45_or_1_cse_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_5_if_return_mult_generic_AC_RND_CONV_false_5_if_and_nl
      = return_extract_51_return_extract_51_or_sva_1 & BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_nl
      = MUX1HOT_s_1_7_2(return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_and_nl,
      return_mult_generic_AC_RND_CONV_false_1_if_return_mult_generic_AC_RND_CONV_false_1_if_and_nl,
      return_mult_generic_AC_RND_CONV_false_2_if_return_mult_generic_AC_RND_CONV_false_2_if_and_nl,
      return_mult_generic_AC_RND_CONV_false_3_if_return_mult_generic_AC_RND_CONV_false_3_if_and_nl,
      return_mult_generic_AC_RND_CONV_false_4_if_return_mult_generic_AC_RND_CONV_false_4_if_and_nl,
      return_mult_generic_AC_RND_CONV_false_5_if_return_mult_generic_AC_RND_CONV_false_5_if_and_nl,
      return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp,
      {(fsm_output[10]) , (fsm_output[12]) , (fsm_output[14]) , (fsm_output[35])
      , (fsm_output[37]) , (fsm_output[39]) , (fsm_output[54])});
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_nl =
      (~ return_extract_12_return_extract_12_or_1_cse_sva_1) & (fsm_output[10]);
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_nl = (return_extract_12_return_extract_12_or_1_cse_sva_1
      & (fsm_output[10])) | (return_extract_44_return_extract_44_or_1_cse_sva_1 &
      (fsm_output[35]));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_2_nl
      = (~ return_extract_13_return_extract_13_or_1_cse_sva_1) & (fsm_output[12]);
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_1_nl =
      (return_extract_13_return_extract_13_or_1_cse_sva_1 & (fsm_output[12])) | (return_extract_45_return_extract_45_or_1_cse_sva_1
      & (fsm_output[37]));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_2_nl =
      ((~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm) & (fsm_output[14]))
      | ((~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm) & (fsm_output[39]));
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_5_nl
      = BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm & (fsm_output[14]);
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_6_nl
      = (~ return_extract_44_return_extract_44_or_1_cse_sva_1) & (fsm_output[35]);
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_8_nl
      = (~ return_extract_45_return_extract_45_or_1_cse_sva_1) & (fsm_output[37]);
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_11_nl
      = BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm & (fsm_output[39]);
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_1_nl
      = MUX1HOT_s_1_10_2(return_extract_15_return_extract_15_nor_cse_sva_mx1, drf_qr_lval_14_smx_0_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_3_r_nan_mux1h_cse, drf_qr_lval_15_smx_0_lpi_3_dfm,
      (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[51]), return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0,
      return_extract_15_return_extract_15_nor_cse_sva_mx2, return_add_generic_AC_RND_CONV_false_16_r_nan_mux1h_cse,
      return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0, (return_mult_generic_AC_RND_CONV_false_6_if_conc_itm_51_0[51]),
      {return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_nl , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_2_nl ,
      return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_1_nl , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_or_2_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_5_nl ,
      return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_6_nl , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_8_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_11_nl
      , (fsm_output[54])});
  assign return_mult_generic_AC_RND_CONV_false_if_mux_5_nl = MUX_s_1_2_2((stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0[50]),
      (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1[50]), fsm_output[35]);
  assign mux_11_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_if_mux_5_nl,
      return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_0, return_mult_generic_AC_RND_CONV_false_if_mux_6_ssc);
  assign return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_nor_nl
      = ~((fsm_output[35]) | return_mult_generic_AC_RND_CONV_false_if_mux_6_ssc);
  assign return_mult_generic_AC_RND_CONV_false_if_and_1_nl = (fsm_output[35]) & (~
      return_mult_generic_AC_RND_CONV_false_if_mux_6_ssc);
  assign return_mult_generic_AC_RND_CONV_false_if_mux1h_nl = MUX1HOT_v_50_3_2((stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0[49:0]),
      (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1[49:0]), return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1,
      {return_mult_generic_AC_RND_CONV_false_if_return_mult_generic_AC_RND_CONV_false_if_nor_nl
      , return_mult_generic_AC_RND_CONV_false_if_and_1_nl , return_mult_generic_AC_RND_CONV_false_if_mux_6_ssc});
  assign return_mult_generic_AC_RND_CONV_false_1_if_and_nl = (~ (fsm_output[37]))
      & (~ return_mult_generic_AC_RND_CONV_false_1_if_mux_6_tmp) & or_dcpl_404;
  assign return_mult_generic_AC_RND_CONV_false_1_if_and_1_nl = (fsm_output[37]) &
      (~ return_mult_generic_AC_RND_CONV_false_1_if_mux_6_tmp) & or_dcpl_404;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_12_nl
      = return_mult_generic_AC_RND_CONV_false_1_if_mux_6_tmp & or_dcpl_404;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_13_nl
      = (~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm) & BUTTERFLY_i_or_4_cse;
  assign return_mult_generic_AC_RND_CONV_false_2_if_and_nl = (~ (fsm_output[39]))
      & BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm & BUTTERFLY_i_or_4_cse;
  assign return_mult_generic_AC_RND_CONV_false_2_if_and_1_nl = (fsm_output[39]) &
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm & BUTTERFLY_i_or_4_cse;
  assign return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_2_nl
      = MUX1HOT_v_51_8_2(({mux_11_nl , return_mult_generic_AC_RND_CONV_false_if_mux1h_nl}),
      stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0, stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0,
      return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm, (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[50:0]),
      return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1,
      (return_mult_generic_AC_RND_CONV_false_6_if_conc_itm_51_0[50:0]), {or_dcpl_548
      , return_mult_generic_AC_RND_CONV_false_1_if_and_nl , return_mult_generic_AC_RND_CONV_false_1_if_and_1_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_12_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_and_13_nl
      , return_mult_generic_AC_RND_CONV_false_2_if_and_nl , return_mult_generic_AC_RND_CONV_false_2_if_and_1_nl
      , (fsm_output[54])});
  assign nl_leading_sign_53_0_rg_mantissa = {return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_1_nl
      , return_mult_generic_AC_RND_CONV_false_if_leading_sign_53_0_rtn_mux1h_2_nl};
  wire [79:0] nl_stage_run_out1_rsci_inst_out1_rsci_idat;
  assign nl_stage_run_out1_rsci_inst_out1_rsci_idat = {out1_rsci_idat_79_64 , out1_rsci_idat_63
      , out1_rsci_idat_62_52 , out1_rsci_idat_51 , out1_rsci_idat_50_0};
  wire  nl_stage_run_run_fsm_inst_for_1_C_2_tr0;
  assign nl_stage_run_run_fsm_inst_for_1_C_2_tr0 = z_out_19[10];
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd16)) mode1_rsci (
      .dat(mode1_rsc_dat),
      .idat(mode1_rsci_idat)
    );
  

`ifdef USE_PDK_ROM
wire [56:0] O_1_out_57;
wire [56:0] O_1_out_1_57;
ROM_1024x142 ROM_1024x142(
.CLK(clk),
.CEN(1'b1),//not sure
.I(z_out_7),
.O({U_ROM_1i10_1o14_out_2,U_ROM_1i10_1o14_out_3,O_1_out_57,O_1_out_1_57})
);

assign O_1_out={z_out_7[0],1'b0,{5{O_1_out_57[56]}},O_1_out_57};
assign O_1_out_1={{5{O_1_out_1_57[56]}},O_1_out_1_57};

`else
  ROM_1i10_1o14_64308806abd59d677de1cc2043c30c27bd  U_ROM_1i10_1o14_486610990d9cceb357c747b53d9fad3232_rg
      (
      .I_1(z_out_7),
      .O_1(U_ROM_1i10_1o14_out_2)
    );
  ROM_1i10_1o14_281e23127cb7ddaedd69e0bbd10d0137bd  U_ROM_1i10_1o14_65c485e62ebcbda02b981400037c62ce32_rg
      (
      .I_1(z_out_7),
      .O_1(U_ROM_1i10_1o14_out_3)
    );
  ROM_1i10_1o64_a49ff3631daca65e62d175dd412366e6bd  U_ROM_1i10_1o64_198d068ad119e36f3a1745eecd5c3e2132_rg
      (
      .I_1(z_out_7),
      .O_1(O_1_out)
    );
  ROM_1i10_1o62_e041a31844d9eff753e17f0437c907cdbd  U_ROM_1i10_1o62_1843679b7562278e9c543f644738904f32_rg
      (
      .I_1(z_out_7),
      .O_1(O_1_out_1)
    );
`endif
    
  mgc_shift_l_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_10_lshift_1_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_10_lshift_1_rg_s[5:0]),
      .z(z_out_15)
    );
  mgc_shift_l_v5 #(.width_a(32'sd55),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd55)) return_add_generic_AC_RND_CONV_false_10_lshift_rg (
      .a(55'b1111111111111111111111111111111111111111111111111111111),
      .s(nl_return_add_generic_AC_RND_CONV_false_10_lshift_rg_s[5:0]),
      .z(z_out_16)
    );
  mgc_shift_l_v5 #(.width_a(32'sd55),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd55)) return_add_generic_AC_RND_CONV_false_15_lshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_15_lshift_rg_a[54:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_15_lshift_rg_s[5:0]),
      .z(z_out_17)
    );
  mgc_shift_l_v5 #(.width_a(32'sd106),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd106)) return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg (
      .a(nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_a[105:0]),
      .s(nl_return_mult_generic_AC_RND_CONV_false_1_if_1_lshift_rg_s[5:0]),
      .z(z_out_18)
    );
  leading_sign_57_0_1_0  leading_sign_57_0_1_0_rg (
      .mantissa(z_out_30),
      .all_same(all_same_out),
      .rtn(rtn_out)
    );
  mgc_shift_r_v5 #(.width_a(32'sd54),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd54)) return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg (
      .a(nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_a[53:0]),
      .s(nl_return_mult_generic_AC_RND_CONV_false_1_else_1_rshift_rg_s[5:0]),
      .z(z_out_42)
    );
  mgc_shift_r_v5 #(.width_a(32'sd57),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd57)) return_add_generic_AC_RND_CONV_false_10_rshift_rg (
      .a(nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_a[56:0]),
      .s(nl_return_add_generic_AC_RND_CONV_false_10_rshift_rg_s[5:0]),
      .z(z_out_43)
    );
  leading_sign_53_0  leading_sign_53_0_rg (
      .mantissa(nl_leading_sign_53_0_rg_mantissa[52:0]),
      .rtn(rtn_out_1)
    );
  stage_run_ap_start_rsci stage_run_ap_start_rsci_inst (
      .ap_start_rsc_dat(ap_start_rsc_dat),
      .ap_start_rsc_vld(ap_start_rsc_vld),
      .ap_start_rsc_rdy(ap_start_rsc_rdy),
      .ap_start_rsci_oswt(reg_ap_start_rsci_iswt0_cse),
      .ap_start_rsci_wen_comp(ap_start_rsci_wen_comp)
    );
  stage_run_ap_done_rsci stage_run_ap_done_rsci_inst (
      .ap_done_rsc_dat(ap_done_rsc_dat),
      .ap_done_rsc_vld(ap_done_rsc_vld),
      .ap_done_rsc_rdy(ap_done_rsc_rdy),
      .ap_done_rsci_oswt(reg_out_u_triosy_obj_iswt0_cse),
      .ap_done_rsci_wen_comp(ap_done_rsci_wen_comp)
    );
  stage_run_wait_dp stage_run_wait_dp_inst (
      .in_f_d_rsci_en_d(in_f_d_rsci_en_d),
      .in_u_rsci_en_d(in_u_rsci_en_d),
      .out_f_d_rsci_en_d(out_f_d_rsci_en_d),
      .out_u_rsci_en_d(out_u_rsci_en_d),
      .run_wen(run_wen),
      .in_f_d_rsci_cgo(reg_in_f_d_rsci_cgo_ir_cse),
      .in_f_d_rsci_cgo_ir_unreg(or_1181_rmff),
      .in_u_rsci_cgo(reg_in_u_rsci_cgo_ir_cse),
      .in_u_rsci_cgo_ir_unreg(or_1180_rmff),
      .out_f_d_rsci_cgo(reg_out_f_d_rsci_cgo_ir_cse),
      .out_f_d_rsci_cgo_ir_unreg(or_1179_rmff),
      .out_u_rsci_cgo(reg_out_u_rsci_cgo_ir_cse),
      .out_u_rsci_cgo_ir_unreg(or_1178_rmff)
    );
  stage_run_out1_rsci stage_run_out1_rsci_inst (
      .out1_rsc_dat(out1_rsc_dat),
      .out1_rsc_vld(out1_rsc_vld),
      .out1_rsc_rdy(out1_rsc_rdy),
      .out1_rsci_oswt(reg_out1_rsci_iswt0_cse),
      .out1_rsci_wen_comp(out1_rsci_wen_comp),
      .out1_rsci_idat(nl_stage_run_out1_rsci_inst_out1_rsci_idat[79:0])
    );
  stage_run_mode1_triosy_obj stage_run_mode1_triosy_obj_inst (
      .mode1_triosy_lz(mode1_triosy_lz),
      .run_wten(run_wten),
      .mode1_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_in_f_d_triosy_obj stage_run_in_f_d_triosy_obj_inst (
      .in_f_d_triosy_lz(in_f_d_triosy_lz),
      .run_wten(run_wten),
      .in_f_d_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_in_u_triosy_obj stage_run_in_u_triosy_obj_inst (
      .in_u_triosy_lz(in_u_triosy_lz),
      .run_wten(run_wten),
      .in_u_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_out_f_d_triosy_obj stage_run_out_f_d_triosy_obj_inst (
      .out_f_d_triosy_lz(out_f_d_triosy_lz),
      .run_wten(run_wten),
      .out_f_d_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_out_u_triosy_obj stage_run_out_u_triosy_obj_inst (
      .out_u_triosy_lz(out_u_triosy_lz),
      .run_wten(run_wten),
      .out_u_triosy_obj_iswt0(reg_out_u_triosy_obj_iswt0_cse)
    );
  stage_run_staller stage_run_staller_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .ap_start_rsci_wen_comp(ap_start_rsci_wen_comp),
      .ap_done_rsci_wen_comp(ap_done_rsci_wen_comp),
      .out1_rsci_wen_comp(out1_rsci_wen_comp)
    );
  stage_run_run_fsm stage_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .for_C_0_tr0(for_i_0_sva),
      .BUTTERFLY_C_24_tr0(and_83_cse),
      .BUTTERFLY_C_24_tr1(nor_158_cse),
      .BUTTERFLY_1_C_24_tr0(and_83_cse),
      .BUTTERFLY_1_C_24_tr1(nor_158_cse),
      .for_1_C_2_tr0(nl_stage_run_run_fsm_inst_for_1_C_2_tr0)
    );
  assign for_1_if_and_ssc = run_wen & (or_tmp_61 | out1_rsci_idat_63_0_mx0c1 | out1_rsci_idat_63_0_mx0c2);
  assign or_1178_rmff = (stage_PE_1_and_cse & (or_dcpl_92 | (fsm_output[30]))) |
      (nor_3_cse & ((fsm_output[35:34]!=2'b00))) | (~(mode_lpi_1_dfm | (~((fsm_output[3])
      | (fsm_output[33]) | or_dcpl_95)))) | (operator_16_false_operator_16_false_nor_cse_sva
      & or_dcpl_11);
  assign or_1179_rmff = (stage_PE_1_and_1_tmp & (or_dcpl_102 | or_dcpl_101 | or_dcpl_99
      | or_dcpl_92)) | (and_dcpl_1 & ((fsm_output[52:51]!=2'b00) | or_dcpl_108 |
      or_dcpl_106 | or_dcpl_105)) | (mode_lpi_1_dfm & ((fsm_output[3]) | (fsm_output[7])
      | (fsm_output[6]) | or_dcpl_95)) | (or_dcpl_115 & or_dcpl_11);
  assign or_1180_rmff = (and_dcpl_146 & (fsm_output[55])) | (stage_PE_1_and_cse &
      ((fsm_output[7:5]!=3'b000))) | (~(mode_lpi_1_dfm | (~((fsm_output[28]) | (fsm_output[8])
      | or_dcpl_118)))) | and_592_cse | (nor_3_cse & ((fsm_output[10:9]!=2'b00)));
  assign or_1181_rmff = (mode_lpi_1_dfm & ((fsm_output[28]) | (fsm_output[32]) |
      (fsm_output[31]) | or_dcpl_118)) | (and_dcpl_1 & ((fsm_output[27:26]!=2'b00)
      | or_dcpl_128 | or_dcpl_126 | or_dcpl_125)) | (stage_PE_1_and_1_tmp & (or_dcpl_136
      | or_dcpl_135 | or_dcpl_133 | or_dcpl_132)) | and_592_cse;
  assign or_200_cse = (fsm_output[32]) | (fsm_output[30]);
  assign or_1205_ssc = (fsm_output[45]) | (fsm_output[31]) | (fsm_output[4]);
  assign or_1206_ssc = (fsm_output[33]) | (fsm_output[5]);
  assign and_654_ssc = inverse_lpi_1_dfm_1 & (fsm_output[6]);
  assign or_1208_ssc = (fsm_output[53]) | (fsm_output[49]) | (fsm_output[41]) | ((~
      inverse_lpi_1_dfm_1) & (fsm_output[6]));
  assign or_1209_ssc = or_dcpl_148 | (fsm_output[43]);
  assign or_219_cse = (fsm_output[7]) | (fsm_output[5]);
  assign or_1231_ssc = (fsm_output[20]) | (fsm_output[6]) | (fsm_output[29]);
  assign or_1232_ssc = (fsm_output[8]) | (fsm_output[30]);
  assign or_1233_ssc = ((~ inverse_lpi_1_dfm_1) & (fsm_output[31])) | (fsm_output[53])
      | (fsm_output[24]) | (fsm_output[16]);
  assign or_1234_ssc = or_dcpl_166 | (fsm_output[18]);
  assign and_720_ssc = inverse_lpi_1_dfm_1 & (fsm_output[31]);
  assign return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_nor_cse
      = ~((~ mode_lpi_1_dfm) | (z_out_27[12]));
  assign return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse
      = ~((z_out_8[11:0]==12'b011111111111));
  assign operator_16_false_and_cse = run_wen & ((fsm_output[1]) | (fsm_output[56])
      | (fsm_output[0]));
  assign t_in_and_cse = run_wen & ((~(nor_158_cse | and_dcpl_210)) | (fsm_output[1]));
  assign mode_and_cse = run_wen & (~(and_dcpl_214 & and_dcpl_211 & (~ (fsm_output[54]))));
  assign stage_PE_1_and_2_cse = run_wen & (~(and_dcpl_213 & and_dcpl_165 & and_dcpl_217));
  assign and_83_cse = (and_2334_cse | (BUTTERFLY_1_n_9_0_sva_1[9])) & t_in_10_0_lpi_1_dfm_1_1
      & (~(t_in_10_0_lpi_1_dfm_1_10 | t_in_10_0_lpi_1_dfm_1_9 | t_in_10_0_lpi_1_dfm_1_8
      | t_in_10_0_lpi_1_dfm_1_7 | t_in_10_0_lpi_1_dfm_1_6 | t_in_10_0_lpi_1_dfm_1_5
      | t_in_10_0_lpi_1_dfm_1_4 | t_in_10_0_lpi_1_dfm_1_3 | t_in_10_0_lpi_1_dfm_1_2));
  assign return_extract_26_m_zero_sva_2 = ~((in_f_d_rsci_q_d[51:0]!=52'b0000000000000000000000000000000000000000000000000000));
  assign return_extract_15_and_3_cse = run_wen & (~(or_dcpl_425 | or_dcpl_420));
  assign return_extract_15_m_zero_mux1h_cse = ~(return_add_generic_AC_RND_CONV_false_4_m_r_51_lpi_3_dfm_1
      | (return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign or_1375_cse = (fsm_output[32]) | (fsm_output[29]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_6_nl = MUX_s_1_2_2(and_dcpl_260,
      and_dcpl_264, fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_cse = run_wen & ((~(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_6_nl
      | and_1013_cse)) | (fsm_output[3]) | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[10])
      | (fsm_output[16]) | (fsm_output[28]) | (fsm_output[30]) | (fsm_output[32])
      | (fsm_output[35]) | (fsm_output[41]) | (fsm_output[43]));
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse = (fsm_output[3])
      | (fsm_output[28]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_6_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[50]),
      and_dcpl_261);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_12_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[50]), and_dcpl_265);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_5_cse = (~ and_dcpl_257)
      & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_6_cse = and_dcpl_257
      & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_7_cse = (~ and_dcpl_258)
      & (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_11_cse = (~ and_dcpl_262)
      & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse = and_dcpl_258
      & (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse = (~ and_dcpl_259)
      & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse = and_dcpl_259
      & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse = and_dcpl_263
      & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse = and_dcpl_262
      & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_13_cse = (~ and_dcpl_263)
      & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_7_cse = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_13_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse = (~ and_dcpl_266)
      & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_16_cse = and_dcpl_266
      & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_21_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1, and_dcpl_261);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_27_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1, and_dcpl_265);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_24_cse = return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_tmp
      & (fsm_output[10]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_23_cse = (~ return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_tmp)
      & (fsm_output[10]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_30_cse = return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp
      & (fsm_output[35]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_29_cse = (~ return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp)
      & (fsm_output[35]);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_cse = run_wen & (~(or_dcpl_488
      | (fsm_output[42]) | (fsm_output[18]) | (fsm_output[17])));
  assign return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_2_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_261);
  assign return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_3_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_265);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_cse = (~ and_dcpl_268)
      & (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_4_cse = (~ and_dcpl_267)
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse = and_dcpl_267
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_cse = and_dcpl_268
      & (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_6_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_17_op1_mu_52_lpi_3_dfm_1,
      stage_PE_1_gm_im_d_mux_cse, and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_cse = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[50]),
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0, and_dcpl_261);
  assign return_add_generic_AC_RND_CONV_false_5_op_smaller_mux_cse = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[50]),
      return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0, and_dcpl_265);
  assign return_add_generic_AC_RND_CONV_false_22_op1_mu_mux_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_22_op1_mu_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0, and_dcpl_261);
  assign return_add_generic_AC_RND_CONV_false_22_op1_mu_mux_1_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_22_op1_mu_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0, and_dcpl_265);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_12_cse = (~ return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp)
      & (fsm_output[10]);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_13_cse = return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp
      & (fsm_output[10]);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_14_cse = (~ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp)
      & (fsm_output[35]);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_and_15_cse = return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp
      & (fsm_output[35]);
  assign BUTTERFLY_1_fiy_mux1h_2_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1,
      (stage_PE_1_x_re_d_sva[52]), and_dcpl_261);
  assign BUTTERFLY_1_fiy_mux1h_6_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1,
      (stage_PE_1_x_re_d_sva[52]), and_dcpl_265);
  assign BUTTERFLY_1_fiy_or_1_cse = (fsm_output[17]) | (fsm_output[42]) | or_dcpl_397;
  assign BUTTERFLY_1_n_and_cse = run_wen & (~(and_dcpl_210 & (~((fsm_output[55])
      | (fsm_output[56]) | (fsm_output[0]))) & and_dcpl_217 & and_dcpl_284));
  assign return_add_generic_AC_RND_CONV_false_10_exp_and_2_cse = (~ and_dcpl_326)
      & (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_10_exp_and_5_cse = and_dcpl_265 & (fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_10_exp_and_4_cse = (~ and_dcpl_265)
      & (fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_10_exp_and_3_cse = and_dcpl_326 & (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_and_cse = (~ inverse_lpi_1_dfm_1)
      & or_dcpl_548;
  assign return_add_generic_AC_RND_CONV_false_9_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_9_op1_smaller_oelse_and_cse
      = z_out_33_52 & return_add_generic_AC_RND_CONV_false_9_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_9_op1_smaller_return_add_generic_AC_RND_CONV_false_9_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_9_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_9_op1_smaller_oelse_and_cse
      | (z_out_23[11]);
  assign return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_and_cse
      = z_out_34_52 & return_add_generic_AC_RND_CONV_false_23_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_25_op1_smaller_return_add_generic_AC_RND_CONV_false_25_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_and_cse
      | (z_out_25[11]);
  assign return_add_generic_AC_RND_CONV_false_17_and_2_m1c = or_dcpl_549 & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  assign return_add_generic_AC_RND_CONV_false_17_and_4_m1c = or_dcpl_566 & (fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_17_and_6_m1c = or_dcpl_568 & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_17_and_3_cse = (~ or_dcpl_566) & (fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_17_and_5_cse = (~ or_dcpl_568) & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_17_and_9_cse = (~ return_add_generic_AC_RND_CONV_false_9_op1_smaller_return_add_generic_AC_RND_CONV_false_9_op1_smaller_or_cse)
      & return_add_generic_AC_RND_CONV_false_17_and_4_m1c;
  assign return_add_generic_AC_RND_CONV_false_17_and_10_cse = return_add_generic_AC_RND_CONV_false_9_op1_smaller_return_add_generic_AC_RND_CONV_false_9_op1_smaller_or_cse
      & return_add_generic_AC_RND_CONV_false_17_and_4_m1c;
  assign return_add_generic_AC_RND_CONV_false_17_and_11_cse = (~ return_add_generic_AC_RND_CONV_false_25_op1_smaller_return_add_generic_AC_RND_CONV_false_25_op1_smaller_or_cse)
      & return_add_generic_AC_RND_CONV_false_17_and_6_m1c;
  assign return_add_generic_AC_RND_CONV_false_17_and_12_cse = return_add_generic_AC_RND_CONV_false_25_op1_smaller_return_add_generic_AC_RND_CONV_false_25_op1_smaller_or_cse
      & return_add_generic_AC_RND_CONV_false_17_and_6_m1c;
  assign return_add_generic_AC_RND_CONV_false_9_e_dif_qelse_return_add_generic_AC_RND_CONV_false_9_e_dif_qelse_and_cse
      = (z_out_25[11]) & (z_out_23[11]);
  assign return_add_generic_AC_RND_CONV_false_21_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_1_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_21_e_dif_sat_or_cse = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_1_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_21_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_8_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_8_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_8_e_dif_sat_or_cse = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_8_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_8_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse = (fsm_output[16])
      | (fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse = (fsm_output[5])
      | (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse = (fsm_output[7])
      | (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_itm = MUX_v_51_2_2(stage_PE_1_gm_im_d_mux_2_cse,
      stage_PE_1_gm_re_d_mux_cse, and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_1_itm = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx1, and_dcpl_258);
  assign return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_2_itm = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx1,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm, and_dcpl_259);
  assign return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_7_itm = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm,
      return_extract_32_mux_4_cse, and_dcpl_262);
  assign return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_8_itm = MUX_v_51_2_2(return_extract_32_mux_4_cse,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm, and_dcpl_263);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse = MUX_v_51_2_2(stage_PE_1_gm_re_d_mux_cse,
      stage_PE_1_gm_im_d_mux_2_cse, and_dcpl_257);
  assign return_extract_32_or_1_tmp = return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx6c1
      | ((~ return_add_generic_AC_RND_CONV_false_13_return_add_generic_AC_RND_CONV_false_13_or_1_tmp)
      & return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx6c2);
  assign and_453_tmp = (~ return_add_generic_AC_RND_CONV_false_13_return_add_generic_AC_RND_CONV_false_13_or_1_tmp)
      & inverse_lpi_1_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_or_3_rgt = (fsm_output[4])
      | (fsm_output[6]) | (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_or_8_rgt = ((~ return_extract_32_or_1_tmp)
      & (fsm_output[30])) | ((~ and_453_tmp) & (fsm_output[31]));
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_or_9_rgt = (return_extract_32_or_1_tmp
      & (fsm_output[30])) | (and_453_tmp & (fsm_output[31]));
  assign return_extract_32_mux_4_cse = MUX_v_51_2_2((in_f_d_rsci_q_d[50:0]), (in_f_d_rsci_q_d[51:1]),
      return_add_generic_AC_RND_CONV_false_13_return_add_generic_AC_RND_CONV_false_13_or_1_tmp);
  assign and_522_cse = return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp
      & z_out_35_52;
  assign or_1144_cse = and_522_cse | (z_out_25[11]);
  assign nl_return_add_generic_AC_RND_CONV_false_5_ma1_lt_ma2_acc_2_nl = ({1'b1 ,
      (O_1_out[51:0])}) + conv_u2u_52_53(~ (O_1_out_1[51:0])) + 53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_5_ma1_lt_ma2_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_5_ma1_lt_ma2_acc_2_nl[52:0];
  assign and_416_cse = return_add_generic_AC_RND_CONV_false_4_e1_eq_e2_equal_tmp
      & (readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_5_ma1_lt_ma2_acc_2_nl));
  assign or_590_cse = and_416_cse | (return_add_generic_AC_RND_CONV_false_4_e_dif_acc_tmp[10]);
  assign or_46_cse = inverse_lpi_1_dfm_1 | (~ mode_lpi_1_dfm);
  assign BUTTERFLY_1_else_3_else_and_ssc = run_wen & (~ return_extract_26_exception_or_3_cse);
  assign and_933_nl = (~ inverse_lpi_1_dfm_1) & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  assign BUTTERFLY_1_else_3_else_mux1h_itm = MUX_v_14_2_2(U_ROM_1i10_1o14_out_2,
      U_ROM_1i10_1o14_out_3, and_933_nl);
  assign or_1540_itm = return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      | or_38_cse;
  assign return_extract_17_and_3_cse = run_wen & (~(or_dcpl_570 | or_dcpl_697 | or_dcpl_694
      | or_dcpl_628 | or_dcpl_693));
  assign return_add_generic_AC_RND_CONV_false_1_op_bigger_mux_4_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_326);
  assign return_add_generic_AC_RND_CONV_false_1_op_bigger_mux_5_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_266);
  assign return_add_generic_AC_RND_CONV_false_10_exp_mux1h_8_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1,
      (stage_PE_1_x_im_d_sva[52]), and_dcpl_326);
  assign return_add_generic_AC_RND_CONV_false_10_exp_mux1h_11_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1,
      (stage_PE_1_x_im_d_sva[52]), and_dcpl_266);
  assign return_add_generic_AC_RND_CONV_false_10_exp_and_6_cse = (~ return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp)
      & (fsm_output[37]);
  assign return_add_generic_AC_RND_CONV_false_10_exp_and_7_cse = return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp
      & (fsm_output[37]);
  assign return_add_generic_AC_RND_CONV_false_11_exp_and_2_cse = (~ and_dcpl_261)
      & (fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_11_exp_and_3_cse = and_dcpl_261 & (fsm_output[16]);
  assign return_extract_1_exception_or_cse = (fsm_output[17]) | (fsm_output[20])
      | (fsm_output[44]);
  assign xor_cse = (out_f_d_rsci_q_d[63]) ^ (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[6]);
  assign xor_2_cse = (out_f_d_rsci_q_d[63]) ^ (stage_PE_1_x_im_d_sva[63]);
  assign xor_3_cse = (in_f_d_rsci_q_d[63]) ^ (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[6]);
  assign xor_4_cse = (in_f_d_rsci_q_d[63]) ^ (stage_PE_1_x_im_d_sva[63]);
  assign return_add_generic_AC_RND_CONV_false_11_and_3_cse = (~ xor_cse) & (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_11_and_4_cse = xor_cse & (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_11_and_5_cse = (~ xor_2_cse) & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_11_and_6_cse = xor_2_cse & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_11_and_15_cse = (~ xor_4_cse) & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_11_and_16_cse = xor_4_cse & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_11_and_13_cse = (~ xor_3_cse) & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_11_and_14_cse = xor_3_cse & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_22_op1_mu_and_cse = run_wen & (~(or_dcpl_610
      | or_dcpl_607 | (fsm_output[33]) | or_dcpl_500 | or_dcpl_697 | or_dcpl_587
      | or_dcpl_840 | or_dcpl_401));
  assign nl_return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl = ({1'b1 ,
      (out_f_d_rsci_q_d[51:0])}) + conv_u2u_52_53(~ (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[51:0]))
      + 53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl[52:0];
  assign return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_and_1_cse
      = (readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_2_ma1_lt_ma2_acc_2_nl))
      & return_add_generic_AC_RND_CONV_false_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_and_1_cse
      | (z_out_24[11]);
  assign nl_return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl = ({1'b1
      , (in_f_d_rsci_q_d[51:0])}) + conv_u2u_52_53(~ (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[51:0]))
      + 53'b00000000000000000000000000000000000000000000000000001;
  assign return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl[52:0];
  assign return_add_generic_AC_RND_CONV_false_13_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_13_op1_smaller_oelse_and_1_itm
      = (readslicef_53_1_52(return_add_generic_AC_RND_CONV_false_15_ma1_lt_ma2_acc_2_nl))
      & return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_13_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_13_op1_smaller_oelse_and_1_itm
      | (z_out_24[11]);
  assign return_add_generic_AC_RND_CONV_false_11_and_24_m1c = or_dcpl_863 & (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_11_and_28_m1c = or_dcpl_876 & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_11_and_23_cse = (~ or_dcpl_863) & (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_11_and_31_cse = (~ return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse)
      & return_add_generic_AC_RND_CONV_false_11_and_24_m1c;
  assign return_add_generic_AC_RND_CONV_false_11_and_32_cse = return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse
      & return_add_generic_AC_RND_CONV_false_11_and_24_m1c;
  assign return_add_generic_AC_RND_CONV_false_10_r_zero_and_cse = run_wen & (~(or_dcpl_465
      | (fsm_output[45]) | (fsm_output[42]) | or_dcpl_749 | or_dcpl_461 | (fsm_output[38])
      | (fsm_output[34]) | or_dcpl_552 | or_dcpl_418 | (fsm_output[19]) | (fsm_output[17])));
  assign return_add_generic_AC_RND_CONV_false_10_or_cse = (fsm_output[19]) | (fsm_output[42])
      | (fsm_output[45]);
  assign return_add_generic_AC_RND_CONV_false_22_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_22_op1_smaller_oelse_and_cse
      = z_out_33_52 & return_add_generic_AC_RND_CONV_false_22_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_22_op1_smaller_return_add_generic_AC_RND_CONV_false_22_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_22_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_22_op1_smaller_oelse_and_cse
      | (z_out_23[11]);
  assign and_494_m1c = or_dcpl_876 & inverse_lpi_1_dfm_1;
  assign return_extract_26_exception_or_3_cse = (fsm_output[8]) | (fsm_output[33]);
  assign and_491_tmp = or_dcpl_911 & inverse_lpi_1_dfm_1;
  assign and_497_tmp = or_dcpl_913 & inverse_lpi_1_dfm_1;
  assign return_extract_26_exception_and_5_m1c = and_491_tmp & (fsm_output[7]);
  assign return_extract_26_exception_and_7_m1c = or_dcpl_912 & (fsm_output[18]);
  assign return_extract_26_exception_and_10_m1c = and_497_tmp & (fsm_output[32]);
  assign return_extract_26_exception_and_12_m1c = or_dcpl_914 & (fsm_output[41]);
  assign return_extract_26_exception_and_6_cse = (~ or_dcpl_912) & (fsm_output[18]);
  assign return_extract_26_exception_and_11_cse = (~ or_dcpl_914) & (fsm_output[41]);
  assign return_extract_26_exception_and_17_cse = (~ return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse)
      & return_extract_26_exception_and_7_m1c;
  assign return_extract_26_exception_and_18_cse = return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse
      & return_extract_26_exception_and_7_m1c;
  assign return_extract_26_exception_and_21_cse = (~ return_add_generic_AC_RND_CONV_false_22_op1_smaller_return_add_generic_AC_RND_CONV_false_22_op1_smaller_or_cse)
      & return_extract_26_exception_and_12_m1c;
  assign return_extract_26_exception_and_22_cse = return_add_generic_AC_RND_CONV_false_22_op1_smaller_return_add_generic_AC_RND_CONV_false_22_op1_smaller_or_cse
      & return_extract_26_exception_and_12_m1c;
  assign return_add_generic_AC_RND_CONV_false_23_op1_nan_and_cse = run_wen & (~(or_dcpl_937
      | or_dcpl_560 | or_dcpl_751 | or_dcpl_125 | or_dcpl_136 | or_dcpl_135 | or_dcpl_133));
  assign stage_PE_1_tmp_re_d_and_ssc = run_wen & ((inverse_lpi_1_dfm_1 & (~ or_dcpl_780))
      | stage_PE_1_tmp_re_d_1_sva_1_mx0c0 | (fsm_output[7]) | stage_PE_1_tmp_re_d_1_sva_1_mx0c4
      | (fsm_output[32]));
  assign return_add_generic_AC_RND_CONV_false_8_exp_and_ssc = run_wen & (~(return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
      | or_dcpl_101 | or_dcpl_558 | or_dcpl_159 | or_dcpl_694 | or_dcpl_713));
  assign return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_and_1_cse
      = z_out_34_52 & return_add_generic_AC_RND_CONV_false_1_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_and_1_cse
      | (z_out_25[11]);
  assign return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_and_cse
      = z_out_34_52 & return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_and_cse
      | (z_out_25[11]);
  assign return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_and_1_cse
      = z_out_34_52 & return_add_generic_AC_RND_CONV_false_14_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_and_1_cse
      | (z_out_25[11]);
  assign return_add_generic_AC_RND_CONV_false_12_and_2_m1c = or_dcpl_911 & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_12_and_6_m1c = or_dcpl_913 & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_10_op2_nan_and_cse = run_wen & (~(or_dcpl_662
      | or_dcpl_126 | (fsm_output[42]) | (fsm_output[10]) | or_dcpl_424 | or_dcpl_1015
      | or_dcpl_712));
  assign return_add_generic_AC_RND_CONV_false_2_not_4_nl = ~ (z_out_6[53]);
  assign return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_and_5_cse
      = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000, (z_out_6[51:0]),
      return_add_generic_AC_RND_CONV_false_2_not_4_nl);
  assign return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse = (fsm_output[15])
      | (fsm_output[40]);
  assign nand_12_cse = ~(return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse
      & (~ (z_out_8[11])));
  assign return_add_generic_AC_RND_CONV_false_12_op_bigger_and_8_cse = (~ return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_tmp)
      & (fsm_output[12]);
  assign return_add_generic_AC_RND_CONV_false_12_op_bigger_and_9_cse = return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_tmp
      & (fsm_output[12]);
  assign return_add_generic_AC_RND_CONV_false_12_res_mant_and_ssc = run_wen & (~(or_dcpl_662
      | or_dcpl_961 | (fsm_output[24]) | (fsm_output[21])));
  assign return_add_generic_AC_RND_CONV_false_12_res_mant_or_cse = (fsm_output[20])
      | (fsm_output[45]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_31_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_22_op1_mu_52_lpi_3_dfm, and_dcpl_261);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_34_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_22_op1_mu_52_lpi_3_dfm, and_dcpl_265);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_34_cse = and_dcpl_260
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse = and_dcpl_264
      & (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_12_op_bigger_and_2_cse = run_wen &
      (~ or_tmp_857);
  assign return_add_generic_AC_RND_CONV_false_12_op_smaller_and_1_cse = run_wen &
      (~((fsm_output[44]) | (fsm_output[19])));
  assign return_add_generic_AC_RND_CONV_false_5_op_smaller_mux_1_cse = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[50]),
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_51_lpi_3_dfm_mx0, and_dcpl_326);
  assign return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_2_cse = MUX_s_1_2_2((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[50]),
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0, and_dcpl_266);
  assign return_add_generic_AC_RND_CONV_false_10_exp_mux_5_cse = MUX_s_1_2_2(drf_qr_lval_13_smx_0_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx0, and_dcpl_326);
  assign return_add_generic_AC_RND_CONV_false_13_mux_25_cse = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0, and_dcpl_266);
  assign return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_3_e_dif_qr_lpi_3_dfm_mx0_10_0[10:6]!=5'b00000)
      | ((z_out_24[11]) & (z_out_25[11]));
  assign return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_cse = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_3_e_dif_qr_lpi_3_dfm_mx0_10_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_1_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_2_if_acc_1_nl =  -z_out_29;
  assign return_mult_generic_AC_RND_CONV_false_2_if_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_2_if_acc_1_nl[12:0];
  assign return_mult_generic_AC_RND_CONV_false_2_if_acc_1_itm_12_1 = readslicef_13_1_12(return_mult_generic_AC_RND_CONV_false_2_if_acc_1_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_if_acc_1_nl =  -z_out_29;
  assign return_mult_generic_AC_RND_CONV_false_if_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_if_acc_1_nl[12:0];
  assign return_mult_generic_AC_RND_CONV_false_if_acc_1_itm_12_1 = readslicef_13_1_12(return_mult_generic_AC_RND_CONV_false_if_acc_1_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_1_if_acc_1_nl =  -z_out_29;
  assign return_mult_generic_AC_RND_CONV_false_1_if_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_1_if_acc_1_nl[12:0];
  assign return_mult_generic_AC_RND_CONV_false_1_if_acc_1_itm_12_1 = readslicef_13_1_12(return_mult_generic_AC_RND_CONV_false_1_if_acc_1_nl);
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0 = return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_mux_28);
  assign return_add_generic_AC_RND_CONV_false_1_mux_29_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva,
      return_add_generic_AC_RND_CONV_false_if_5_or_3, z_out_6[53]);
  assign return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs_mx1w0 = return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_1_mux_29_nl);
  assign return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0 = return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva
      | (~ return_add_generic_AC_RND_CONV_false_mux_28);
  assign nl_return_mult_generic_AC_RND_CONV_false_5_if_acc_1_nl =  -z_out_29;
  assign return_mult_generic_AC_RND_CONV_false_5_if_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_5_if_acc_1_nl[12:0];
  assign return_mult_generic_AC_RND_CONV_false_5_if_acc_1_itm_12_1 = readslicef_13_1_12(return_mult_generic_AC_RND_CONV_false_5_if_acc_1_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_3_if_acc_1_nl =  -z_out_29;
  assign return_mult_generic_AC_RND_CONV_false_3_if_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_3_if_acc_1_nl[12:0];
  assign return_mult_generic_AC_RND_CONV_false_3_if_acc_1_itm_12_1 = readslicef_13_1_12(return_mult_generic_AC_RND_CONV_false_3_if_acc_1_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_4_if_acc_1_nl =  -z_out_29;
  assign return_mult_generic_AC_RND_CONV_false_4_if_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_4_if_acc_1_nl[12:0];
  assign return_mult_generic_AC_RND_CONV_false_4_if_acc_1_itm_12_1 = readslicef_13_1_12(return_mult_generic_AC_RND_CONV_false_4_if_acc_1_nl);
  assign nl_return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl =  -(z_out_29[11:0]);
  assign return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl = nl_return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl[11:0];
  assign return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1 = readslicef_12_1_11(return_mult_generic_AC_RND_CONV_false_6_if_acc_1_nl);
  assign return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx1w0 = operator_11_true_return_24_sva
      | (~ return_add_generic_AC_RND_CONV_false_mux_28);
  assign operator_16_false_1_operator_16_false_1_and_mdf_sva_1 = (mode1_rsci_idat==16'b0000000000000001);
  assign operator_16_false_operator_16_false_nor_tmp = ~((mode1_rsci_idat!=16'b0000000000000000));
  assign mode_lpi_1_dfm_mx0w0 = operator_16_false_1_operator_16_false_1_and_mdf_sva_1
      | operator_16_false_operator_16_false_nor_tmp;
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_8 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_8,
      m_in_15_1_lpi_1_dfm_1_9, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_7 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_7,
      m_in_15_1_lpi_1_dfm_1_8, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_6 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_6,
      m_in_15_1_lpi_1_dfm_1_7, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_5 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_5,
      m_in_15_1_lpi_1_dfm_1_6, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_4 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_4,
      m_in_15_1_lpi_1_dfm_1_5, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_3 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_3,
      m_in_15_1_lpi_1_dfm_1_4, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_2 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_2,
      m_in_15_1_lpi_1_dfm_1_3, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_1 = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_1,
      m_in_15_1_lpi_1_dfm_1_2, mode_lpi_1_dfm);
  assign stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_0 = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_9,
      m_in_15_1_lpi_1_dfm_1_1, mode_lpi_1_dfm);
  assign stage_PE_1_and_1_tmp = mode_lpi_1_dfm & inverse_lpi_1_dfm_1;
  assign stage_PE_1_and_cse = (~ mode_lpi_1_dfm) & inverse_lpi_1_dfm_1;
  assign return_extract_3_m_zero_sva_mx1w0 = ~((out_f_d_rsci_q_d[51:0]!=52'b0000000000000000000000000000000000000000000000000000));
  assign BUTTERFLY_i_div_psp_sva_1 = div_9_u9_u16(BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2,
      {stage_PE_1_index_const_15_lpi_2_dfm , stage_PE_1_index_const_14_11_lpi_2_dfm_3
      , stage_PE_1_index_const_14_11_lpi_2_dfm_2 , stage_PE_1_index_const_14_11_lpi_2_dfm_1
      , stage_PE_1_index_const_14_11_lpi_2_dfm_0 , stage_PE_1_index_const_10_lpi_2_dfm
      , stage_PE_1_index_const_9_1_lpi_2_dfm_8 , stage_PE_1_index_const_9_1_lpi_2_dfm_7
      , stage_PE_1_index_const_9_1_lpi_2_dfm_6 , stage_PE_1_index_const_9_1_lpi_2_dfm_5
      , stage_PE_1_index_const_9_1_lpi_2_dfm_4 , stage_PE_1_index_const_9_1_lpi_2_dfm_3
      , stage_PE_1_index_const_9_1_lpi_2_dfm_2 , stage_PE_1_index_const_9_1_lpi_2_dfm_1
      , stage_PE_1_index_const_9_1_lpi_2_dfm_0 , stage_PE_1_index_const_0_lpi_2_dfm});
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (z_out_37[10:1]), return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1));
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_1_nl = ~(MUX_v_10_2_2(10'b0000000000,
      z_out_20, return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1));
  assign return_add_generic_AC_RND_CONV_false_4_mux_18_nl = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_nl,
      return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_1_nl, z_out_6[53]);
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_qr_10_1_lpi_3_dfm_1 = ~(MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_4_mux_18_nl,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_4_e_r_qelse_or_svs_1));
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_2_nl = ~((z_out_37[0])
      & return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1);
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nor_nl = ~((z_out_28[0])
      | (~ return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1));
  assign return_add_generic_AC_RND_CONV_false_4_mux_19_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nand_2_nl,
      return_add_generic_AC_RND_CONV_false_4_e_r_qelse_nor_nl, z_out_6[53]);
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1 = ~(return_add_generic_AC_RND_CONV_false_4_mux_19_nl
      | return_add_generic_AC_RND_CONV_false_4_e_r_qelse_or_svs_1);
  assign return_add_generic_AC_RND_CONV_false_2_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_23_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva | return_add_generic_AC_RND_CONV_false_2_r_nan_and_2;
  assign and_358_nl = (or_dcpl_203 | and_dcpl_166 | return_add_generic_AC_RND_CONV_false_14_op2_inf_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva | return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva)
      & inverse_lpi_1_dfm_1;
  assign and_366_nl = (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_2_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
      & or_dcpl_431 & (~ return_add_generic_AC_RND_CONV_false_23_op1_inf_sva) & (~(return_add_generic_AC_RND_CONV_false_23_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_inf_sva | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva))
      & and_dcpl_241;
  assign return_extract_15_return_extract_15_nor_cse_sva_mx1 = MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_2_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[51]), (stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_0[0]),
      {and_358_nl , and_366_nl , (~ inverse_lpi_1_dfm_1)});
  assign return_add_generic_AC_RND_CONV_false_6_r_sign_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm,
      (~ stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0), or_918_cse);
  assign return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_and_nl
      = (({return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm
      , return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm
      , return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm}) == ({return_add_generic_AC_RND_CONV_false_6_op2_mu_52_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_50_mx0 , return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_49_0_mx0
      , return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1})) & return_add_generic_AC_RND_CONV_false_6_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_6_mux_6_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_r_sign_mux_nl,
      return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_nor_2,
      return_add_generic_AC_RND_CONV_false_6_if_2_return_add_generic_AC_RND_CONV_false_6_if_2_and_nl);
  assign stage_d_mul_return_d_2_63_sva_1 = inverse_lpi_1_dfm_1 ^ return_add_generic_AC_RND_CONV_false_6_mux_6_nl;
  assign return_add_generic_AC_RND_CONV_false_15_r_nan_or_mx2w0 = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | (return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva & return_add_generic_AC_RND_CONV_false_11_do_sub_sva);
  assign and_367_nl = (or_dcpl_278 | and_dcpl_166 | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op1_inf_sva | return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva)
      & inverse_lpi_1_dfm_1;
  assign and_374_nl = (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_15_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
      & or_dcpl_431 & (~ return_add_generic_AC_RND_CONV_false_10_op2_nan_sva) & (~(return_add_generic_AC_RND_CONV_false_10_op2_inf_sva
      | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva | return_add_generic_AC_RND_CONV_false_10_op1_inf_sva))
      & and_dcpl_241;
  assign return_extract_15_return_extract_15_nor_cse_sva_mx2 = MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_15_r_nan_or_mx2w0,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[51]), (stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_0[0]),
      {and_367_nl , and_374_nl , (~ inverse_lpi_1_dfm_1)});
  assign return_add_generic_AC_RND_CONV_false_19_r_sign_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm,
      (~ stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0), or_920_cse);
  assign return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_and_nl
      = (({return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm
      , return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm , drf_qr_lval_13_smx_0_lpi_3_dfm})
      == ({return_add_generic_AC_RND_CONV_false_19_op2_mu_52_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50_mx0
      , return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0_mx0 ,
      return_add_generic_AC_RND_CONV_false_19_op2_mu_0_lpi_3_dfm_1})) & return_add_generic_AC_RND_CONV_false_19_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_19_mux_6_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_19_r_sign_mux_nl,
      return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_nor_2,
      return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_and_nl);
  assign stage_d_mul_return_d_5_63_sva_1 = inverse_lpi_1_dfm_1 ^ return_add_generic_AC_RND_CONV_false_19_mux_6_nl;
  assign return_add_generic_AC_RND_CONV_false_4_m_r_51_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_and_5_cse[51])
      & (~ all_same_out);
  assign return_add_generic_AC_RND_CONV_false_4_if_7_not_5_nl = ~ all_same_out;
  assign return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_and_5_cse[50:0]),
      return_add_generic_AC_RND_CONV_false_4_if_7_not_5_nl);
  assign return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_tmp
      = (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1!=11'b00000000000);
  assign return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp
      = (return_mult_generic_AC_RND_CONV_false_3_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w6!=11'b00000000000);
  assign nl_return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt = ({1'b1 ,
      (~ (O_1_out[61:52]))}) + conv_u2s_10_11(O_1_out_1[61:52]) + 11'b00000000001;
  assign return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt = nl_return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt[10:0];
  assign return_add_generic_AC_RND_CONV_false_4_e_dif_qif_acc_pmx_lpi_3_dfm_mx0_9_0
      = MUX_v_10_2_2((return_add_generic_AC_RND_CONV_false_4_e_dif_acc_tmp[9:0]),
      (return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt[9:0]), return_add_generic_AC_RND_CONV_false_4_e_dif_acc_tmp[10]);
  assign return_add_generic_AC_RND_CONV_false_17_op1_mu_52_lpi_3_dfm_1 = (O_1_out[51])
      | return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_or_tmp;
  assign stage_PE_1_gm_re_d_mux_cse = MUX_v_51_2_2((O_1_out[50:0]), (O_1_out[51:1]),
      return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_or_tmp);
  assign return_add_generic_AC_RND_CONV_false_17_op1_mu_0_lpi_3_dfm_1 = (O_1_out[0])
      & return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_or_tmp;
  assign stage_PE_1_gm_im_d_mux_cse = MUX_s_1_2_2(return_extract_9_return_extract_9_or_1_cse_sva_1,
      (O_1_out_1[51]), return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_if_1_return_add_generic_AC_RND_CONV_false_4_op2_normal_return_extract_9_nor_tmp);
  assign stage_PE_1_gm_im_d_mux_2_cse = MUX_v_51_2_2((O_1_out_1[51:1]), (O_1_out_1[50:0]),
      return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_if_1_return_add_generic_AC_RND_CONV_false_4_op2_normal_return_extract_9_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_17_op2_mu_0_lpi_3_dfm_1 = (O_1_out_1[0])
      & (~ return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_if_1_return_add_generic_AC_RND_CONV_false_4_op2_normal_return_extract_9_nor_tmp);
  assign drf_qr_lval_4_smx_9_0_lpi_3_dfm_mx0 = MUX_v_10_2_2((O_1_out_1[61:52]), (O_1_out[61:52]),
      and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_4_op_smaller_qr_0_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_17_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_17_op2_mu_0_lpi_3_dfm_1, and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_4_sticky_bit_and_cse = return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_6_cse
      & (~ (z_out_16[54]));
  assign return_add_generic_AC_RND_CONV_false_4_sticky_bit_and_52_cse = return_add_generic_AC_RND_CONV_false_4_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_16[2]));
  assign return_add_generic_AC_RND_CONV_false_4_res_mant_3_0_sva_1 = return_add_generic_AC_RND_CONV_false_4_sticky_bit_and_cse
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[50]) & (~ (z_out_16[53])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[49]) & (~ (z_out_16[52])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[48]) & (~ (z_out_16[51])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[47]) & (~ (z_out_16[50])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[46]) & (~ (z_out_16[49])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[45]) & (~ (z_out_16[48])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[44]) & (~ (z_out_16[47])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[43]) & (~ (z_out_16[46])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[42]) & (~ (z_out_16[45])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[41]) & (~ (z_out_16[44])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[40]) & (~ (z_out_16[43])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[39]) & (~ (z_out_16[42])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[38]) & (~ (z_out_16[41])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[37]) & (~ (z_out_16[40])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[36]) & (~ (z_out_16[39])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[35]) & (~ (z_out_16[38])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[34]) & (~ (z_out_16[37])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[33]) & (~ (z_out_16[36])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[32]) & (~ (z_out_16[35])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[31]) & (~ (z_out_16[34])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[30]) & (~ (z_out_16[33])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[29]) & (~ (z_out_16[32])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[28]) & (~ (z_out_16[31])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[27]) & (~ (z_out_16[30])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[26]) & (~ (z_out_16[29])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[25]) & (~ (z_out_16[28])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[24]) & (~ (z_out_16[27])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[23]) & (~ (z_out_16[26])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[22]) & (~ (z_out_16[25])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[21]) & (~ (z_out_16[24])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[20]) & (~ (z_out_16[23])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[19]) & (~ (z_out_16[22])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[18]) & (~ (z_out_16[21])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[17]) & (~ (z_out_16[20])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[16]) & (~ (z_out_16[19])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[15]) & (~ (z_out_16[18])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[14]) & (~ (z_out_16[17])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[13]) & (~ (z_out_16[16])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[12]) & (~ (z_out_16[15])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[11]) & (~ (z_out_16[14])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[10]) & (~ (z_out_16[13])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[9]) & (~ (z_out_16[12])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[8]) & (~ (z_out_16[11])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[7]) & (~ (z_out_16[10])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[6]) & (~ (z_out_16[9])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[5]) & (~ (z_out_16[8])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[4]) & (~ (z_out_16[7])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[3]) & (~ (z_out_16[6])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[2]) & (~ (z_out_16[5])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[1]) & (~ (z_out_16[4])))
      | ((return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse[0]) & (~ (z_out_16[3])))
      | return_add_generic_AC_RND_CONV_false_4_sticky_bit_and_52_cse;
  assign return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_if_1_return_add_generic_AC_RND_CONV_false_4_op2_normal_return_extract_9_nor_tmp
      = ~((O_1_out_1[61:52]!=10'b0000000000));
  assign nl_return_add_generic_AC_RND_CONV_false_4_acc_2_nl =  -(z_out_37[10:0]);
  assign return_add_generic_AC_RND_CONV_false_4_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_4_acc_2_nl[10:0];
  assign return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1 = readslicef_11_1_10(return_add_generic_AC_RND_CONV_false_4_acc_2_nl);
  assign return_add_generic_AC_RND_CONV_false_4_if_5_return_add_generic_AC_RND_CONV_false_4_if_5_nor_cse
      = ~((z_out_37[11:0]!=12'b000000000000));
  assign return_add_generic_AC_RND_CONV_false_4_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1
      | return_add_generic_AC_RND_CONV_false_4_if_5_return_add_generic_AC_RND_CONV_false_4_if_5_nor_cse;
  assign return_add_generic_AC_RND_CONV_false_4_mux_15_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1,
      return_add_generic_AC_RND_CONV_false_4_if_5_or_1_nl, z_out_6[53]);
  assign return_add_generic_AC_RND_CONV_false_4_e_r_qelse_or_svs_1 = all_same_out
      | (~ return_add_generic_AC_RND_CONV_false_4_mux_15_nl);
  assign return_add_generic_AC_RND_CONV_false_4_mux_10_itm = MUX_v_6_2_2((drf_qr_lval_4_smx_9_0_lpi_3_dfm_mx0[5:0]),
      rtn_out, return_add_generic_AC_RND_CONV_false_4_acc_2_itm_10_1);
  assign return_add_generic_AC_RND_CONV_false_17_do_sub_sva_1 = ~((O_1_out[63]) ^
      inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_4_e_dif_sat_or_2_nl = (return_add_generic_AC_RND_CONV_false_4_e_dif_qif_acc_pmx_lpi_3_dfm_mx0_9_0[9:6]!=4'b0000)
      | ((return_add_generic_AC_RND_CONV_false_18_e_dif_qif_acc_sdt[10]) & (return_add_generic_AC_RND_CONV_false_4_e_dif_acc_tmp[10]));
  assign return_add_generic_AC_RND_CONV_false_4_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_4_e_dif_qif_acc_pmx_lpi_3_dfm_mx0_9_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_4_e_dif_sat_or_2_nl);
  assign nl_BUTTERFLY_i_9_0_sva_1 = conv_u2u_9_10(BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2)
      + (z_out_21[9:0]);
  assign BUTTERFLY_i_9_0_sva_1 = nl_BUTTERFLY_i_9_0_sva_1[9:0];
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx1 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1,
      and_dcpl_258);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1,
      and_dcpl_259);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx5 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1,
      and_dcpl_262);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx6 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1,
      and_dcpl_263);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx1 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_op2_mu_52_lpi_3_dfm_1, drf_qr_lval_13_smx_0_lpi_3_dfm,
      and_dcpl_258);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx2 =
      MUX_s_1_2_2(drf_qr_lval_13_smx_0_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_op2_mu_52_lpi_3_dfm_1,
      and_dcpl_259);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx6 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_13_op1_mu_52_lpi_3_dfm_1,
      drf_qr_lval_13_smx_0_lpi_3_dfm, and_dcpl_262);
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx7 =
      MUX_s_1_2_2(drf_qr_lval_13_smx_0_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_13_op1_mu_52_lpi_3_dfm_1,
      and_dcpl_263);
  assign return_extract_9_return_extract_9_or_1_cse_sva_1 = (O_1_out_1[61:52]!=10'b0000000000);
  assign and_2331_cse = return_extract_13_m_zero_return_extract_13_m_zero_nor_tmp
      & return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_1_return_add_generic_AC_RND_CONV_false_6_op2_normal_return_extract_13_nor_tmp;
  assign and_411_nl = (~(operator_11_true_return_17_sva | operator_11_true_13_operator_11_true_13_and_tmp))
      & (~(return_extract_17_return_extract_17_nor_cse_sva & return_extract_17_m_zero_sva))
      & (~(and_2331_cse | return_mult_generic_AC_RND_CONV_false_1_exp_ovf_return_mult_generic_AC_RND_CONV_false_1_exp_ovf_or_tmp));
  assign drf_qr_lval_14_smx_0_lpi_3_dfm_mx1 = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_1_r_nan_sva_1,
      (z_out_6[51]), and_411_nl);
  assign and_2332_cse = return_extract_24_m_zero_sva & return_extract_15_return_extract_15_nor_cse_sva;
  assign and_415_nl = (~(operator_11_true_return_17_sva | operator_11_true_44_operator_11_true_44_and_tmp))
      & (~(return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp
      & return_extract_44_m_zero_return_extract_44_m_zero_nor_tmp)) & (~(and_2332_cse
      | return_mult_generic_AC_RND_CONV_false_3_exp_ovf_return_mult_generic_AC_RND_CONV_false_3_exp_ovf_or_tmp));
  assign drf_qr_lval_14_smx_0_lpi_3_dfm_mx3 = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_3_r_nan_sva_1,
      (z_out_6[51]), and_415_nl);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nand_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (z_out_37[10:1]), return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10_1));
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nand_1_nl = ~(MUX_v_10_2_2(10'b0000000000,
      z_out_20, return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10_1));
  assign return_add_generic_AC_RND_CONV_false_17_mux_18_nl = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nand_nl,
      return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nand_1_nl, z_out_6[53]);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qelse_qr_10_1_lpi_3_dfm_1 =
      ~(MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_17_mux_18_nl, 10'b1111111111,
      return_add_generic_AC_RND_CONV_false_17_e_r_qelse_or_svs_1));
  assign BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_tmp = (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2==9'b011111111);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nand_2_nl = ~((z_out_37[0])
      & return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10_1);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nor_nl = ~((z_out_28[0])
      | (~ return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10_1));
  assign return_add_generic_AC_RND_CONV_false_17_mux_19_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nand_2_nl,
      return_add_generic_AC_RND_CONV_false_17_e_r_qelse_nor_nl, z_out_6[53]);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm_1 = ~(return_add_generic_AC_RND_CONV_false_17_mux_19_nl
      | return_add_generic_AC_RND_CONV_false_17_e_r_qelse_or_svs_1);
  assign return_add_generic_AC_RND_CONV_false_9_if_2_return_add_generic_AC_RND_CONV_false_9_if_2_and_1_mx2w0
      = return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 & (stage_PE_1_x_re_d_sva[63]);
  assign return_add_generic_AC_RND_CONV_false_12_if_2_return_add_generic_AC_RND_CONV_false_12_if_2_nor_mx4w0
      = ~(return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva
      | (~ (stage_PE_1_x_im_d_sva[63])));
  assign return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_tmp
      = (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w3!=11'b00000000000);
  assign return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp
      = (return_mult_generic_AC_RND_CONV_false_4_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w2!=11'b00000000000);
  assign return_add_generic_AC_RND_CONV_false_7_if_2_return_add_generic_AC_RND_CONV_false_7_if_2_and_1_mx1w0
      = return_extract_15_return_extract_15_nor_cse_sva & return_add_generic_AC_RND_CONV_false_18_e_r_qr_0_lpi_3_dfm;
  assign return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_and_cse
      = z_out_35_52 & return_add_generic_AC_RND_CONV_false_7_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_7_op1_smaller_return_add_generic_AC_RND_CONV_false_7_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_and_cse
      | (z_out_25[11]);
  assign return_add_generic_AC_RND_CONV_false_7_r_sign_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_18_e_r_qr_0_lpi_3_dfm,
      return_extract_15_return_extract_15_nor_cse_sva, return_add_generic_AC_RND_CONV_false_7_op1_smaller_return_add_generic_AC_RND_CONV_false_7_op1_smaller_or_cse);
  assign nand_108_nl = ~(return_add_generic_AC_RND_CONV_false_7_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm , return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm
      , return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_49_0 , return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1})));
  assign return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_if_2_return_add_generic_AC_RND_CONV_false_7_if_2_and_1_mx1w0,
      return_add_generic_AC_RND_CONV_false_7_r_sign_mux_1_nl, nand_108_nl);
  assign return_add_generic_AC_RND_CONV_false_8_if_2_return_add_generic_AC_RND_CONV_false_8_if_2_and_1_mx2w0
      = return_extract_15_return_extract_15_nor_cse_sva & return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm;
  assign return_add_generic_AC_RND_CONV_false_20_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_20_op1_smaller_oelse_and_cse
      = z_out_31_52 & return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_20_op1_smaller_return_add_generic_AC_RND_CONV_false_20_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_20_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_20_op1_smaller_oelse_and_cse
      | (z_out_26[11]);
  assign return_add_generic_AC_RND_CONV_false_20_r_sign_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm,
      return_extract_15_return_extract_15_nor_cse_sva, return_add_generic_AC_RND_CONV_false_20_op1_smaller_return_add_generic_AC_RND_CONV_false_20_op1_smaller_or_cse);
  assign nand_109_nl = ~((({return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm
      , return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm , return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_49_0
      , return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1
      , return_add_generic_AC_RND_CONV_false_20_op2_mu_1_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_20_op2_mu_1_50_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_20_op2_mu_1_0_lpi_3_dfm_1})) & return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp);
  assign return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_if_2_return_add_generic_AC_RND_CONV_false_8_if_2_and_1_mx2w0,
      return_add_generic_AC_RND_CONV_false_20_r_sign_mux_1_nl, nand_109_nl);
  assign return_add_generic_AC_RND_CONV_false_2_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_2_e_dif_qr_lpi_3_dfm_mx0_10_0[10:6]!=5'b00000)
      | ((z_out_23[11]) & (z_out_24[11]));
  assign return_add_generic_AC_RND_CONV_false_2_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_2_e_dif_qr_lpi_3_dfm_mx0_10_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_2_e_dif_sat_or_1_nl);
  assign return_mult_generic_AC_RND_CONV_false_1_oelse_3_return_mult_generic_AC_RND_CONV_false_1_if_3_nor_nl
      = ~((~ return_mult_generic_AC_RND_CONV_false_1_zero_m_return_mult_generic_AC_RND_CONV_false_1_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_1_r_zero_return_mult_generic_AC_RND_CONV_false_1_r_zero_nor_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_1_lor_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (z_out_6[50:0]), return_mult_generic_AC_RND_CONV_false_1_oelse_3_return_mult_generic_AC_RND_CONV_false_1_if_3_nor_nl);
  assign return_mult_generic_AC_RND_CONV_false_3_oelse_3_return_mult_generic_AC_RND_CONV_false_3_if_3_nor_nl
      = ~((~ return_mult_generic_AC_RND_CONV_false_3_zero_m_return_mult_generic_AC_RND_CONV_false_3_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_3_r_zero_return_mult_generic_AC_RND_CONV_false_3_r_zero_nor_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_3_lor_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (z_out_6[50:0]), return_mult_generic_AC_RND_CONV_false_3_oelse_3_return_mult_generic_AC_RND_CONV_false_3_if_3_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx1 = MUX_v_51_2_2((out_f_d_rsci_q_d[50:0]),
      (out_f_d_rsci_q_d[51:1]), return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2 = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx1,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm, and_dcpl_258);
  assign return_mult_generic_AC_RND_CONV_false_oelse_3_return_mult_generic_AC_RND_CONV_false_if_3_nor_nl
      = ~((~ return_mult_generic_AC_RND_CONV_false_zero_m_return_mult_generic_AC_RND_CONV_false_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_r_zero_return_mult_generic_AC_RND_CONV_false_r_zero_nor_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_lor_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (z_out_6[50:0]), return_mult_generic_AC_RND_CONV_false_oelse_3_return_mult_generic_AC_RND_CONV_false_if_3_nor_nl);
  assign return_mult_generic_AC_RND_CONV_false_4_oelse_3_return_mult_generic_AC_RND_CONV_false_4_if_3_nor_nl
      = ~((~ return_mult_generic_AC_RND_CONV_false_4_zero_m_return_mult_generic_AC_RND_CONV_false_4_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_4_r_zero_return_mult_generic_AC_RND_CONV_false_4_r_zero_nor_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_4_lor_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (z_out_6[50:0]), return_mult_generic_AC_RND_CONV_false_4_oelse_3_return_mult_generic_AC_RND_CONV_false_4_if_3_nor_nl);
  assign and_1589_cse = and_dcpl_348 & (fsm_output[37]);
  assign or_1670_ssc = return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
      | or_dcpl_423 | or_dcpl_716 | or_dcpl_136 | (fsm_output[9]) | (fsm_output[36])
      | or_dcpl_793 | and_1589_cse | (and_dcpl_349 & (fsm_output[12]));
  assign and_468_cse = return_add_generic_AC_RND_CONV_false_6_e1_eq_e2_equal_tmp
      & z_out_32_52;
  assign or_918_cse = and_468_cse | (z_out_24[11]);
  assign or_1673_ssc = or_918_cse & (fsm_output[12]);
  assign and_470_cse = z_out_32_52 & return_add_generic_AC_RND_CONV_false_19_e1_eq_e2_equal_tmp;
  assign or_920_cse = and_470_cse | (z_out_24[11]);
  assign or_1678_ssc = or_920_cse & (fsm_output[37]);
  assign return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp
      = (out_f_d_rsci_q_d[62:52]!=11'b00000000000);
  assign operator_11_true_24_operator_11_true_24_and_tmp = (out_f_d_rsci_q_d[62:52]==11'b11111111111);
  assign operator_11_true_33_operator_11_true_33_and_tmp = (in_f_d_rsci_q_d[62:52]==11'b11111111111);
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_5_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (z_out_37[10:1]), return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1));
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_7_nl = ~(MUX_v_10_2_2(10'b0000000000,
      z_out_20, return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1));
  assign return_add_generic_AC_RND_CONV_false_5_mux_25_nl = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_5_nl,
      return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_7_nl, z_out_6[53]);
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qelse_qr_10_1_lpi_3_dfm_1 = ~(MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_5_mux_25_nl,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_svs_1));
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_3_nl = ~((z_out_37[0])
      & return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1);
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nor_1_nl = ~((z_out_28[0])
      | (~ return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1));
  assign return_add_generic_AC_RND_CONV_false_5_mux_23_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nand_3_nl,
      return_add_generic_AC_RND_CONV_false_5_e_r_qelse_nor_1_nl, z_out_6[53]);
  assign return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1 = ~(return_add_generic_AC_RND_CONV_false_5_mux_23_nl
      | return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_svs_1);
  assign operator_11_true_return_17_sva_mx0w0 = (return_add_generic_AC_RND_CONV_false_5_e_r_qelse_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_5_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm
      & (~ (z_out_16[54]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[50])
      & (~ (z_out_16[53]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49])
      & (~ (z_out_16[52]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[48])
      & (~ (z_out_16[51]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[47])
      & (~ (z_out_16[50]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[46])
      & (~ (z_out_16[49]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[45])
      & (~ (z_out_16[48]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[44])
      & (~ (z_out_16[47]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[43])
      & (~ (z_out_16[46]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[42])
      & (~ (z_out_16[45]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[41])
      & (~ (z_out_16[44]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[40])
      & (~ (z_out_16[43]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[39])
      & (~ (z_out_16[42]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[38])
      & (~ (z_out_16[41]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[37])
      & (~ (z_out_16[40]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[36])
      & (~ (z_out_16[39]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[35])
      & (~ (z_out_16[38]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[34])
      & (~ (z_out_16[37]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[33])
      & (~ (z_out_16[36]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[32])
      & (~ (z_out_16[35]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[31])
      & (~ (z_out_16[34]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[30])
      & (~ (z_out_16[33]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[29])
      & (~ (z_out_16[32]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[28])
      & (~ (z_out_16[31]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[27])
      & (~ (z_out_16[30]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[26])
      & (~ (z_out_16[29]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[25])
      & (~ (z_out_16[28]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[24])
      & (~ (z_out_16[27]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[23])
      & (~ (z_out_16[26]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[22])
      & (~ (z_out_16[25]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[21])
      & (~ (z_out_16[24]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[20])
      & (~ (z_out_16[23]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[19])
      & (~ (z_out_16[22]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[18])
      & (~ (z_out_16[21]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[17])
      & (~ (z_out_16[20]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[16])
      & (~ (z_out_16[19]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[15])
      & (~ (z_out_16[18]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[14])
      & (~ (z_out_16[17]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[13])
      & (~ (z_out_16[16]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[12])
      & (~ (z_out_16[15]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[11])
      & (~ (z_out_16[14]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[10])
      & (~ (z_out_16[13]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[9])
      & (~ (z_out_16[12]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[8])
      & (~ (z_out_16[11]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[7])
      & (~ (z_out_16[10]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[6])
      & (~ (z_out_16[9]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[5])
      & (~ (z_out_16[8]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[4])
      & (~ (z_out_16[7]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[3])
      & (~ (z_out_16[6]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[2])
      & (~ (z_out_16[5]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[1])
      & (~ (z_out_16[4]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[0])
      & (~ (z_out_16[3]))) | return_add_generic_AC_RND_CONV_false_5_sticky_bit_and_54;
  assign return_add_generic_AC_RND_CONV_false_5_if_5_or_2_nl = return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1
      | return_add_generic_AC_RND_CONV_false_4_if_5_return_add_generic_AC_RND_CONV_false_4_if_5_nor_cse;
  assign return_add_generic_AC_RND_CONV_false_5_mux_27_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1,
      return_add_generic_AC_RND_CONV_false_5_if_5_or_2_nl, z_out_6[53]);
  assign return_add_generic_AC_RND_CONV_false_18_e_r_qelse_or_svs_1 = all_same_out
      | (~ return_add_generic_AC_RND_CONV_false_5_mux_27_nl);
  assign return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm_mx1 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_260);
  assign return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm_mx4 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_20_op2_mu_1_0_lpi_3_dfm_1, and_dcpl_264);
  assign return_add_generic_AC_RND_CONV_false_op2_mu_52_lpi_3_dfm_1 = (out_f_d_rsci_q_d[51])
      | return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp;
  assign return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm_mx0w4 = (stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_1[0])
      & (~ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva);
  assign return_add_generic_AC_RND_CONV_false_13_op1_mu_52_lpi_3_dfm_1 = (in_f_d_rsci_q_d[51])
      | return_add_generic_AC_RND_CONV_false_13_return_add_generic_AC_RND_CONV_false_13_or_1_tmp;
  assign stage_d_mul_return_d_63_sva_1 = return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm
      ^ return_add_generic_AC_RND_CONV_false_17_mux_6_itm;
  assign stage_d_mul_return_d_4_63_sva_1 = stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0 ^
      return_add_generic_AC_RND_CONV_false_18_mux_itm;
  assign nl_return_add_generic_AC_RND_CONV_false_acc_2_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_1_acc_2_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_1_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_1_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_1_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_1_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_9_acc_2_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_9_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_9_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_9_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_9_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_10_acc_2_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_10_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_10_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_10_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_10_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_11_acc_2_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_11_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_11_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_11_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_12_acc_2_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_12_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_12_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_12_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_12_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_13_acc_2_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_13_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_13_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_13_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_13_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_14_acc_2_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_14_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_14_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_14_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_14_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_22_acc_2_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_22_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_22_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_22_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_22_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_23_acc_2_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_23_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_23_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_23_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_24_acc_2_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_24_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_24_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_24_acc_2_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_25_acc_2_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_25_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_25_acc_2_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_25_acc_2_nl);
  assign drf_qr_lval_smx_lpi_3_dfm_mx0_10_5 = MUX_v_6_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_0[5:0]),
      (out_f_d_rsci_q_d[62:57]), and_dcpl_258);
  assign drf_qr_lval_smx_lpi_3_dfm_mx0_4_0 = MUX_v_5_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_1[56:52]),
      (out_f_d_rsci_q_d[56:52]), and_dcpl_258);
  assign return_add_generic_AC_RND_CONV_false_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_24,
      z_out_23, z_out_24[11]);
  assign return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1 = (out_f_d_rsci_q_d[0])
      & return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp;
  assign return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1 = (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[0])
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_e1_eq_e2_equal_tmp = (out_f_d_rsci_q_d[62:52])
      == ({(stage_PE_1_tmp_im_d_1_sva_1_rsp_0[5:0]) , (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[56:52])});
  assign return_add_generic_AC_RND_CONV_false_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx1
      & (~ (z_out_16[54]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[50])
      & (~ (z_out_16[53]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[49])
      & (~ (z_out_16[52]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[48])
      & (~ (z_out_16[51]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[47])
      & (~ (z_out_16[50]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[46])
      & (~ (z_out_16[49]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[45])
      & (~ (z_out_16[48]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[44])
      & (~ (z_out_16[47]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[43])
      & (~ (z_out_16[46]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[42])
      & (~ (z_out_16[45]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[41])
      & (~ (z_out_16[44]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[40])
      & (~ (z_out_16[43]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[39])
      & (~ (z_out_16[42]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[38])
      & (~ (z_out_16[41]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[37])
      & (~ (z_out_16[40]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[36])
      & (~ (z_out_16[39]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[35])
      & (~ (z_out_16[38]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[34])
      & (~ (z_out_16[37]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[33])
      & (~ (z_out_16[36]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[32])
      & (~ (z_out_16[35]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[31])
      & (~ (z_out_16[34]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[30])
      & (~ (z_out_16[33]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[29])
      & (~ (z_out_16[32]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[28])
      & (~ (z_out_16[31]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[27])
      & (~ (z_out_16[30]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[26])
      & (~ (z_out_16[29]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[25])
      & (~ (z_out_16[28]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[24])
      & (~ (z_out_16[27]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[23])
      & (~ (z_out_16[26]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[22])
      & (~ (z_out_16[25]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[21])
      & (~ (z_out_16[24]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[20])
      & (~ (z_out_16[23]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[19])
      & (~ (z_out_16[22]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[18])
      & (~ (z_out_16[21]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[17])
      & (~ (z_out_16[20]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[16])
      & (~ (z_out_16[19]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[15])
      & (~ (z_out_16[18]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[14])
      & (~ (z_out_16[17]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[13])
      & (~ (z_out_16[16]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[12])
      & (~ (z_out_16[15]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[11])
      & (~ (z_out_16[14]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[10])
      & (~ (z_out_16[13]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[9])
      & (~ (z_out_16[12]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[8])
      & (~ (z_out_16[11]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[7])
      & (~ (z_out_16[10]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[6])
      & (~ (z_out_16[9]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[5])
      & (~ (z_out_16[8]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[4])
      & (~ (z_out_16[7]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[3])
      & (~ (z_out_16[6]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[2])
      & (~ (z_out_16[5]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[1])
      & (~ (z_out_16[4]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[0])
      & (~ (z_out_16[3]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx1
      & (~ (z_out_16[2])));
  assign return_add_generic_AC_RND_CONV_false_2_e_dif_qr_lpi_3_dfm_mx0_10_0 = MUX_v_11_2_2((z_out_24[10:0]),
      (z_out_23[10:0]), z_out_24[11]);
  assign return_add_generic_AC_RND_CONV_false_2_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx1
      & (~ (z_out_17[54]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[50])
      & (~ (z_out_17[53]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[49])
      & (~ (z_out_17[52]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[48])
      & (~ (z_out_17[51]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[47])
      & (~ (z_out_17[50]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[46])
      & (~ (z_out_17[49]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[45])
      & (~ (z_out_17[48]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[44])
      & (~ (z_out_17[47]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[43])
      & (~ (z_out_17[46]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[42])
      & (~ (z_out_17[45]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[41])
      & (~ (z_out_17[44]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[40])
      & (~ (z_out_17[43]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[39])
      & (~ (z_out_17[42]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[38])
      & (~ (z_out_17[41]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[37])
      & (~ (z_out_17[40]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[36])
      & (~ (z_out_17[39]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[35])
      & (~ (z_out_17[38]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[34])
      & (~ (z_out_17[37]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[33])
      & (~ (z_out_17[36]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[32])
      & (~ (z_out_17[35]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[31])
      & (~ (z_out_17[34]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[30])
      & (~ (z_out_17[33]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[29])
      & (~ (z_out_17[32]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[28])
      & (~ (z_out_17[31]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[27])
      & (~ (z_out_17[30]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[26])
      & (~ (z_out_17[29]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[25])
      & (~ (z_out_17[28]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[24])
      & (~ (z_out_17[27]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[23])
      & (~ (z_out_17[26]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[22])
      & (~ (z_out_17[25]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[21])
      & (~ (z_out_17[24]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[20])
      & (~ (z_out_17[23]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[19])
      & (~ (z_out_17[22]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[18])
      & (~ (z_out_17[21]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[17])
      & (~ (z_out_17[20]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[16])
      & (~ (z_out_17[19]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[15])
      & (~ (z_out_17[18]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[14])
      & (~ (z_out_17[17]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[13])
      & (~ (z_out_17[16]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[12])
      & (~ (z_out_17[15]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[11])
      & (~ (z_out_17[14]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[10])
      & (~ (z_out_17[13]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[9])
      & (~ (z_out_17[12]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[8])
      & (~ (z_out_17[11]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[7])
      & (~ (z_out_17[10]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[6])
      & (~ (z_out_17[9]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[5])
      & (~ (z_out_17[8]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[4])
      & (~ (z_out_17[7]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[3])
      & (~ (z_out_17[6]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[2])
      & (~ (z_out_17[5]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[1])
      & (~ (z_out_17[4]))) | ((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx2[0])
      & (~ (z_out_17[3]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx1
      & (~ (z_out_17[2])));
  assign return_add_generic_AC_RND_CONV_false_mux_26_itm_4_0 = MUX_v_5_2_2(drf_qr_lval_smx_lpi_3_dfm_mx0_4_0,
      (rtn_out[4:0]), return_add_generic_AC_RND_CONV_false_acc_2_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_e_dif_sat_or_cse = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_e_dif_sat_or_1_nl);
  assign and_2333_cse = return_extract_12_m_zero_return_extract_12_m_zero_nor_tmp
      & return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp;
  assign and_460_nl = (~(operator_11_true_return_15_sva | return_mult_generic_AC_RND_CONV_false_exp_ovf_return_mult_generic_AC_RND_CONV_false_exp_ovf_or_tmp))
      & (~(return_extract_15_return_extract_15_nor_cse_sva & return_extract_15_m_zero_sva))
      & (~(and_2333_cse | operator_11_true_12_operator_11_true_12_and_tmp));
  assign return_add_generic_AC_RND_CONV_false_11_mux_2_itm_mx3 = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_r_nan_sva_1,
      (z_out_6[51]), and_460_nl);
  assign and_464_nl = (~(return_extract_17_return_extract_17_nor_cse_sva & return_extract_1_m_zero_sva))
      & (~(return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_tmp
      & return_extract_45_m_zero_return_extract_45_m_zero_nor_tmp)) & (~(return_mult_generic_AC_RND_CONV_false_4_exp_ovf_return_mult_generic_AC_RND_CONV_false_4_exp_ovf_or_tmp
      | operator_11_true_45_operator_11_true_45_and_tmp | operator_11_true_return_24_sva));
  assign return_add_generic_AC_RND_CONV_false_11_mux_2_itm_mx9 = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_4_r_nan_sva_1,
      (z_out_6[51]), and_464_nl);
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w3_10_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_2_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_2_exception_sva_1);
  assign or_265_nl = or_dcpl_203 | or_dcpl_199 | and_dcpl_166;
  assign return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs, or_265_nl);
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w3_0 = (return_add_generic_AC_RND_CONV_false_6_mux_35
      & (~ return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_nl)) | return_add_generic_AC_RND_CONV_false_2_exception_sva_1;
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w9_10_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_2_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_15_exception_sva_1);
  assign or_340_nl = or_dcpl_278 | or_dcpl_275 | and_dcpl_166;
  assign return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_2_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs, or_340_nl);
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w9_0 = (return_add_generic_AC_RND_CONV_false_6_mux_35
      & (~ return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_2_nl)) | return_add_generic_AC_RND_CONV_false_15_exception_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_1_else_2_else_else_mux_nl = MUX_v_11_2_2((return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[10:0]),
      (z_out_36[10:0]), return_mult_generic_AC_RND_CONV_false_1_e_incr_lpi_3_dfm_2);
  assign return_mult_generic_AC_RND_CONV_false_1_else_2_else_return_mult_generic_AC_RND_CONV_false_1_else_2_else_and_nl
      = MUX_v_11_2_2(11'b00000000000, return_mult_generic_AC_RND_CONV_false_1_else_2_else_else_mux_nl,
      return_mult_generic_AC_RND_CONV_false_1_zero_m_return_mult_generic_AC_RND_CONV_false_1_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_1_r_zero_return_mult_generic_AC_RND_CONV_false_1_r_zero_nor_mdf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w3
      = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_1_else_2_else_return_mult_generic_AC_RND_CONV_false_1_else_2_else_and_nl,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_1_lor_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_3_else_2_else_else_mux_nl = MUX_v_11_2_2((return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[10:0]),
      (z_out_36[10:0]), return_mult_generic_AC_RND_CONV_false_3_e_incr_lpi_3_dfm_2);
  assign return_mult_generic_AC_RND_CONV_false_3_else_2_else_return_mult_generic_AC_RND_CONV_false_3_else_2_else_and_nl
      = MUX_v_11_2_2(11'b00000000000, return_mult_generic_AC_RND_CONV_false_3_else_2_else_else_mux_nl,
      return_mult_generic_AC_RND_CONV_false_3_zero_m_return_mult_generic_AC_RND_CONV_false_3_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_3_r_zero_return_mult_generic_AC_RND_CONV_false_3_r_zero_nor_mdf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_3_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w6
      = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_3_else_2_else_return_mult_generic_AC_RND_CONV_false_3_else_2_else_and_nl,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_3_lor_lpi_3_dfm_1);
  assign and_1615_cse = return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse
      & (fsm_output[7]);
  assign and_1626_cse = return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse
      & (fsm_output[32]);
  assign drf_qr_lval_1_smx_lpi_3_dfm_mx1 = MUX_v_11_2_2((out_f_d_rsci_q_d[62:52]),
      (stage_PE_1_x_im_d_sva[62:52]), and_dcpl_259);
  assign return_add_generic_AC_RND_CONV_false_11_if_2_return_add_generic_AC_RND_CONV_false_11_if_2_nor_mx2w0
      = ~(return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 | (~ (stage_PE_1_x_re_d_sva[63])));
  assign return_add_generic_AC_RND_CONV_false_10_if_2_return_add_generic_AC_RND_CONV_false_10_if_2_and_1_mx5w0
      = return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva
      & (stage_PE_1_x_im_d_sva[63]);
  assign return_add_generic_AC_RND_CONV_false_6_do_sub_sva_1 = ~(return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm
      ^ stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0);
  assign return_add_generic_AC_RND_CONV_false_13_return_add_generic_AC_RND_CONV_false_13_or_1_tmp
      = (in_f_d_rsci_q_d[62:52]!=11'b00000000000);
  assign return_add_generic_AC_RND_CONV_false_1_op1_nan_sva_mx3w0 = operator_11_true_return_1_sva
      & (~ return_extract_1_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_9_op2_nan_sva_mx7w0 = operator_11_true_return_1_sva
      & (~ return_extract_15_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_9_op1_nan_sva_1 = operator_11_true_return_24_sva
      & (~ return_extract_24_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_9_op1_inf_sva_1 = operator_11_true_return_24_sva
      & return_extract_24_m_zero_sva;
  assign return_extract_2_and_1_tmp = operator_11_true_return_1_sva & return_extract_1_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_2_r_nan_and_2 = return_add_generic_AC_RND_CONV_false_23_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_14_op2_inf_sva & return_add_generic_AC_RND_CONV_false_11_do_sub_sva;
  assign nl_operator_33_true_1_acc_nl = conv_s2u_11_12(z_out_1[11:1]) + 12'b000000000001;
  assign operator_33_true_1_acc_nl = nl_operator_33_true_1_acc_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_5_cse
      = MUX_v_12_2_2(12'b000000000000, operator_33_true_1_acc_nl, return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva);
  assign return_add_generic_AC_RND_CONV_false_if_5_or_nl = return_add_generic_AC_RND_CONV_false_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_mux_16_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_exception_sva_1 = return_add_generic_AC_RND_CONV_false_9_op1_inf_sva_1
      | return_extract_2_and_1_tmp | return_add_generic_AC_RND_CONV_false_9_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_1_op1_nan_sva_mx3w0 | return_add_generic_AC_RND_CONV_false_mux_16_nl;
  assign return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_or_2_cse
      = (z_out_1[0]) | (~ return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva);
  assign return_add_generic_AC_RND_CONV_false_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_10_op2_nan_sva_1 = operator_11_true_return_15_sva
      & (~ return_extract_17_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_9_op2_inf_sva_1 = operator_11_true_return_1_sva
      & return_extract_15_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_10_op2_inf_sva_1 = operator_11_true_return_15_sva
      & return_extract_17_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_1_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_25,
      z_out_24, z_out_25[11]);
  assign return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1 = (stage_PE_1_x_im_d_sva[0])
      & return_add_generic_AC_RND_CONV_false_10_unequal_tmp;
  assign return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0
      = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx1, and_dcpl_259);
  assign return_add_generic_AC_RND_CONV_false_1_e1_eq_e2_equal_tmp = (stage_PE_1_x_im_d_sva[62:52])
      == (out_f_d_rsci_q_d[62:52]);
  assign return_add_generic_AC_RND_CONV_false_1_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx2
      & (~ (z_out_16[54]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_16[53]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_16[52]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_16[51]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_16[50]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_16[49]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_16[48]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_16[47]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_16[46]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_16[45]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_16[44]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_16[43]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_16[42]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_16[41]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_16[40]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_16[39]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_16[38]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_16[37]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_16[36]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_16[35]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_16[34]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_16[33]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_16[32]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_16[31]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_16[30]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_16[29]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_16[28]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_16[27]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_16[26]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_16[25]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_16[24]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_16[23]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_16[22]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_16[21]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_16[20]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_16[19]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_16[18]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_16[17]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_16[16]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_16[15]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_16[14]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_16[13]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_16[12]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_16[11]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_16[10]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_16[9]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_16[8]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_16[7]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_16[6]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_16[5]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_16[4]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_16[3]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2
      & (~ (z_out_16[2])));
  assign return_add_generic_AC_RND_CONV_false_3_e_dif_qr_lpi_3_dfm_mx0_10_0 = MUX_v_11_2_2((z_out_25[10:0]),
      (z_out_24[10:0]), z_out_25[11]);
  assign return_add_generic_AC_RND_CONV_false_3_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx2
      & (~ (z_out_17[54]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_17[53]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_17[52]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_17[51]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_17[50]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_17[49]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_17[48]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_17[47]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_17[46]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_17[45]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_17[44]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_17[43]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_17[42]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_17[41]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_17[40]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_17[39]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_17[38]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_17[37]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_17[36]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_17[35]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_17[34]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_17[33]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_17[32]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_17[31]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_17[30]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_17[29]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_17[28]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_17[27]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_17[26]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_17[25]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_17[24]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_17[23]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_17[22]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_17[21]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_17[20]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_17[19]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_17[18]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_17[17]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_17[16]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_17[15]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_17[14]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_17[13]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_17[12]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_17[11]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_17[10]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_17[9]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_17[8]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_17[7]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_17[6]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_17[5]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_17[4]))) | ((return_add_generic_AC_RND_CONV_false_1_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_17[3]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2
      & (~ (z_out_17[2])));
  assign drf_qr_lval_11_smx_lpi_3_dfm_mx2 = MUX_v_11_2_2((in_f_d_rsci_q_d[62:52]),
      (stage_PE_1_x_im_d_sva[62:52]), and_dcpl_263);
  assign return_add_generic_AC_RND_CONV_false_1_if_5_or_nl = return_add_generic_AC_RND_CONV_false_1_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_1_mux_16_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_1_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_1_if_5_or_nl, z_out_6[53]);
  assign return_add_generic_AC_RND_CONV_false_1_exception_sva_1 = return_extract_2_and_1_tmp
      | return_add_generic_AC_RND_CONV_false_9_op1_inf_sva_1 | return_add_generic_AC_RND_CONV_false_1_op1_nan_sva_mx3w0
      | return_add_generic_AC_RND_CONV_false_9_op1_nan_sva_1 | return_add_generic_AC_RND_CONV_false_1_mux_16_nl;
  assign return_add_generic_AC_RND_CONV_false_1_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_1_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_1_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_1_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_1_mux_25_itm_4_0 = MUX_v_5_2_2(reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1,
      (return_add_generic_AC_RND_CONV_false_10_ls_sva[4:0]), return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva);
  assign return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1 = operator_11_true_44_operator_11_true_44_and_tmp
      & return_extract_44_m_zero_return_extract_44_m_zero_nor_tmp;
  assign return_add_generic_AC_RND_CONV_false_6_op2_nan_sva_1 = operator_11_true_13_operator_11_true_13_and_tmp
      & (~ return_extract_13_m_zero_return_extract_13_m_zero_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1 = operator_11_true_45_operator_11_true_45_and_tmp
      & (~ return_extract_45_m_zero_return_extract_45_m_zero_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 = operator_11_true_return_15_sva
      & (~ return_extract_1_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_22_op2_nan_sva_1 = operator_11_true_return_1_sva
      & (~ return_extract_24_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_6_op2_inf_sva_1 = operator_11_true_13_operator_11_true_13_and_tmp
      & return_extract_13_m_zero_return_extract_13_m_zero_nor_tmp;
  assign return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1 = operator_11_true_45_operator_11_true_45_and_tmp
      & return_extract_45_m_zero_return_extract_45_m_zero_nor_tmp;
  assign return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1 = operator_11_true_return_15_sva
      & return_extract_1_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_22_op2_inf_sva_1 = operator_11_true_return_1_sva
      & return_extract_24_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_2_if_7_return_add_generic_AC_RND_CONV_false_2_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_2_exception_sva_1 | return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva);
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0w0 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[50:0]),
      return_add_generic_AC_RND_CONV_false_2_if_7_return_add_generic_AC_RND_CONV_false_2_if_7_nor_nl);
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0 = MUX_v_51_2_2(stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_1,
      stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0w0, inverse_lpi_1_dfm_1);
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx1_50 = MUX_s_1_2_2((stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_1[50]),
      (stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0w0[50]), inverse_lpi_1_dfm_1);
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_5 = MUX_v_6_2_2((stage_PE_1_tmp_re_d_1_sva_1_63_57[5:0]),
      (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w3_10_1[9:4]), inverse_lpi_1_dfm_1);
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_4_1 = MUX_v_4_2_2((stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_0[5:2]),
      (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w3_10_1[3:0]), inverse_lpi_1_dfm_1);
  assign stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0 = MUX_s_1_2_2((stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_0[1]),
      stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w3_0, inverse_lpi_1_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_else_2_else_else_mux_nl = MUX_v_11_2_2((return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[10:0]),
      (z_out_36[10:0]), return_mult_generic_AC_RND_CONV_false_e_incr_lpi_3_dfm_2);
  assign return_mult_generic_AC_RND_CONV_false_else_2_else_return_mult_generic_AC_RND_CONV_false_else_2_else_and_nl
      = MUX_v_11_2_2(11'b00000000000, return_mult_generic_AC_RND_CONV_false_else_2_else_else_mux_nl,
      return_mult_generic_AC_RND_CONV_false_zero_m_return_mult_generic_AC_RND_CONV_false_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_r_zero_return_mult_generic_AC_RND_CONV_false_r_zero_nor_mdf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1 = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_else_2_else_return_mult_generic_AC_RND_CONV_false_else_2_else_and_nl,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_lor_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_6_op1_inf_sva_1 = operator_11_true_12_operator_11_true_12_and_tmp
      & return_extract_12_m_zero_return_extract_12_m_zero_nor_tmp;
  assign return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_1 = operator_11_true_12_operator_11_true_12_and_tmp
      & (~ return_extract_12_m_zero_return_extract_12_m_zero_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp
      = ~((stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_5!=6'b000000) | (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_4_1!=4'b0000)
      | stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0);
  assign return_add_generic_AC_RND_CONV_false_2_e_r_qelse_not_5_nl = ~ return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0;
  assign return_add_generic_AC_RND_CONV_false_2_e_r_qelse_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(10'b0000000000,
      z_out_9, return_add_generic_AC_RND_CONV_false_2_e_r_qelse_not_5_nl);
  assign return_add_generic_AC_RND_CONV_false_2_if_5_or_nl = return_add_generic_AC_RND_CONV_false_2_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_2_mux_10_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_2_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_2_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_2_exception_sva_1 = return_add_generic_AC_RND_CONV_false_23_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_inf_sva | return_add_generic_AC_RND_CONV_false_23_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva | return_add_generic_AC_RND_CONV_false_2_mux_10_nl;
  assign return_add_generic_AC_RND_CONV_false_2_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_2_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_mult_generic_AC_RND_CONV_false_if_1_aelse_return_mult_generic_AC_RND_CONV_false_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_if_acc_1_itm_12_1) | (z_out_18[105]);
  assign return_mult_generic_AC_RND_CONV_false_if_if_not_nl = ~ (z_out_29[12]);
  assign return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1 = MUX_v_12_2_2(12'b000000000000,
      (z_out_29[11:0]), return_mult_generic_AC_RND_CONV_false_if_if_not_nl);
  assign return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1 = ~((z_out_27[9:6]==4'b1111));
  assign return_mult_generic_AC_RND_CONV_false_e_incr_lpi_3_dfm_2 = ~((~(((z_out_18[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((z_out_18[51]) | return_mult_generic_AC_RND_CONV_false_if_1_aelse_return_mult_generic_AC_RND_CONV_false_if_1_aelse_or_2))
      | (z_out_18[105]))) | (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_zero_m_return_mult_generic_AC_RND_CONV_false_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_r_zero_return_mult_generic_AC_RND_CONV_false_r_zero_nor_mdf_sva_1
      = ~(and_2333_cse | return_mult_generic_AC_RND_CONV_false_op2_zero_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_r_nan_sva_1 = return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_1
      | (operator_11_true_return_15_sva & (~ return_extract_15_m_zero_sva)) | (return_add_generic_AC_RND_CONV_false_6_op1_inf_sva_1
      & return_mult_generic_AC_RND_CONV_false_op2_zero_sva_1) | (and_2333_cse & return_mult_generic_AC_RND_CONV_false_op2_inf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_exp_ovf_oif_aelse_nor_cse = ~((return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[11])
      | (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[0]));
  assign return_mult_generic_AC_RND_CONV_false_exp_ovf_return_mult_generic_AC_RND_CONV_false_exp_ovf_or_tmp
      = ((return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[10:1]==10'b1111111111)
      & return_mult_generic_AC_RND_CONV_false_exp_ovf_oif_aelse_nor_cse & return_mult_generic_AC_RND_CONV_false_e_incr_lpi_3_dfm_2)
      | (z_out_36[11]);
  assign return_mult_generic_AC_RND_CONV_false_lor_lpi_3_dfm_1 = return_add_generic_AC_RND_CONV_false_6_op1_inf_sva_1
      | return_mult_generic_AC_RND_CONV_false_op2_inf_sva_1 | return_mult_generic_AC_RND_CONV_false_exp_ovf_return_mult_generic_AC_RND_CONV_false_exp_ovf_or_tmp
      | return_mult_generic_AC_RND_CONV_false_r_nan_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_return_mult_generic_AC_RND_CONV_false_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_if_1_and_1_tmp_1 | (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_and_2_nl = return_mult_generic_AC_RND_CONV_false_if_1_and_1_tmp_1
      & (~ (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_res_bef_rnd_3_53_1_lpi_3_dfm_1 = MUX1HOT_v_53_3_2((z_out_18[104:52]),
      (z_out_18[103:51]), (z_out_42[53:1]), {return_mult_generic_AC_RND_CONV_false_return_mult_generic_AC_RND_CONV_false_nor_nl
      , return_mult_generic_AC_RND_CONV_false_and_2_nl , (z_out_27[12])});
  assign return_mult_generic_AC_RND_CONV_false_op2_inf_sva_1 = operator_11_true_return_15_sva
      & return_extract_15_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_op2_zero_sva_1 = return_extract_15_return_extract_15_nor_cse_sva
      & return_extract_15_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_1_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_if_acc_1_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva, z_out_27[12]);
  assign return_mult_generic_AC_RND_CONV_false_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_do_shift_left_1_mux_1_nl
      & (~ (z_out_18[105]));
  assign return_extract_12_return_extract_12_or_1_cse_sva_1 = (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_5!=6'b000000)
      | (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_4_1!=4'b0000) | stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0;
  assign return_extract_12_m_zero_return_extract_12_m_zero_nor_tmp = ~(return_extract_15_return_extract_15_nor_cse_sva_mx1
      | stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx1_50 | (stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0[49:0]!=50'b00000000000000000000000000000000000000000000000000));
  assign operator_11_true_12_operator_11_true_12_and_tmp = (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_5==6'b111111)
      & (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_4_1==4'b1111) & stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0;
  assign return_mult_generic_AC_RND_CONV_false_if_or_3_cse = (~ (z_out_27[5])) |
      return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_if_not_nl = ~ return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_if_nand_1_cse = ~(MUX_v_4_2_2(4'b0000,
      (z_out_27[4:1]), return_mult_generic_AC_RND_CONV_false_if_not_nl));
  assign return_mult_generic_AC_RND_CONV_false_if_or_cse = (~ (z_out_27[0])) | return_mult_generic_AC_RND_CONV_false_if_nor_ovfl_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_4_else_2_else_else_mux_nl = MUX_v_11_2_2((return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[10:0]),
      (z_out_36[10:0]), return_mult_generic_AC_RND_CONV_false_4_e_incr_lpi_3_dfm_2);
  assign return_mult_generic_AC_RND_CONV_false_4_else_2_else_return_mult_generic_AC_RND_CONV_false_4_else_2_else_and_nl
      = MUX_v_11_2_2(11'b00000000000, return_mult_generic_AC_RND_CONV_false_4_else_2_else_else_mux_nl,
      return_mult_generic_AC_RND_CONV_false_4_zero_m_return_mult_generic_AC_RND_CONV_false_4_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_4_r_zero_return_mult_generic_AC_RND_CONV_false_4_r_zero_nor_mdf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_4_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w2
      = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_4_else_2_else_return_mult_generic_AC_RND_CONV_false_4_else_2_else_and_nl,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_4_lor_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_and_cse
      = z_out_31_52 & return_add_generic_AC_RND_CONV_false_8_e1_eq_e2_equal_tmp;
  assign return_add_generic_AC_RND_CONV_false_8_op1_smaller_return_add_generic_AC_RND_CONV_false_8_op1_smaller_or_cse
      = return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_and_cse
      | (z_out_26[11]);
  assign return_add_generic_AC_RND_CONV_false_8_r_sign_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm,
      return_extract_15_return_extract_15_nor_cse_sva, return_add_generic_AC_RND_CONV_false_8_op1_smaller_return_add_generic_AC_RND_CONV_false_8_op1_smaller_or_cse);
  assign nand_114_nl = ~(return_add_generic_AC_RND_CONV_false_8_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm
      , return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm , return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1})));
  assign return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva_mx1
      = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_if_2_return_add_generic_AC_RND_CONV_false_8_if_2_and_1_mx2w0,
      return_add_generic_AC_RND_CONV_false_8_r_sign_mux_1_nl, nand_114_nl);
  assign return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp
      = ~((stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_5!=6'b000000) | (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_4_1!=4'b0000)
      | stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0);
  assign return_add_generic_AC_RND_CONV_false_21_r_sign_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_18_e_r_qr_0_lpi_3_dfm,
      return_extract_15_return_extract_15_nor_cse_sva, or_1144_cse);
  assign nand_115_nl = ~(return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm , drf_qr_lval_13_smx_0_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm , return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1})
      == ({return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_20_op2_mu_1_51_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_20_op2_mu_1_50_1_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_20_op2_mu_1_0_lpi_3_dfm_1})));
  assign return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva_mx2
      = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_if_2_return_add_generic_AC_RND_CONV_false_7_if_2_and_1_mx1w0,
      return_add_generic_AC_RND_CONV_false_21_r_sign_mux_1_nl, nand_115_nl);
  assign return_add_generic_AC_RND_CONV_false_19_op1_nan_sva_1 = operator_11_true_44_operator_11_true_44_and_tmp
      & (~ return_extract_44_m_zero_return_extract_44_m_zero_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_15_if_7_return_add_generic_AC_RND_CONV_false_15_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_15_exception_sva_1 | return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva);
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx0w3 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[50:0]),
      return_add_generic_AC_RND_CONV_false_15_if_7_return_add_generic_AC_RND_CONV_false_15_if_7_nor_nl);
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1 = MUX_v_51_2_2(stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_1,
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx0w3, inverse_lpi_1_dfm_1);
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx2_50 = MUX_s_1_2_2((stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_1[50]),
      (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx0w3[50]), inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_3_mux_16_mx0_4_0 = MUX_v_5_2_2(drf_qr_lval_11_smx_lpi_3_dfm_4_0,
      (return_add_generic_AC_RND_CONV_false_10_ls_sva[4:0]), return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1);
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0 = MUX_s_1_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_0[6]),
      return_add_generic_AC_RND_CONV_false_12_mux_itm, inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_3_if_7_return_add_generic_AC_RND_CONV_false_3_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_3_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0w0 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[50:0]),
      return_add_generic_AC_RND_CONV_false_3_if_7_return_add_generic_AC_RND_CONV_false_3_if_7_nor_nl);
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0 = MUX_v_51_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_1[50:0]),
      stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0w0, inverse_lpi_1_dfm_1);
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50 = MUX_s_1_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_1[50]),
      (stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0w0[50]), inverse_lpi_1_dfm_1);
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_3_exception_sva_1);
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5 = MUX_v_6_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_0[5:0]),
      (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1[9:4]), inverse_lpi_1_dfm_1);
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1 = MUX_v_4_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_1[56:53]),
      (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1[3:0]), inverse_lpi_1_dfm_1);
  assign or_278_nl = or_dcpl_216 | return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
      | operator_11_true_return_26_sva | and_dcpl_166;
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_2_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs, or_278_nl);
  assign return_add_generic_AC_RND_CONV_false_3_e_r_return_add_generic_AC_RND_CONV_false_3_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_6_mux_35 & (~ return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_2_nl))
      | return_add_generic_AC_RND_CONV_false_3_exception_sva_1;
  assign stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0 = MUX_s_1_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_1[52]),
      return_add_generic_AC_RND_CONV_false_3_e_r_return_add_generic_AC_RND_CONV_false_3_e_r_or_1_nl,
      inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_3_r_nan_or_1_nl = operator_11_true_return_26_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_10_unequal_tmp;
  assign and_502_nl = (or_dcpl_216 | and_dcpl_166 | return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
      | or_dcpl_1069) & inverse_lpi_1_dfm_1;
  assign and_510_nl = (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_3_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
      & or_dcpl_431 & (~ return_add_generic_AC_RND_CONV_false_10_op2_nan_sva) & (~(return_add_generic_AC_RND_CONV_false_10_op2_inf_sva
      | return_add_generic_AC_RND_CONV_false_10_op1_inf_sva | operator_11_true_return_26_sva))
      & and_dcpl_385;
  assign return_add_generic_AC_RND_CONV_false_3_r_nan_mux1h_cse = MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_3_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[51]), (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[51]),
      {and_502_nl , and_510_nl , (~ inverse_lpi_1_dfm_1)});
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_not_7_nl = ~ return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
  assign return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(10'b0000000000,
      z_out_9, return_add_generic_AC_RND_CONV_false_e_r_qelse_not_7_nl);
  assign return_add_generic_AC_RND_CONV_false_3_if_5_or_nl = return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_3_mux_10_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_3_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_3_exception_sva_1 = return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | operator_11_true_return_26_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_3_mux_10_nl;
  assign return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_3_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_6_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_24,
      z_out_25, z_out_24[11]);
  assign return_add_generic_AC_RND_CONV_false_6_op2_mu_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_extract_13_return_extract_13_or_1_cse_sva_1,
      return_add_generic_AC_RND_CONV_false_3_r_nan_mux1h_cse, return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_1_return_add_generic_AC_RND_CONV_false_6_op2_normal_return_extract_13_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_50_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_3_r_nan_mux1h_cse,
      stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50, return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_1_return_add_generic_AC_RND_CONV_false_6_op2_normal_return_extract_13_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_49_0_mx0 =
      MUX_v_50_2_2((stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0[50:1]), (stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0[49:0]),
      return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_1_return_add_generic_AC_RND_CONV_false_6_op2_normal_return_extract_13_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1 = (stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0[0])
      & (~ return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_1_return_add_generic_AC_RND_CONV_false_6_op2_normal_return_extract_13_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_6_op2_mu_52_lpi_3_dfm_mx0, and_dcpl_349);
  assign return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_50_mx0
      = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_50_mx0, and_dcpl_349);
  assign return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0
      = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm,
      return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_49_0_mx0, and_dcpl_349);
  assign return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_0_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm,
      return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1, and_dcpl_349);
  assign return_add_generic_AC_RND_CONV_false_6_e1_eq_e2_equal_tmp = ({BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_1
      , reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd , reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1
      , reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2 , reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3})
      == ({stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5 , stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1
      , stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0});
  assign return_add_generic_AC_RND_CONV_false_6_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_16[54]))) | (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_50_mx0
      & (~ (z_out_16[53]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[49])
      & (~ (z_out_16[52]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[48])
      & (~ (z_out_16[51]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[47])
      & (~ (z_out_16[50]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[46])
      & (~ (z_out_16[49]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[45])
      & (~ (z_out_16[48]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[44])
      & (~ (z_out_16[47]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[43])
      & (~ (z_out_16[46]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[42])
      & (~ (z_out_16[45]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[41])
      & (~ (z_out_16[44]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[40])
      & (~ (z_out_16[43]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[39])
      & (~ (z_out_16[42]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[38])
      & (~ (z_out_16[41]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[37])
      & (~ (z_out_16[40]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[36])
      & (~ (z_out_16[39]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[35])
      & (~ (z_out_16[38]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[34])
      & (~ (z_out_16[37]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[33])
      & (~ (z_out_16[36]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[32])
      & (~ (z_out_16[35]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[31])
      & (~ (z_out_16[34]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[30])
      & (~ (z_out_16[33]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[29])
      & (~ (z_out_16[32]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[28])
      & (~ (z_out_16[31]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[27])
      & (~ (z_out_16[30]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[26])
      & (~ (z_out_16[29]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[25])
      & (~ (z_out_16[28]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[24])
      & (~ (z_out_16[27]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[23])
      & (~ (z_out_16[26]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[22])
      & (~ (z_out_16[25]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[21])
      & (~ (z_out_16[24]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[20])
      & (~ (z_out_16[23]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[19])
      & (~ (z_out_16[22]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[18])
      & (~ (z_out_16[21]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[17])
      & (~ (z_out_16[20]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[16])
      & (~ (z_out_16[19]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[15])
      & (~ (z_out_16[18]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[14])
      & (~ (z_out_16[17]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[13])
      & (~ (z_out_16[16]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[12])
      & (~ (z_out_16[15]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[11])
      & (~ (z_out_16[14]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[10])
      & (~ (z_out_16[13]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[9])
      & (~ (z_out_16[12]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[8])
      & (~ (z_out_16[11]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[7])
      & (~ (z_out_16[10]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[6])
      & (~ (z_out_16[9]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[5])
      & (~ (z_out_16[8]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[4])
      & (~ (z_out_16[7]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[3])
      & (~ (z_out_16[6]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[2])
      & (~ (z_out_16[5]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[1])
      & (~ (z_out_16[4]))) | ((return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[0])
      & (~ (z_out_16[3]))) | (return_add_generic_AC_RND_CONV_false_6_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_16[2])));
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_1_if_acc_1_itm_12_1) | (z_out_18[105]);
  assign return_mult_generic_AC_RND_CONV_false_1_e_incr_lpi_3_dfm_2 = ~((~(((z_out_18[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((z_out_18[51]) | return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_or_2))
      | (z_out_18[105]))) | (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_1_zero_m_return_mult_generic_AC_RND_CONV_false_1_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_1_r_zero_return_mult_generic_AC_RND_CONV_false_1_r_zero_nor_mdf_sva_1
      = ~(and_2331_cse | return_mult_generic_AC_RND_CONV_false_1_op2_zero_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_1_r_nan_sva_1 = return_add_generic_AC_RND_CONV_false_6_op2_nan_sva_1
      | (operator_11_true_return_17_sva & (~ return_extract_17_m_zero_sva)) | (return_add_generic_AC_RND_CONV_false_6_op2_inf_sva_1
      & return_mult_generic_AC_RND_CONV_false_1_op2_zero_sva_1) | (and_2331_cse &
      return_mult_generic_AC_RND_CONV_false_1_op2_inf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_1_exp_ovf_return_mult_generic_AC_RND_CONV_false_1_exp_ovf_or_tmp
      = ((return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[10:1]==10'b1111111111)
      & return_mult_generic_AC_RND_CONV_false_exp_ovf_oif_aelse_nor_cse & return_mult_generic_AC_RND_CONV_false_1_e_incr_lpi_3_dfm_2)
      | (z_out_36[11]);
  assign return_mult_generic_AC_RND_CONV_false_1_lor_lpi_3_dfm_1 = return_add_generic_AC_RND_CONV_false_6_op2_inf_sva_1
      | return_mult_generic_AC_RND_CONV_false_1_op2_inf_sva_1 | return_mult_generic_AC_RND_CONV_false_1_exp_ovf_return_mult_generic_AC_RND_CONV_false_1_exp_ovf_or_tmp
      | return_mult_generic_AC_RND_CONV_false_1_r_nan_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_1_return_mult_generic_AC_RND_CONV_false_1_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_tmp_1 | (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_1_and_2_nl = return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_tmp_1
      & (~ (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_1_res_bef_rnd_3_53_1_lpi_3_dfm_1 =
      MUX1HOT_v_53_3_2((z_out_18[104:52]), (z_out_18[103:51]), (z_out_42[53:1]),
      {return_mult_generic_AC_RND_CONV_false_1_return_mult_generic_AC_RND_CONV_false_1_nor_nl
      , return_mult_generic_AC_RND_CONV_false_1_and_2_nl , (z_out_27[12])});
  assign return_mult_generic_AC_RND_CONV_false_1_op2_inf_sva_1 = operator_11_true_return_17_sva
      & return_extract_17_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_1_op2_zero_sva_1 = return_extract_17_return_extract_17_nor_cse_sva
      & return_extract_17_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_mux_1_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_1_if_acc_1_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva, z_out_27[12]);
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_mux_1_nl
      & (~ (z_out_18[105]));
  assign return_extract_13_return_extract_13_or_1_cse_sva_1 = (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5!=6'b000000)
      | (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1!=4'b0000) | stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0;
  assign return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_1_return_add_generic_AC_RND_CONV_false_6_op2_normal_return_extract_13_nor_tmp
      = ~((stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5!=6'b000000) | (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1!=4'b0000)
      | stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0);
  assign return_extract_13_m_zero_return_extract_13_m_zero_nor_tmp = ~(return_add_generic_AC_RND_CONV_false_3_r_nan_mux1h_cse
      | stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50 | (stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0[49:0]!=50'b00000000000000000000000000000000000000000000000000));
  assign return_add_generic_AC_RND_CONV_false_6_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_6_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_6_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_6_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_6_e_dif_sat_or_1_nl);
  assign operator_11_true_13_operator_11_true_13_and_tmp = (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5==6'b111111)
      & (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1==4'b1111) & stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0;
  assign return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_52_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1,
      and_dcpl_260);
  assign return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_51_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0,
      and_dcpl_260);
  assign return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_49_0,
      return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_260);
  assign return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_2_if_acc_1_itm_12_1) | (z_out_18[105]);
  assign return_mult_generic_AC_RND_CONV_false_2_e_incr_lpi_3_dfm_2 = ~((~(((z_out_18[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((z_out_18[51]) | return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_or_2))
      | (z_out_18[105]))) | (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_2_zero_m_return_mult_generic_AC_RND_CONV_false_2_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_2_r_zero_return_mult_generic_AC_RND_CONV_false_2_r_zero_nor_mdf_sva_1
      = ~(return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 | (return_extract_19_return_extract_19_nor_tmp
      & return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp));
  assign return_mult_generic_AC_RND_CONV_false_2_else_2_else_else_mux_nl = MUX_v_11_2_2((return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[10:0]),
      (z_out_36[10:0]), return_mult_generic_AC_RND_CONV_false_2_e_incr_lpi_3_dfm_2);
  assign return_mult_generic_AC_RND_CONV_false_2_else_2_else_return_mult_generic_AC_RND_CONV_false_2_else_2_else_and_nl
      = MUX_v_11_2_2(11'b00000000000, return_mult_generic_AC_RND_CONV_false_2_else_2_else_else_mux_nl,
      return_mult_generic_AC_RND_CONV_false_2_zero_m_return_mult_generic_AC_RND_CONV_false_2_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_2_r_zero_return_mult_generic_AC_RND_CONV_false_2_r_zero_nor_mdf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1 =
      MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_2_else_2_else_return_mult_generic_AC_RND_CONV_false_2_else_2_else_and_nl,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_2_lor_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[0])
      & operator_11_true_return_15_sva;
  assign return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1 = return_mult_generic_AC_RND_CONV_false_2_m_r_51_lpi_3_dfm_mx1
      | return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0 = MUX_s_1_2_2((return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1[50]),
      return_mult_generic_AC_RND_CONV_false_2_m_r_51_lpi_3_dfm_mx1, return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_1_tmp);
  assign return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0 = MUX_v_50_2_2((return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1[49:0]),
      (return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1[50:1]), return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_1_tmp);
  assign return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1 = (return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1[0])
      & return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_1_tmp;
  assign and_514_nl = return_mult_generic_AC_RND_CONV_false_2_zero_m_return_mult_generic_AC_RND_CONV_false_2_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_2_r_zero_return_mult_generic_AC_RND_CONV_false_2_r_zero_nor_mdf_sva_1
      & (~(operator_11_true_19_operator_11_true_19_and_tmp | return_mult_generic_AC_RND_CONV_false_2_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_2_exp_ovf_oif_aelse_and_tmp
      | (z_out_36[11])));
  assign return_mult_generic_AC_RND_CONV_false_2_m_r_51_lpi_3_dfm_mx1 = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_2_r_nan_sva_1,
      (z_out_6[51]), and_514_nl);
  assign return_mult_generic_AC_RND_CONV_false_2_oelse_3_return_mult_generic_AC_RND_CONV_false_2_if_3_nor_nl
      = ~((~ return_mult_generic_AC_RND_CONV_false_2_zero_m_return_mult_generic_AC_RND_CONV_false_2_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_2_r_zero_return_mult_generic_AC_RND_CONV_false_2_r_zero_nor_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_2_lor_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (z_out_6[50:0]), return_mult_generic_AC_RND_CONV_false_2_oelse_3_return_mult_generic_AC_RND_CONV_false_2_if_3_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_7_e1_eq_e2_equal_tmp = ({BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1
      , BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2}) == (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1);
  assign return_add_generic_AC_RND_CONV_false_8_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_26,
      z_out_23, z_out_26[11]);
  assign return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[0])
      & return_add_generic_AC_RND_CONV_false_10_do_sub_sva;
  assign return_add_generic_AC_RND_CONV_false_8_e1_eq_e2_equal_tmp = ({BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1
      , reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd , reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1})
      == (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1);
  assign return_add_generic_AC_RND_CONV_false_7_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_52_lpi_3_dfm_mx0
      & (~ (z_out_16[54]))) | (return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_51_lpi_3_dfm_mx0
      & (~ (z_out_16[53]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_16[52]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_16[51]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_16[50]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_16[49]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_16[48]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_16[47]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_16[46]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_16[45]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_16[44]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_16[43]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_16[42]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_16[41]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_16[40]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_16[39]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_16[38]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_16[37]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_16[36]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_16[35]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_16[34]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_16[33]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_16[32]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_16[31]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_16[30]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_16[29]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_16[28]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_16[27]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_16[26]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_16[25]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_16[24]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_16[23]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_16[22]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_16[21]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_16[20]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_16[19]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_16[18]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_16[17]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_16[16]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_16[15]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_16[14]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_16[13]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_16[12]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_16[11]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_16[10]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_16[9]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_16[8]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_16[7]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_16[6]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_16[5]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_16[4]))) | ((return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_16[3]))) | (return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm_mx1
      & (~ (z_out_16[2])));
  assign return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_1_tmp
      = (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1!=11'b00000000000);
  assign return_mult_generic_AC_RND_CONV_false_2_r_nan_sva_1 = (operator_11_true_19_operator_11_true_19_and_tmp
      & (~ return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp)) | (return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1
      & return_mult_generic_AC_RND_CONV_false_2_op2_inf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_2_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_2_exp_ovf_oif_aelse_and_tmp
      = (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[10:1]==10'b1111111111)
      & return_mult_generic_AC_RND_CONV_false_exp_ovf_oif_aelse_nor_cse & return_mult_generic_AC_RND_CONV_false_2_e_incr_lpi_3_dfm_2;
  assign return_mult_generic_AC_RND_CONV_false_2_lor_lpi_3_dfm_1 = return_mult_generic_AC_RND_CONV_false_2_op2_inf_sva_1
      | return_mult_generic_AC_RND_CONV_false_2_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_2_exp_ovf_oif_aelse_and_tmp
      | (z_out_36[11]) | return_mult_generic_AC_RND_CONV_false_2_r_nan_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_2_return_mult_generic_AC_RND_CONV_false_2_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_2_if_1_and_1_tmp_1 | (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_2_and_2_nl = return_mult_generic_AC_RND_CONV_false_2_if_1_and_1_tmp_1
      & (~ (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_2_res_bef_rnd_3_53_1_lpi_3_dfm_1 =
      MUX1HOT_v_53_3_2((z_out_18[104:52]), (z_out_18[103:51]), (z_out_42[53:1]),
      {return_mult_generic_AC_RND_CONV_false_2_return_mult_generic_AC_RND_CONV_false_2_nor_nl
      , return_mult_generic_AC_RND_CONV_false_2_and_2_nl , (z_out_27[12])});
  assign return_mult_generic_AC_RND_CONV_false_2_op2_inf_sva_1 = operator_11_true_19_operator_11_true_19_and_tmp
      & return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp;
  assign return_extract_19_return_extract_19_nor_tmp = ~((return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1);
  assign return_extract_19_m_zero_return_extract_19_m_zero_nor_tmp = ~(return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_mux_1_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_2_if_acc_1_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva, z_out_27[12]);
  assign return_mult_generic_AC_RND_CONV_false_2_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_mux_1_nl
      & (~ (z_out_18[105]));
  assign return_extract_19_return_extract_19_or_sva_1 = (return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_6_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | (return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva & return_add_generic_AC_RND_CONV_false_11_do_sub_sva);
  assign and_521_nl = (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
      & or_dcpl_431 & and_dcpl_399 & (~(return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva));
  assign return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[51]), and_521_nl);
  assign return_add_generic_AC_RND_CONV_false_6_if_7_return_add_generic_AC_RND_CONV_false_6_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_6_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[50:0]),
      return_add_generic_AC_RND_CONV_false_6_if_7_return_add_generic_AC_RND_CONV_false_6_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_6_exception_sva_1);
  assign or_290_nl = or_dcpl_228 | or_dcpl_225 | and_dcpl_166;
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_5_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs, or_290_nl);
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_6_mux_35
      & (~ return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_5_nl)) | return_add_generic_AC_RND_CONV_false_6_exception_sva_1;
  assign operator_11_true_19_operator_11_true_19_and_tmp = (return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_6_if_5_or_nl = return_add_generic_AC_RND_CONV_false_6_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_6_mux_16_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_6_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_6_exception_sva_1 = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_6_mux_16_nl;
  assign return_add_generic_AC_RND_CONV_false_6_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_51_lpi_3_dfm_mx3 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm, return_add_generic_AC_RND_CONV_false_20_op2_mu_1_51_lpi_3_dfm_mx0,
      and_dcpl_264);
  assign return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_52_lpi_3_dfm_mx3 =
      MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm, return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1,
      and_dcpl_264);
  assign return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_9_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_9_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_9_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_9_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[49:0]),
      return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_261);
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_149_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[49])
      & (~ (z_out_16[52]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_141_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[48])
      & (~ (z_out_16[51]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_133_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[47])
      & (~ (z_out_16[50]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_125_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[46])
      & (~ (z_out_16[49]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_117_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[45])
      & (~ (z_out_16[48]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_109_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[44])
      & (~ (z_out_16[47]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_101_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[43])
      & (~ (z_out_16[46]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_93_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[42])
      & (~ (z_out_16[45]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_85_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[41])
      & (~ (z_out_16[44]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_77_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[40])
      & (~ (z_out_16[43]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_69_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[39])
      & (~ (z_out_16[42]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_61_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[38])
      & (~ (z_out_16[41]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_155_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[37])
      & (~ (z_out_16[40]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_147_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[36])
      & (~ (z_out_16[39]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_139_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[35])
      & (~ (z_out_16[38]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_131_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[34])
      & (~ (z_out_16[37]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_123_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[33])
      & (~ (z_out_16[36]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_115_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[32])
      & (~ (z_out_16[35]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_107_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[31])
      & (~ (z_out_16[34]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_99_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[30])
      & (~ (z_out_16[33]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_91_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[29])
      & (~ (z_out_16[32]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_83_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[28])
      & (~ (z_out_16[31]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_75_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[27])
      & (~ (z_out_16[30]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_67_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[26])
      & (~ (z_out_16[29]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_59_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[25])
      & (~ (z_out_16[28]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_153_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[24])
      & (~ (z_out_16[27]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_145_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[23])
      & (~ (z_out_16[26]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_137_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[22])
      & (~ (z_out_16[25]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_129_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[21])
      & (~ (z_out_16[24]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_121_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[20])
      & (~ (z_out_16[23]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_113_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[19])
      & (~ (z_out_16[22]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_105_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[18])
      & (~ (z_out_16[21]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_97_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[17])
      & (~ (z_out_16[20]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_89_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[16])
      & (~ (z_out_16[19]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_81_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[15])
      & (~ (z_out_16[18]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_73_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[14])
      & (~ (z_out_16[17]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_65_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[13])
      & (~ (z_out_16[16]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_57_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[12])
      & (~ (z_out_16[15]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_151_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[11])
      & (~ (z_out_16[14]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_143_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[10])
      & (~ (z_out_16[13]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_135_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[9])
      & (~ (z_out_16[12]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_127_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[8])
      & (~ (z_out_16[11]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_119_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[7])
      & (~ (z_out_16[10]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_111_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[6])
      & (~ (z_out_16[9]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_103_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[5])
      & (~ (z_out_16[8]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_95_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[4])
      & (~ (z_out_16[7]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_87_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[3])
      & (~ (z_out_16[6]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_79_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[2])
      & (~ (z_out_16[5]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_71_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[1])
      & (~ (z_out_16[4]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_63_cse = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[0])
      & (~ (z_out_16[3]));
  assign return_add_generic_AC_RND_CONV_false_8_res_mant_3_0_sva_1 = return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_54
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_56 | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_149_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_141_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_133_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_125_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_117_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_109_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_101_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_93_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_85_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_77_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_69_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_61_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_155_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_147_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_139_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_131_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_123_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_115_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_107_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_99_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_91_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_83_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_75_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_67_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_59_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_153_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_145_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_137_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_129_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_121_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_113_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_105_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_97_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_89_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_81_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_73_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_65_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_57_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_151_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_143_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_135_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_127_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_119_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_111_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_103_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_95_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_87_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_79_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_71_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_63_cse | return_add_generic_AC_RND_CONV_false_5_sticky_bit_and_54;
  assign return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_7_exception_sva_1);
  assign or_299_nl = or_dcpl_237 | or_dcpl_235;
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_7_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs, or_299_nl);
  assign return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_6_mux_35
      & (~ return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_7_nl)) | return_add_generic_AC_RND_CONV_false_7_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_7_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_9_op2_nan_sva_mx7w0
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_9_op2_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_16_do_sub_sva);
  assign and_529_nl = (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_7_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
      & or_dcpl_431 & and_dcpl_408;
  assign return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[51]), and_529_nl);
  assign return_add_generic_AC_RND_CONV_false_7_if_7_return_add_generic_AC_RND_CONV_false_7_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_7_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[50:0]),
      return_add_generic_AC_RND_CONV_false_7_if_7_return_add_generic_AC_RND_CONV_false_7_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_9_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_23,
      z_out_25, z_out_23[11]);
  assign return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1 = (stage_PE_1_x_re_d_sva[0])
      & return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva;
  assign return_extract_25_return_extract_25_or_2_nl = (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_extract_25_return_extract_25_or_2_nl,
      return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1[50]), return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0 = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1[50:1]),
      (return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1[49:0]), return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1[0])
      & (~ return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_9_e1_eq_e2_equal_tmp = (stage_PE_1_x_re_d_sva[62:52])
      == ({return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1});
  assign return_add_generic_AC_RND_CONV_false_11_e_dif_qr_lpi_3_dfm_mx0_10_0 = MUX_v_11_2_2((z_out_23[10:0]),
      (z_out_25[10:0]), z_out_23[11]);
  assign return_add_generic_AC_RND_CONV_false_9_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_22_op1_mu_mux_cse
      & (~ (z_out_17[54]))) | (return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_cse
      & (~ (z_out_17[53]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_17[52]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_17[51]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_17[50]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_17[49]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_17[48]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_17[47]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_17[46]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_17[45]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_17[44]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_17[43]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_17[42]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_17[41]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_17[40]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_17[39]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_17[38]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_17[37]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_17[36]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_17[35]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_17[34]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_17[33]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_17[32]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_17[31]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_17[30]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_17[29]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_17[28]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_17[27]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_17[26]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_17[25]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_17[24]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_17[23]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_17[22]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_17[21]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_17[20]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_17[19]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_17[18]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_17[17]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_17[16]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_17[15]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_17[14]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_17[13]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_17[12]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_17[11]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_17[10]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_17[9]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_17[8]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_17[7]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_17[6]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_17[5]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_17[4]))) | ((return_add_generic_AC_RND_CONV_false_9_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_17[3]))) | (return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_2_cse
      & (~ (z_out_17[2])));
  assign return_add_generic_AC_RND_CONV_false_9_return_add_generic_AC_RND_CONV_false_9_if_1_return_add_generic_AC_RND_CONV_false_9_op2_normal_return_extract_25_nor_tmp
      = ~((return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_7_if_5_or_nl = return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_7_mux_18_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_7_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_7_exception_sva_1 = return_add_generic_AC_RND_CONV_false_9_op2_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_9_op2_nan_sva_mx7w0
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_7_mux_18_nl;
  assign return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_7_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_2_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[49])
      & (~ (z_out_16[52]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_3_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[48])
      & (~ (z_out_16[51]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_4_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[47])
      & (~ (z_out_16[50]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_5_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[46])
      & (~ (z_out_16[49]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_6_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[45])
      & (~ (z_out_16[48]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_7_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[44])
      & (~ (z_out_16[47]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_8_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[43])
      & (~ (z_out_16[46]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_9_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[42])
      & (~ (z_out_16[45]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_10_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[41])
      & (~ (z_out_16[44]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_11_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[40])
      & (~ (z_out_16[43]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_12_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[39])
      & (~ (z_out_16[42]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_13_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[38])
      & (~ (z_out_16[41]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_14_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[37])
      & (~ (z_out_16[40]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_15_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[36])
      & (~ (z_out_16[39]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_16_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[35])
      & (~ (z_out_16[38]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_17_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[34])
      & (~ (z_out_16[37]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_18_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[33])
      & (~ (z_out_16[36]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_19_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[32])
      & (~ (z_out_16[35]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_20_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[31])
      & (~ (z_out_16[34]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_21_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[30])
      & (~ (z_out_16[33]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_22_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[29])
      & (~ (z_out_16[32]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_23_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[28])
      & (~ (z_out_16[31]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_24_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[27])
      & (~ (z_out_16[30]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_25_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[26])
      & (~ (z_out_16[29]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_26_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[25])
      & (~ (z_out_16[28]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_27_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[24])
      & (~ (z_out_16[27]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_28_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[23])
      & (~ (z_out_16[26]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_29_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[22])
      & (~ (z_out_16[25]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_30_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[21])
      & (~ (z_out_16[24]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_31_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[20])
      & (~ (z_out_16[23]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_32_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[19])
      & (~ (z_out_16[22]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_33_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[18])
      & (~ (z_out_16[21]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_34_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[17])
      & (~ (z_out_16[20]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_35_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[16])
      & (~ (z_out_16[19]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_36_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[15])
      & (~ (z_out_16[18]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_37_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[14])
      & (~ (z_out_16[17]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_38_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[13])
      & (~ (z_out_16[16]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_39_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[12])
      & (~ (z_out_16[15]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_40_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[11])
      & (~ (z_out_16[14]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_41_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[10])
      & (~ (z_out_16[13]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_42_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[9])
      & (~ (z_out_16[12]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_43_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[8])
      & (~ (z_out_16[11]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_44_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[7])
      & (~ (z_out_16[10]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_45_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[6])
      & (~ (z_out_16[9]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_46_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[5])
      & (~ (z_out_16[8]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_47_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[4])
      & (~ (z_out_16[7]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_48_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[3])
      & (~ (z_out_16[6]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_49_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[2])
      & (~ (z_out_16[5]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_50_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[1])
      & (~ (z_out_16[4]));
  assign return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_51_cse = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[0])
      & (~ (z_out_16[3]));
  assign return_add_generic_AC_RND_CONV_false_11_res_mant_3_0_sva_1 = return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_54
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_56 | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_2_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_3_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_4_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_5_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_6_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_7_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_8_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_9_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_10_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_11_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_12_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_13_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_14_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_15_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_16_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_17_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_18_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_19_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_20_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_21_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_22_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_23_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_24_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_25_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_26_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_27_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_28_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_29_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_30_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_31_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_32_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_33_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_34_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_35_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_36_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_37_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_38_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_39_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_40_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_41_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_42_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_43_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_44_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_45_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_46_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_47_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_48_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_49_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_50_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_51_cse | return_add_generic_AC_RND_CONV_false_5_sticky_bit_and_54;
  assign return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_8_exception_sva_1);
  assign or_308_nl = return_add_generic_AC_RND_CONV_false_8_r_inf_lpi_3_dfm_2 | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva
      | or_dcpl_244;
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_9_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs, or_308_nl);
  assign return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_6_mux_35
      & (~ return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_9_nl)) | return_add_generic_AC_RND_CONV_false_8_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_8_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_8_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | (return_add_generic_AC_RND_CONV_false_8_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva & return_add_generic_AC_RND_CONV_false_14_op2_inf_sva);
  assign and_534_nl = (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_8_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
      & or_dcpl_431 & and_dcpl_413;
  assign return_add_generic_AC_RND_CONV_false_8_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[51]), and_534_nl);
  assign return_add_generic_AC_RND_CONV_false_8_if_7_return_add_generic_AC_RND_CONV_false_8_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_8_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[50:0]),
      return_add_generic_AC_RND_CONV_false_8_if_7_return_add_generic_AC_RND_CONV_false_8_if_7_nor_nl);
  assign return_extract_27_return_extract_27_or_2_nl = (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_extract_27_return_extract_27_or_2_nl,
      return_add_generic_AC_RND_CONV_false_8_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_10_op2_mu_1_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_m_r_51_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1[50]), return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_10_op2_mu_1_50_1_lpi_3_dfm_mx0 = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1[50:1]),
      (return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1[49:0]), return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1[0])
      & (~ return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49:0]),
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_326);
  assign return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_equal_tmp = (stage_PE_1_x_im_d_sva[62:52])
      == ({return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1});
  assign return_add_generic_AC_RND_CONV_false_10_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_10_exp_mux_5_cse
      & (~ (z_out_16[54]))) | (return_add_generic_AC_RND_CONV_false_5_op_smaller_mux_1_cse
      & (~ (z_out_16[53]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_16[52]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_16[51]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_16[50]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_16[49]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_16[48]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_16[47]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_16[46]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_16[45]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_16[44]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_16[43]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_16[42]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_16[41]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_16[40]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_16[39]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_16[38]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_16[37]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_16[36]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_16[35]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_16[34]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_16[33]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_16[32]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_16[31]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_16[30]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_16[29]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_16[28]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_16[27]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_16[26]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_16[25]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_16[24]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_16[23]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_16[22]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_16[21]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_16[20]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_16[19]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_16[18]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_16[17]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_16[16]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_16[15]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_16[14]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_16[13]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_16[12]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_16[11]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_16[10]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_16[9]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_16[8]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_16[7]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_16[6]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_16[5]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_16[4]))) | ((return_add_generic_AC_RND_CONV_false_10_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_16[3]))) | (return_add_generic_AC_RND_CONV_false_1_op_bigger_mux_4_cse
      & (~ (z_out_16[2])));
  assign return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_if_1_return_add_generic_AC_RND_CONV_false_10_op2_normal_return_extract_27_nor_tmp
      = ~((return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_8_op1_nan_sva_1 = operator_11_true_return_17_sva
      & (~ return_extract_1_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_8_op1_inf_sva_1 = operator_11_true_return_17_sva
      & return_extract_1_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_8_if_5_or_nl = return_add_generic_AC_RND_CONV_false_8_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_8_mux_14_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_8_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_8_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_8_exception_sva_1 = return_add_generic_AC_RND_CONV_false_8_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_8_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_8_mux_14_nl;
  assign return_add_generic_AC_RND_CONV_false_8_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_8_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_12_res_mant_3_0_sva_1 = return_add_generic_AC_RND_CONV_false_12_sticky_bit_and_54
      | return_add_generic_AC_RND_CONV_false_12_sticky_bit_and_56 | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_149_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_141_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_133_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_125_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_117_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_109_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_101_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_93_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_85_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_77_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_69_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_61_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_155_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_147_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_139_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_131_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_123_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_115_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_107_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_99_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_91_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_83_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_75_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_67_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_59_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_153_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_145_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_137_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_129_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_121_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_113_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_105_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_97_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_89_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_81_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_73_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_65_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_57_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_151_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_143_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_135_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_127_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_119_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_111_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_103_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_95_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_87_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_79_cse | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_71_cse
      | return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_63_cse | return_add_generic_AC_RND_CONV_false_12_sticky_bit_and_58;
  assign return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp
      = (return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_5_cse[9:0]==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_or_2_cse
      & (return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_5_cse[11:10]==2'b00);
  assign return_add_generic_AC_RND_CONV_false_9_if_5_or_nl = return_add_generic_AC_RND_CONV_false_9_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_9_mux_17_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_9_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_9_exception_sva_1 = return_add_generic_AC_RND_CONV_false_23_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_9_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_23_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_9_op2_nan_sva_mx7w0 | return_add_generic_AC_RND_CONV_false_9_mux_17_nl;
  assign return_add_generic_AC_RND_CONV_false_9_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_9_exception_sva_1
      | operator_11_true_return_24_sva;
  assign return_add_generic_AC_RND_CONV_false_9_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_9_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_10_if_5_or_nl = return_add_generic_AC_RND_CONV_false_10_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_10_mux_17_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_10_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_10_exception_sva_1 = return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_10_mux_17_nl;
  assign return_add_generic_AC_RND_CONV_false_10_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_10_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_10_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_10_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_11_if_5_or_nl = return_add_generic_AC_RND_CONV_false_11_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_11_mux_10_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_11_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_11_exception_sva_1 = return_add_generic_AC_RND_CONV_false_23_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_inf_sva | return_add_generic_AC_RND_CONV_false_23_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva | return_add_generic_AC_RND_CONV_false_11_mux_10_nl;
  assign return_add_generic_AC_RND_CONV_false_11_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_11_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_11_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_12_if_5_or_nl = return_add_generic_AC_RND_CONV_false_12_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_12_mux_10_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_12_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_12_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_12_exception_sva_1 = return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_12_mux_10_nl;
  assign return_add_generic_AC_RND_CONV_false_12_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_12_exception_sva_1
      | operator_11_true_return_24_sva;
  assign return_add_generic_AC_RND_CONV_false_12_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_12_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign nl_return_add_generic_AC_RND_CONV_false_4_e_dif_acc_tmp = ({1'b1 , (~ (O_1_out_1[61:52]))})
      + conv_u2s_10_11(O_1_out[61:52]) + 11'b00000000001;
  assign return_add_generic_AC_RND_CONV_false_4_e_dif_acc_tmp = nl_return_add_generic_AC_RND_CONV_false_4_e_dif_acc_tmp[10:0];
  assign return_add_generic_AC_RND_CONV_false_4_e1_eq_e2_equal_tmp = (O_1_out[61:52])
      == (O_1_out_1[61:52]);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_12_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[50]),
      (stage_PE_1_gm_im_d_mux_2_cse[50]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_13_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[49]),
      (stage_PE_1_gm_im_d_mux_2_cse[49]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_14_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[48]),
      (stage_PE_1_gm_im_d_mux_2_cse[48]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_15_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[47]),
      (stage_PE_1_gm_im_d_mux_2_cse[47]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_16_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[46]),
      (stage_PE_1_gm_im_d_mux_2_cse[46]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_17_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[45]),
      (stage_PE_1_gm_im_d_mux_2_cse[45]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_18_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[44]),
      (stage_PE_1_gm_im_d_mux_2_cse[44]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_19_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[43]),
      (stage_PE_1_gm_im_d_mux_2_cse[43]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_20_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[42]),
      (stage_PE_1_gm_im_d_mux_2_cse[42]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_21_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[41]),
      (stage_PE_1_gm_im_d_mux_2_cse[41]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_22_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[40]),
      (stage_PE_1_gm_im_d_mux_2_cse[40]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_23_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[39]),
      (stage_PE_1_gm_im_d_mux_2_cse[39]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_24_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[38]),
      (stage_PE_1_gm_im_d_mux_2_cse[38]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_25_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[37]),
      (stage_PE_1_gm_im_d_mux_2_cse[37]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_26_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[36]),
      (stage_PE_1_gm_im_d_mux_2_cse[36]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_27_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[35]),
      (stage_PE_1_gm_im_d_mux_2_cse[35]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_28_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[34]),
      (stage_PE_1_gm_im_d_mux_2_cse[34]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_29_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[33]),
      (stage_PE_1_gm_im_d_mux_2_cse[33]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_30_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[32]),
      (stage_PE_1_gm_im_d_mux_2_cse[32]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_31_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[31]),
      (stage_PE_1_gm_im_d_mux_2_cse[31]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_32_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[30]),
      (stage_PE_1_gm_im_d_mux_2_cse[30]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_33_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[29]),
      (stage_PE_1_gm_im_d_mux_2_cse[29]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_34_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[28]),
      (stage_PE_1_gm_im_d_mux_2_cse[28]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_35_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[27]),
      (stage_PE_1_gm_im_d_mux_2_cse[27]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_36_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[26]),
      (stage_PE_1_gm_im_d_mux_2_cse[26]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_37_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[25]),
      (stage_PE_1_gm_im_d_mux_2_cse[25]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_38_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[24]),
      (stage_PE_1_gm_im_d_mux_2_cse[24]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_39_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[23]),
      (stage_PE_1_gm_im_d_mux_2_cse[23]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_40_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[22]),
      (stage_PE_1_gm_im_d_mux_2_cse[22]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_41_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[21]),
      (stage_PE_1_gm_im_d_mux_2_cse[21]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_42_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[20]),
      (stage_PE_1_gm_im_d_mux_2_cse[20]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_43_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[19]),
      (stage_PE_1_gm_im_d_mux_2_cse[19]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_44_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[18]),
      (stage_PE_1_gm_im_d_mux_2_cse[18]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_45_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[17]),
      (stage_PE_1_gm_im_d_mux_2_cse[17]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_46_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[16]),
      (stage_PE_1_gm_im_d_mux_2_cse[16]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_47_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[15]),
      (stage_PE_1_gm_im_d_mux_2_cse[15]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_48_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[14]),
      (stage_PE_1_gm_im_d_mux_2_cse[14]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_49_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[13]),
      (stage_PE_1_gm_im_d_mux_2_cse[13]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_50_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[12]),
      (stage_PE_1_gm_im_d_mux_2_cse[12]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_51_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[11]),
      (stage_PE_1_gm_im_d_mux_2_cse[11]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_52_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[10]),
      (stage_PE_1_gm_im_d_mux_2_cse[10]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_53_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[9]),
      (stage_PE_1_gm_im_d_mux_2_cse[9]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_54_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[8]),
      (stage_PE_1_gm_im_d_mux_2_cse[8]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_55_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[7]),
      (stage_PE_1_gm_im_d_mux_2_cse[7]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_56_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[6]),
      (stage_PE_1_gm_im_d_mux_2_cse[6]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_57_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[5]),
      (stage_PE_1_gm_im_d_mux_2_cse[5]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_58_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[4]),
      (stage_PE_1_gm_im_d_mux_2_cse[4]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_59_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[3]),
      (stage_PE_1_gm_im_d_mux_2_cse[3]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_60_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[2]),
      (stage_PE_1_gm_im_d_mux_2_cse[2]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_61_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[1]),
      (stage_PE_1_gm_im_d_mux_2_cse[1]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_62_nl = MUX_s_1_2_2((stage_PE_1_gm_re_d_mux_cse[0]),
      (stage_PE_1_gm_im_d_mux_2_cse[0]), and_dcpl_257);
  assign return_add_generic_AC_RND_CONV_false_17_res_mant_3_0_sva_1 = return_add_generic_AC_RND_CONV_false_4_sticky_bit_and_cse
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_12_nl & (~ (z_out_16[53])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_13_nl & (~ (z_out_16[52])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_14_nl & (~ (z_out_16[51])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_15_nl & (~ (z_out_16[50])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_16_nl & (~ (z_out_16[49])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_17_nl & (~ (z_out_16[48])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_18_nl & (~ (z_out_16[47])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_19_nl & (~ (z_out_16[46])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_20_nl & (~ (z_out_16[45])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_21_nl & (~ (z_out_16[44])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_22_nl & (~ (z_out_16[43])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_23_nl & (~ (z_out_16[42])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_24_nl & (~ (z_out_16[41])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_25_nl & (~ (z_out_16[40])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_26_nl & (~ (z_out_16[39])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_27_nl & (~ (z_out_16[38])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_28_nl & (~ (z_out_16[37])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_29_nl & (~ (z_out_16[36])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_30_nl & (~ (z_out_16[35])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_31_nl & (~ (z_out_16[34])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_32_nl & (~ (z_out_16[33])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_33_nl & (~ (z_out_16[32])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_34_nl & (~ (z_out_16[31])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_35_nl & (~ (z_out_16[30])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_36_nl & (~ (z_out_16[29])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_37_nl & (~ (z_out_16[28])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_38_nl & (~ (z_out_16[27])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_39_nl & (~ (z_out_16[26])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_40_nl & (~ (z_out_16[25])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_41_nl & (~ (z_out_16[24])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_42_nl & (~ (z_out_16[23])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_43_nl & (~ (z_out_16[22])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_44_nl & (~ (z_out_16[21])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_45_nl & (~ (z_out_16[20])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_46_nl & (~ (z_out_16[19])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_47_nl & (~ (z_out_16[18])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_48_nl & (~ (z_out_16[17])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_49_nl & (~ (z_out_16[16])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_50_nl & (~ (z_out_16[15])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_51_nl & (~ (z_out_16[14])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_52_nl & (~ (z_out_16[13])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_53_nl & (~ (z_out_16[12])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_54_nl & (~ (z_out_16[11])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_55_nl & (~ (z_out_16[10])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_56_nl & (~ (z_out_16[9])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_57_nl & (~ (z_out_16[8])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_58_nl & (~ (z_out_16[7])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_59_nl & (~ (z_out_16[6])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_60_nl & (~ (z_out_16[5])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_61_nl & (~ (z_out_16[4])))
      | (return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_62_nl & (~ (z_out_16[3])))
      | return_add_generic_AC_RND_CONV_false_4_sticky_bit_and_52_cse;
  assign nl_return_add_generic_AC_RND_CONV_false_17_acc_2_nl =  -(z_out_37[10:0]);
  assign return_add_generic_AC_RND_CONV_false_17_acc_2_nl = nl_return_add_generic_AC_RND_CONV_false_17_acc_2_nl[10:0];
  assign return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10_1 = readslicef_11_1_10(return_add_generic_AC_RND_CONV_false_17_acc_2_nl);
  assign return_add_generic_AC_RND_CONV_false_17_if_5_or_1_nl = return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10_1
      | return_add_generic_AC_RND_CONV_false_4_if_5_return_add_generic_AC_RND_CONV_false_4_if_5_nor_cse;
  assign return_add_generic_AC_RND_CONV_false_17_mux_15_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10_1,
      return_add_generic_AC_RND_CONV_false_17_if_5_or_1_nl, z_out_6[53]);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_qelse_or_svs_1 = all_same_out
      | (~ return_add_generic_AC_RND_CONV_false_17_mux_15_nl);
  assign return_add_generic_AC_RND_CONV_false_17_mux_10_itm = MUX_v_6_2_2((drf_qr_lval_4_smx_9_0_lpi_3_dfm_mx0[5:0]),
      rtn_out, return_add_generic_AC_RND_CONV_false_17_acc_2_itm_10_1);
  assign return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_or_tmp
      = (O_1_out[61:52]!=10'b0000000000);
  assign drf_qr_lval_16_smx_lpi_3_dfm_mx0_10_5 = MUX_v_6_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_0[5:0]),
      (in_f_d_rsci_q_d[62:57]), and_dcpl_262);
  assign drf_qr_lval_16_smx_lpi_3_dfm_mx0_4_0 = MUX_v_5_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_1[56:52]),
      (in_f_d_rsci_q_d[56:52]), and_dcpl_262);
  assign return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1 = (in_f_d_rsci_q_d[0])
      & return_add_generic_AC_RND_CONV_false_13_return_add_generic_AC_RND_CONV_false_13_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0
      = MUX_v_51_2_2(return_extract_32_mux_4_cse, return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm,
      and_dcpl_262);
  assign return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp = (in_f_d_rsci_q_d[62:52])
      == ({(stage_PE_1_tmp_im_d_1_sva_1_rsp_0[5:0]) , (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[56:52])});
  assign return_add_generic_AC_RND_CONV_false_13_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx6
      & (~ (z_out_16[54]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_16[53]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_16[52]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_16[51]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_16[50]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_16[49]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_16[48]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_16[47]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_16[46]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_16[45]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_16[44]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_16[43]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_16[42]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_16[41]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_16[40]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_16[39]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_16[38]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_16[37]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_16[36]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_16[35]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_16[34]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_16[33]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_16[32]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_16[31]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_16[30]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_16[29]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_16[28]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_16[27]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_16[26]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_16[25]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_16[24]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_16[23]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_16[22]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_16[21]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_16[20]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_16[19]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_16[18]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_16[17]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_16[16]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_16[15]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_16[14]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_16[13]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_16[12]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_16[11]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_16[10]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_16[9]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_16[8]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_16[7]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_16[6]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_16[5]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_16[4]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_16[3]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx5
      & (~ (z_out_16[2])));
  assign return_add_generic_AC_RND_CONV_false_15_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx6
      & (~ (z_out_17[54]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_17[53]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_17[52]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_17[51]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_17[50]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_17[49]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_17[48]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_17[47]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_17[46]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_17[45]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_17[44]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_17[43]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_17[42]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_17[41]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_17[40]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_17[39]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_17[38]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_17[37]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_17[36]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_17[35]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_17[34]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_17[33]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_17[32]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_17[31]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_17[30]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_17[29]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_17[28]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_17[27]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_17[26]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_17[25]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_17[24]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_17[23]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_17[22]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_17[21]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_17[20]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_17[19]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_17[18]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_17[17]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_17[16]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_17[15]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_17[14]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_17[13]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_17[12]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_17[11]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_17[10]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_17[9]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_17[8]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_17[7]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_17[6]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_17[5]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_17[4]))) | ((return_add_generic_AC_RND_CONV_false_13_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_17[3]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx5
      & (~ (z_out_17[2])));
  assign return_add_generic_AC_RND_CONV_false_13_mux_28_itm_4_0 = MUX_v_5_2_2(drf_qr_lval_16_smx_lpi_3_dfm_mx0_4_0,
      (rtn_out[4:0]), return_add_generic_AC_RND_CONV_false_13_acc_2_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_13_if_5_or_nl = return_add_generic_AC_RND_CONV_false_13_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_13_mux_16_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_13_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_13_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_13_exception_sva_1 = return_add_generic_AC_RND_CONV_false_9_op2_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_9_op2_nan_sva_mx7w0
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_13_mux_16_nl;
  assign return_add_generic_AC_RND_CONV_false_13_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_13_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_13_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_13_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0
      = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm,
      return_extract_32_mux_4_cse, and_dcpl_263);
  assign return_add_generic_AC_RND_CONV_false_14_e1_eq_e2_equal_tmp = (stage_PE_1_x_im_d_sva[62:52])
      == (in_f_d_rsci_q_d[62:52]);
  assign return_add_generic_AC_RND_CONV_false_14_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx7
      & (~ (z_out_16[54]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_16[53]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_16[52]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_16[51]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_16[50]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_16[49]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_16[48]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_16[47]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_16[46]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_16[45]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_16[44]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_16[43]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_16[42]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_16[41]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_16[40]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_16[39]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_16[38]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_16[37]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_16[36]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_16[35]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_16[34]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_16[33]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_16[32]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_16[31]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_16[30]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_16[29]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_16[28]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_16[27]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_16[26]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_16[25]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_16[24]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_16[23]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_16[22]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_16[21]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_16[20]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_16[19]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_16[18]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_16[17]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_16[16]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_16[15]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_16[14]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_16[13]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_16[12]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_16[11]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_16[10]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_16[9]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_16[8]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_16[7]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_16[6]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_16[5]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_16[4]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_16[3]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx6
      & (~ (z_out_16[2])));
  assign return_add_generic_AC_RND_CONV_false_16_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm_mx7
      & (~ (z_out_17[54]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[50])
      & (~ (z_out_17[53]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_17[52]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_17[51]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_17[50]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_17[49]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_17[48]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_17[47]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_17[46]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_17[45]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_17[44]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_17[43]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_17[42]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_17[41]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_17[40]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_17[39]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_17[38]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_17[37]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_17[36]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_17[35]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_17[34]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_17[33]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_17[32]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_17[31]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_17[30]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_17[29]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_17[28]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_17[27]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_17[26]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_17[25]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_17[24]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_17[23]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_17[22]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_17[21]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_17[20]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_17[19]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_17[18]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_17[17]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_17[16]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_17[15]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_17[14]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_17[13]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_17[12]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_17[11]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_17[10]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_17[9]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_17[8]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_17[7]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_17[6]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_17[5]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_17[4]))) | ((return_add_generic_AC_RND_CONV_false_14_op_smaller_qr_51_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_17[3]))) | (return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx6
      & (~ (z_out_17[2])));
  assign return_add_generic_AC_RND_CONV_false_14_if_5_or_nl = return_add_generic_AC_RND_CONV_false_14_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_14_mux_16_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_14_if_5_or_nl, z_out_6[53]);
  assign return_add_generic_AC_RND_CONV_false_14_exception_sva_1 = return_add_generic_AC_RND_CONV_false_9_op2_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_9_op2_nan_sva_mx7w0
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_14_mux_16_nl;
  assign return_add_generic_AC_RND_CONV_false_14_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_14_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_14_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_14_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_5 = MUX_v_6_2_2((stage_PE_1_tmp_re_d_1_sva_1_63_57[5:0]),
      (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w9_10_1[9:4]), inverse_lpi_1_dfm_1);
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_4_1 = MUX_v_4_2_2((stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_0[5:2]),
      (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w9_10_1[3:0]), inverse_lpi_1_dfm_1);
  assign stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0 = MUX_s_1_2_2((stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_0[1]),
      stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w9_0, inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_15_if_5_or_nl = return_add_generic_AC_RND_CONV_false_15_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_15_mux_10_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_15_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_15_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_15_exception_sva_1 = return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_15_mux_10_nl;
  assign return_add_generic_AC_RND_CONV_false_15_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_15_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_mult_generic_AC_RND_CONV_false_3_if_1_aelse_return_mult_generic_AC_RND_CONV_false_3_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_3_if_acc_1_itm_12_1) | (z_out_18[105]);
  assign return_mult_generic_AC_RND_CONV_false_3_e_incr_lpi_3_dfm_2 = ~((~(((z_out_18[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((z_out_18[51]) | return_mult_generic_AC_RND_CONV_false_3_if_1_aelse_return_mult_generic_AC_RND_CONV_false_3_if_1_aelse_or_2))
      | (z_out_18[105]))) | (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_3_zero_m_return_mult_generic_AC_RND_CONV_false_3_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_3_r_zero_return_mult_generic_AC_RND_CONV_false_3_r_zero_nor_mdf_sva_1
      = ~(return_mult_generic_AC_RND_CONV_false_3_op1_zero_sva_1 | and_2332_cse);
  assign return_mult_generic_AC_RND_CONV_false_3_r_nan_sva_1 = return_add_generic_AC_RND_CONV_false_19_op1_nan_sva_1
      | (operator_11_true_return_17_sva & (~ return_extract_24_m_zero_sva)) | (return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1
      & and_2332_cse) | (return_mult_generic_AC_RND_CONV_false_3_op1_zero_sva_1 &
      return_mult_generic_AC_RND_CONV_false_3_op2_inf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_3_exp_ovf_return_mult_generic_AC_RND_CONV_false_3_exp_ovf_or_tmp
      = ((return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[10:1]==10'b1111111111)
      & return_mult_generic_AC_RND_CONV_false_exp_ovf_oif_aelse_nor_cse & return_mult_generic_AC_RND_CONV_false_3_e_incr_lpi_3_dfm_2)
      | (z_out_36[11]);
  assign return_mult_generic_AC_RND_CONV_false_3_lor_lpi_3_dfm_1 = return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1
      | return_mult_generic_AC_RND_CONV_false_3_op2_inf_sva_1 | return_mult_generic_AC_RND_CONV_false_3_exp_ovf_return_mult_generic_AC_RND_CONV_false_3_exp_ovf_or_tmp
      | return_mult_generic_AC_RND_CONV_false_3_r_nan_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_3_return_mult_generic_AC_RND_CONV_false_3_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_3_if_1_and_1_tmp_1 | (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_3_and_2_nl = return_mult_generic_AC_RND_CONV_false_3_if_1_and_1_tmp_1
      & (~ (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_3_res_bef_rnd_3_53_1_lpi_3_dfm_1 =
      MUX1HOT_v_53_3_2((z_out_18[104:52]), (z_out_18[103:51]), (z_out_42[53:1]),
      {return_mult_generic_AC_RND_CONV_false_3_return_mult_generic_AC_RND_CONV_false_3_nor_nl
      , return_mult_generic_AC_RND_CONV_false_3_and_2_nl , (z_out_27[12])});
  assign return_mult_generic_AC_RND_CONV_false_3_op2_inf_sva_1 = operator_11_true_return_17_sva
      & return_extract_24_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_3_op1_zero_sva_1 = return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp
      & return_extract_44_m_zero_return_extract_44_m_zero_nor_tmp;
  assign return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_mux_1_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_3_if_acc_1_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva, z_out_27[12]);
  assign return_mult_generic_AC_RND_CONV_false_3_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_mux_1_nl
      & (~ (z_out_18[105]));
  assign return_extract_44_return_extract_44_or_1_cse_sva_1 = (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_5!=6'b000000)
      | (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_4_1!=4'b0000) | stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0;
  assign return_extract_44_m_zero_return_extract_44_m_zero_nor_tmp = ~(return_extract_15_return_extract_15_nor_cse_sva_mx2
      | stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx2_50 | (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1[49:0]!=50'b00000000000000000000000000000000000000000000000000));
  assign operator_11_true_44_operator_11_true_44_and_tmp = (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_5==6'b111111)
      & (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_4_1==4'b1111) & stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0;
  assign return_add_generic_AC_RND_CONV_false_16_if_7_return_add_generic_AC_RND_CONV_false_16_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_16_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0w0 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[50:0]),
      return_add_generic_AC_RND_CONV_false_16_if_7_return_add_generic_AC_RND_CONV_false_16_if_7_nor_nl);
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0 = MUX_v_51_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_1[50:0]),
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0w0, inverse_lpi_1_dfm_1);
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50 = MUX_s_1_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_1[50]),
      (stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0w0[50]), inverse_lpi_1_dfm_1);
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_16_exception_sva_1);
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5 = MUX_v_6_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_0[5:0]),
      (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1[9:4]), inverse_lpi_1_dfm_1);
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1 = MUX_v_4_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_1[56:53]),
      (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1[3:0]), inverse_lpi_1_dfm_1);
  assign or_351_nl = or_dcpl_289 | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva
      | operator_11_true_return_26_sva | and_dcpl_166;
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_13_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs, or_351_nl);
  assign return_add_generic_AC_RND_CONV_false_16_e_r_return_add_generic_AC_RND_CONV_false_16_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_6_mux_35 & (~ return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_13_nl))
      | return_add_generic_AC_RND_CONV_false_16_exception_sva_1;
  assign stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0 = MUX_s_1_2_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_1[52]),
      return_add_generic_AC_RND_CONV_false_16_e_r_return_add_generic_AC_RND_CONV_false_16_e_r_or_1_nl,
      inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_16_r_nan_or_1_nl = operator_11_true_return_26_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva | return_add_generic_AC_RND_CONV_false_10_unequal_tmp;
  assign and_535_nl = (or_dcpl_289 | and_dcpl_166 | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva
      | or_dcpl_1069) & inverse_lpi_1_dfm_1;
  assign and_542_nl = (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_16_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
      & or_dcpl_431 & (~ return_add_generic_AC_RND_CONV_false_22_op1_inf_sva) & (~(return_add_generic_AC_RND_CONV_false_14_op2_inf_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva | operator_11_true_return_26_sva))
      & and_dcpl_385;
  assign return_add_generic_AC_RND_CONV_false_16_r_nan_mux1h_cse = MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_16_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[51]), (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[51]),
      {and_535_nl , and_542_nl , (~ inverse_lpi_1_dfm_1)});
  assign return_add_generic_AC_RND_CONV_false_16_if_5_or_nl = return_add_generic_AC_RND_CONV_false_16_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_16_mux_10_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_16_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_16_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_16_exception_sva_1 = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_inf_sva | operator_11_true_return_26_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva | return_add_generic_AC_RND_CONV_false_16_mux_10_nl;
  assign return_add_generic_AC_RND_CONV_false_16_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_16_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_19_op2_mu_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_extract_45_return_extract_45_or_1_cse_sva_1,
      return_add_generic_AC_RND_CONV_false_16_r_nan_mux1h_cse, return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_16_r_nan_mux1h_cse,
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50, return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0_mx0 =
      MUX_v_50_2_2((stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0[50:1]), (stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0[49:0]),
      return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_19_op2_mu_0_lpi_3_dfm_1 = (stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0[0])
      & (~ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_50_mx0
      = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm,
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50_mx0, and_dcpl_348);
  assign return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0
      = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm,
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0_mx0, and_dcpl_348);
  assign return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_0_lpi_3_dfm_mx0 =
      MUX_s_1_2_2(drf_qr_lval_13_smx_0_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_19_op2_mu_0_lpi_3_dfm_1,
      and_dcpl_348);
  assign return_add_generic_AC_RND_CONV_false_19_e1_eq_e2_equal_tmp = ({BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_1
      , reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd , reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1
      , reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2 , reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3})
      == ({stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5 , stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1
      , stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0});
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_mux_1_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_19_op2_mu_52_lpi_3_dfm_mx0, and_dcpl_348);
  assign return_add_generic_AC_RND_CONV_false_19_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_11_op_smaller_mux_1_nl
      & (~ (z_out_16[54]))) | (return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_50_mx0
      & (~ (z_out_16[53]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[49])
      & (~ (z_out_16[52]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[48])
      & (~ (z_out_16[51]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[47])
      & (~ (z_out_16[50]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[46])
      & (~ (z_out_16[49]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[45])
      & (~ (z_out_16[48]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[44])
      & (~ (z_out_16[47]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[43])
      & (~ (z_out_16[46]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[42])
      & (~ (z_out_16[45]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[41])
      & (~ (z_out_16[44]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[40])
      & (~ (z_out_16[43]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[39])
      & (~ (z_out_16[42]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[38])
      & (~ (z_out_16[41]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[37])
      & (~ (z_out_16[40]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[36])
      & (~ (z_out_16[39]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[35])
      & (~ (z_out_16[38]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[34])
      & (~ (z_out_16[37]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[33])
      & (~ (z_out_16[36]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[32])
      & (~ (z_out_16[35]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[31])
      & (~ (z_out_16[34]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[30])
      & (~ (z_out_16[33]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[29])
      & (~ (z_out_16[32]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[28])
      & (~ (z_out_16[31]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[27])
      & (~ (z_out_16[30]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[26])
      & (~ (z_out_16[29]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[25])
      & (~ (z_out_16[28]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[24])
      & (~ (z_out_16[27]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[23])
      & (~ (z_out_16[26]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[22])
      & (~ (z_out_16[25]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[21])
      & (~ (z_out_16[24]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[20])
      & (~ (z_out_16[23]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[19])
      & (~ (z_out_16[22]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[18])
      & (~ (z_out_16[21]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[17])
      & (~ (z_out_16[20]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[16])
      & (~ (z_out_16[19]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[15])
      & (~ (z_out_16[18]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[14])
      & (~ (z_out_16[17]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[13])
      & (~ (z_out_16[16]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[12])
      & (~ (z_out_16[15]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[11])
      & (~ (z_out_16[14]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[10])
      & (~ (z_out_16[13]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[9])
      & (~ (z_out_16[12]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[8])
      & (~ (z_out_16[11]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[7])
      & (~ (z_out_16[10]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[6])
      & (~ (z_out_16[9]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[5])
      & (~ (z_out_16[8]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[4])
      & (~ (z_out_16[7]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[3])
      & (~ (z_out_16[6]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[2])
      & (~ (z_out_16[5]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[1])
      & (~ (z_out_16[4]))) | ((return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_51_1_lpi_3_dfm_49_0_mx0[0])
      & (~ (z_out_16[3]))) | (return_add_generic_AC_RND_CONV_false_19_op_smaller_qr_0_lpi_3_dfm_mx0
      & (~ (z_out_16[2])));
  assign return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_4_if_acc_1_itm_12_1) | (z_out_18[105]);
  assign return_mult_generic_AC_RND_CONV_false_4_e_incr_lpi_3_dfm_2 = ~((~(((z_out_18[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((z_out_18[51]) | return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_or_2))
      | (z_out_18[105]))) | (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_4_zero_m_return_mult_generic_AC_RND_CONV_false_4_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_4_r_zero_return_mult_generic_AC_RND_CONV_false_4_r_zero_nor_mdf_sva_1
      = ~(return_mult_generic_AC_RND_CONV_false_4_op1_zero_sva_1 | return_mult_generic_AC_RND_CONV_false_4_op2_zero_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_4_r_nan_sva_1 = return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1
      | (operator_11_true_return_24_sva & (~ return_extract_1_m_zero_sva)) | (return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1
      & return_mult_generic_AC_RND_CONV_false_4_op2_zero_sva_1) | (return_mult_generic_AC_RND_CONV_false_4_op1_zero_sva_1
      & return_mult_generic_AC_RND_CONV_false_4_op2_inf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_4_exp_ovf_return_mult_generic_AC_RND_CONV_false_4_exp_ovf_or_tmp
      = ((return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[10:1]==10'b1111111111)
      & return_mult_generic_AC_RND_CONV_false_exp_ovf_oif_aelse_nor_cse & return_mult_generic_AC_RND_CONV_false_4_e_incr_lpi_3_dfm_2)
      | (z_out_36[11]);
  assign return_mult_generic_AC_RND_CONV_false_4_lor_lpi_3_dfm_1 = return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1
      | return_mult_generic_AC_RND_CONV_false_4_op2_inf_sva_1 | return_mult_generic_AC_RND_CONV_false_4_exp_ovf_return_mult_generic_AC_RND_CONV_false_4_exp_ovf_or_tmp
      | return_mult_generic_AC_RND_CONV_false_4_r_nan_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_4_return_mult_generic_AC_RND_CONV_false_4_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_4_if_1_and_1_tmp_1 | (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_4_and_2_nl = return_mult_generic_AC_RND_CONV_false_4_if_1_and_1_tmp_1
      & (~ (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_4_res_bef_rnd_3_53_1_lpi_3_dfm_1 =
      MUX1HOT_v_53_3_2((z_out_18[104:52]), (z_out_18[103:51]), (z_out_42[53:1]),
      {return_mult_generic_AC_RND_CONV_false_4_return_mult_generic_AC_RND_CONV_false_4_nor_nl
      , return_mult_generic_AC_RND_CONV_false_4_and_2_nl , (z_out_27[12])});
  assign return_mult_generic_AC_RND_CONV_false_4_op2_inf_sva_1 = operator_11_true_return_24_sva
      & return_extract_1_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_4_op1_zero_sva_1 = return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_tmp
      & return_extract_45_m_zero_return_extract_45_m_zero_nor_tmp;
  assign return_mult_generic_AC_RND_CONV_false_4_op2_zero_sva_1 = return_extract_17_return_extract_17_nor_cse_sva
      & return_extract_1_m_zero_sva;
  assign return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_mux_1_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_4_if_acc_1_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva, z_out_27[12]);
  assign return_mult_generic_AC_RND_CONV_false_4_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_mux_1_nl
      & (~ (z_out_18[105]));
  assign return_extract_45_return_extract_45_or_1_cse_sva_1 = (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5!=6'b000000)
      | (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1!=4'b0000) | stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0;
  assign return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_1_return_add_generic_AC_RND_CONV_false_19_op2_normal_return_extract_45_nor_tmp
      = ~((stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5!=6'b000000) | (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1!=4'b0000)
      | stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0);
  assign return_extract_45_m_zero_return_extract_45_m_zero_nor_tmp = ~(return_add_generic_AC_RND_CONV_false_16_r_nan_mux1h_cse
      | stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx1_50 | (stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0[49:0]!=50'b00000000000000000000000000000000000000000000000000));
  assign operator_11_true_45_operator_11_true_45_and_tmp = (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5==6'b111111)
      & (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1==4'b1111) & stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0;
  assign return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_49_0,
      return_add_generic_AC_RND_CONV_false_20_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_264);
  assign return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_5_if_acc_1_itm_12_1) | (z_out_18[105]);
  assign return_mult_generic_AC_RND_CONV_false_5_e_incr_lpi_3_dfm_2 = ~((~(((z_out_18[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((z_out_18[51]) | return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_or_2))
      | (z_out_18[105]))) | (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_5_zero_m_return_mult_generic_AC_RND_CONV_false_5_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_5_r_zero_return_mult_generic_AC_RND_CONV_false_5_r_zero_nor_mdf_sva_1
      = ~(return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 | (return_extract_51_return_extract_51_nor_tmp
      & return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp));
  assign return_mult_generic_AC_RND_CONV_false_5_else_2_else_else_mux_nl = MUX_v_11_2_2((return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[10:0]),
      (z_out_36[10:0]), return_mult_generic_AC_RND_CONV_false_5_e_incr_lpi_3_dfm_2);
  assign return_mult_generic_AC_RND_CONV_false_5_else_2_else_return_mult_generic_AC_RND_CONV_false_5_else_2_else_and_nl
      = MUX_v_11_2_2(11'b00000000000, return_mult_generic_AC_RND_CONV_false_5_else_2_else_else_mux_nl,
      return_mult_generic_AC_RND_CONV_false_5_zero_m_return_mult_generic_AC_RND_CONV_false_5_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_5_r_zero_return_mult_generic_AC_RND_CONV_false_5_r_zero_nor_mdf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1 =
      MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_5_else_2_else_return_mult_generic_AC_RND_CONV_false_5_else_2_else_and_nl,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_5_lor_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[0])
      & operator_11_true_return_15_sva;
  assign return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1 = return_mult_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_mx1
      | return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp;
  assign return_add_generic_AC_RND_CONV_false_20_op2_mu_1_51_lpi_3_dfm_mx0 = MUX_s_1_2_2((return_mult_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[50]),
      return_mult_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_mx1, return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp);
  assign return_add_generic_AC_RND_CONV_false_20_op2_mu_1_50_1_lpi_3_dfm_mx0 = MUX_v_50_2_2((return_mult_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[49:0]),
      (return_mult_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[50:1]), return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp);
  assign return_add_generic_AC_RND_CONV_false_20_op2_mu_1_0_lpi_3_dfm_1 = (return_mult_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1[0])
      & return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp;
  assign and_546_nl = return_mult_generic_AC_RND_CONV_false_5_zero_m_return_mult_generic_AC_RND_CONV_false_5_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_5_r_zero_return_mult_generic_AC_RND_CONV_false_5_r_zero_nor_mdf_sva_1
      & (~(operator_11_true_51_operator_11_true_51_and_tmp | (z_out_36[11]) | return_mult_generic_AC_RND_CONV_false_5_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_5_exp_ovf_oif_aelse_and_tmp));
  assign return_mult_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_mx1 = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_5_r_nan_sva_1,
      (z_out_6[51]), and_546_nl);
  assign return_mult_generic_AC_RND_CONV_false_5_oelse_3_return_mult_generic_AC_RND_CONV_false_5_if_3_nor_nl
      = ~((~ return_mult_generic_AC_RND_CONV_false_5_zero_m_return_mult_generic_AC_RND_CONV_false_5_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_5_r_zero_return_mult_generic_AC_RND_CONV_false_5_r_zero_nor_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_5_lor_lpi_3_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (z_out_6[50:0]), return_mult_generic_AC_RND_CONV_false_5_oelse_3_return_mult_generic_AC_RND_CONV_false_5_if_3_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_20_e1_eq_e2_equal_tmp = ({BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1
      , reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd , reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1})
      == (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1);
  assign return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[0])
      & return_add_generic_AC_RND_CONV_false_10_do_sub_sva;
  assign return_add_generic_AC_RND_CONV_false_21_e1_eq_e2_equal_tmp = ({BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1
      , BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2}) == (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1);
  assign return_add_generic_AC_RND_CONV_false_20_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_52_lpi_3_dfm_mx3
      & (~ (z_out_16[54]))) | (return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_51_lpi_3_dfm_mx3
      & (~ (z_out_16[53]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_16[52]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_16[51]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_16[50]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_16[49]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_16[48]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_16[47]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_16[46]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_16[45]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_16[44]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_16[43]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_16[42]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_16[41]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_16[40]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_16[39]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_16[38]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_16[37]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_16[36]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_16[35]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_16[34]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_16[33]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_16[32]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_16[31]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_16[30]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_16[29]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_16[28]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_16[27]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_16[26]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_16[25]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_16[24]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_16[23]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_16[22]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_16[21]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_16[20]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_16[19]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_16[18]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_16[17]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_16[16]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_16[15]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_16[14]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_16[13]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_16[12]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_16[11]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_16[10]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_16[9]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_16[8]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_16[7]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_16[6]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_16[5]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_16[4]))) | ((return_add_generic_AC_RND_CONV_false_20_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_16[3]))) | (return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm_mx4
      & (~ (z_out_16[2])));
  assign return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_1_tmp
      = (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1!=11'b00000000000);
  assign return_mult_generic_AC_RND_CONV_false_5_r_nan_sva_1 = (operator_11_true_51_operator_11_true_51_and_tmp
      & (~ return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp)) | (return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1
      & return_mult_generic_AC_RND_CONV_false_5_op2_inf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_5_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_5_exp_ovf_oif_aelse_and_tmp
      = (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1[10:1]==10'b1111111111)
      & return_mult_generic_AC_RND_CONV_false_exp_ovf_oif_aelse_nor_cse & return_mult_generic_AC_RND_CONV_false_5_e_incr_lpi_3_dfm_2;
  assign return_mult_generic_AC_RND_CONV_false_5_lor_lpi_3_dfm_1 = return_mult_generic_AC_RND_CONV_false_5_op2_inf_sva_1
      | return_mult_generic_AC_RND_CONV_false_5_exp_ovf_oif_aif_return_mult_generic_AC_RND_CONV_false_5_exp_ovf_oif_aelse_and_tmp
      | (z_out_36[11]) | return_mult_generic_AC_RND_CONV_false_5_r_nan_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_5_return_mult_generic_AC_RND_CONV_false_5_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_5_if_1_and_1_tmp_1 | (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_5_and_2_nl = return_mult_generic_AC_RND_CONV_false_5_if_1_and_1_tmp_1
      & (~ (z_out_27[12]));
  assign return_mult_generic_AC_RND_CONV_false_5_res_bef_rnd_3_53_1_lpi_3_dfm_1 =
      MUX1HOT_v_53_3_2((z_out_18[104:52]), (z_out_18[103:51]), (z_out_42[53:1]),
      {return_mult_generic_AC_RND_CONV_false_5_return_mult_generic_AC_RND_CONV_false_5_nor_nl
      , return_mult_generic_AC_RND_CONV_false_5_and_2_nl , (z_out_27[12])});
  assign return_mult_generic_AC_RND_CONV_false_5_op2_inf_sva_1 = operator_11_true_51_operator_11_true_51_and_tmp
      & return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp;
  assign return_extract_51_return_extract_51_nor_tmp = ~((return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1);
  assign return_extract_51_m_zero_return_extract_51_m_zero_nor_tmp = ~(return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_mux_1_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_5_if_acc_1_itm_12_1,
      return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva, z_out_27[12]);
  assign return_mult_generic_AC_RND_CONV_false_5_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_mux_1_nl
      & (~ (z_out_18[105]));
  assign return_extract_51_return_extract_51_or_sva_1 = (return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1;
  assign and_551_nl = (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
      & or_dcpl_431 & and_dcpl_399 & (~(return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva));
  assign return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_15_r_nan_or_mx2w0,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[51]), and_551_nl);
  assign return_add_generic_AC_RND_CONV_false_19_if_7_return_add_generic_AC_RND_CONV_false_19_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_19_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[50:0]),
      return_add_generic_AC_RND_CONV_false_19_if_7_return_add_generic_AC_RND_CONV_false_19_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_19_exception_sva_1);
  assign or_358_nl = or_dcpl_296 | or_dcpl_275 | and_dcpl_166;
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_15_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs, or_358_nl);
  assign return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_6_mux_35
      & (~ return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_15_nl)) | return_add_generic_AC_RND_CONV_false_19_exception_sva_1;
  assign operator_11_true_51_operator_11_true_51_and_tmp = (return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_19_if_5_or_nl = return_add_generic_AC_RND_CONV_false_19_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_19_mux_16_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_19_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_19_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_19_exception_sva_1 = return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_19_mux_16_nl;
  assign return_add_generic_AC_RND_CONV_false_19_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49:0]),
      return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_265);
  assign return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_20_exception_sva_1);
  assign or_364_nl = or_dcpl_302 | or_dcpl_235;
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_17_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs, or_364_nl);
  assign return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_6_mux_35
      & (~ return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_17_nl)) | return_add_generic_AC_RND_CONV_false_20_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_20_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_22_op2_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_22_op2_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_16_do_sub_sva);
  assign and_554_nl = (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_20_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
      & or_dcpl_431 & and_dcpl_408;
  assign return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_20_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[51]), and_554_nl);
  assign return_add_generic_AC_RND_CONV_false_20_if_7_return_add_generic_AC_RND_CONV_false_20_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_20_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[50:0]),
      return_add_generic_AC_RND_CONV_false_20_if_7_return_add_generic_AC_RND_CONV_false_20_if_7_nor_nl);
  assign return_extract_57_return_extract_57_or_2_nl = (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_extract_57_return_extract_57_or_2_nl,
      return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1[50]), return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0 = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1[50:1]),
      (return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1[49:0]), return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1[0])
      & (~ return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_22_e1_eq_e2_equal_tmp = (stage_PE_1_x_re_d_sva[62:52])
      == ({return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1});
  assign return_add_generic_AC_RND_CONV_false_22_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_22_op1_mu_mux_1_cse
      & (~ (z_out_17[54]))) | (return_add_generic_AC_RND_CONV_false_5_op_smaller_mux_cse
      & (~ (z_out_17[53]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_17[52]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_17[51]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_17[50]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_17[49]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_17[48]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_17[47]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_17[46]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_17[45]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_17[44]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_17[43]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_17[42]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_17[41]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_17[40]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_17[39]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_17[38]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_17[37]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_17[36]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_17[35]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_17[34]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_17[33]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_17[32]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_17[31]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_17[30]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_17[29]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_17[28]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_17[27]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_17[26]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_17[25]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_17[24]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_17[23]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_17[22]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_17[21]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_17[20]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_17[19]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_17[18]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_17[17]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_17[16]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_17[15]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_17[14]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_17[13]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_17[12]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_17[11]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_17[10]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_17[9]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_17[8]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_17[7]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_17[6]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_17[5]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_17[4]))) | ((return_add_generic_AC_RND_CONV_false_22_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_17[3]))) | (return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_3_cse
      & (~ (z_out_17[2])));
  assign return_add_generic_AC_RND_CONV_false_22_return_add_generic_AC_RND_CONV_false_22_if_1_return_add_generic_AC_RND_CONV_false_22_op2_normal_return_extract_57_nor_tmp
      = ~((return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_20_if_5_or_nl = return_add_generic_AC_RND_CONV_false_20_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_20_mux_18_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_20_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_20_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_20_exception_sva_1 = return_add_generic_AC_RND_CONV_false_22_op2_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_22_op2_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_20_mux_18_nl;
  assign return_add_generic_AC_RND_CONV_false_20_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_20_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_3_e_r_qelse_qr_10_1_lpi_3_dfm_1,
      10'b1111111111, return_add_generic_AC_RND_CONV_false_21_exception_sva_1);
  assign or_368_nl = return_add_generic_AC_RND_CONV_false_21_r_inf_lpi_3_dfm_2 |
      return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | or_dcpl_244;
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_19_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs, or_368_nl);
  assign return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_6_mux_35
      & (~ return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_19_nl)) | return_add_generic_AC_RND_CONV_false_21_exception_sva_1;
  assign return_add_generic_AC_RND_CONV_false_21_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_21_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | (return_add_generic_AC_RND_CONV_false_21_op1_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva & return_add_generic_AC_RND_CONV_false_14_op2_inf_sva);
  assign and_557_nl = (~((~((~ (operator_33_true_12_acc_psp_sva[11])) & return_add_generic_AC_RND_CONV_false_21_else_4_unequal_tmp))
      & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva))
      & or_dcpl_431 & and_dcpl_413;
  assign return_add_generic_AC_RND_CONV_false_21_m_r_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_r_nan_or_1_nl,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[51]), and_557_nl);
  assign return_add_generic_AC_RND_CONV_false_21_if_7_return_add_generic_AC_RND_CONV_false_21_if_7_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_21_exception_sva_1 | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1 = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      (return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0[50:0]),
      return_add_generic_AC_RND_CONV_false_21_if_7_return_add_generic_AC_RND_CONV_false_21_if_7_nor_nl);
  assign return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0 = MUX_v_12_2_2(z_out_25,
      z_out_23, z_out_25[11]);
  assign return_extract_59_return_extract_59_or_2_nl = (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_extract_59_return_extract_59_or_2_nl,
      return_add_generic_AC_RND_CONV_false_21_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_m_r_51_lpi_3_dfm_mx0,
      (return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1[50]), return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0 = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1[50:1]),
      (return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1[49:0]), return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1 = (return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1[0])
      & (~ return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp);
  assign return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0
      = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[49:0]),
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0, and_dcpl_266);
  assign return_add_generic_AC_RND_CONV_false_23_e1_eq_e2_equal_tmp = (stage_PE_1_x_im_d_sva[62:52])
      == ({return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1 , return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1});
  assign return_add_generic_AC_RND_CONV_false_23_res_mant_3_0_sva_1 = (return_add_generic_AC_RND_CONV_false_13_mux_25_cse
      & (~ (z_out_16[54]))) | (return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_2_cse
      & (~ (z_out_16[53]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[49])
      & (~ (z_out_16[52]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[48])
      & (~ (z_out_16[51]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[47])
      & (~ (z_out_16[50]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[46])
      & (~ (z_out_16[49]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[45])
      & (~ (z_out_16[48]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[44])
      & (~ (z_out_16[47]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[43])
      & (~ (z_out_16[46]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[42])
      & (~ (z_out_16[45]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[41])
      & (~ (z_out_16[44]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[40])
      & (~ (z_out_16[43]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[39])
      & (~ (z_out_16[42]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[38])
      & (~ (z_out_16[41]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[37])
      & (~ (z_out_16[40]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[36])
      & (~ (z_out_16[39]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[35])
      & (~ (z_out_16[38]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[34])
      & (~ (z_out_16[37]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[33])
      & (~ (z_out_16[36]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[32])
      & (~ (z_out_16[35]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[31])
      & (~ (z_out_16[34]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[30])
      & (~ (z_out_16[33]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[29])
      & (~ (z_out_16[32]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[28])
      & (~ (z_out_16[31]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[27])
      & (~ (z_out_16[30]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[26])
      & (~ (z_out_16[29]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[25])
      & (~ (z_out_16[28]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[24])
      & (~ (z_out_16[27]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[23])
      & (~ (z_out_16[26]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[22])
      & (~ (z_out_16[25]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[21])
      & (~ (z_out_16[24]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[20])
      & (~ (z_out_16[23]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[19])
      & (~ (z_out_16[22]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[18])
      & (~ (z_out_16[21]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[17])
      & (~ (z_out_16[20]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[16])
      & (~ (z_out_16[19]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[15])
      & (~ (z_out_16[18]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[14])
      & (~ (z_out_16[17]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[13])
      & (~ (z_out_16[16]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[12])
      & (~ (z_out_16[15]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[11])
      & (~ (z_out_16[14]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[10])
      & (~ (z_out_16[13]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[9])
      & (~ (z_out_16[12]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[8])
      & (~ (z_out_16[11]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[7])
      & (~ (z_out_16[10]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[6])
      & (~ (z_out_16[9]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[5])
      & (~ (z_out_16[8]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[4])
      & (~ (z_out_16[7]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[3])
      & (~ (z_out_16[6]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[2])
      & (~ (z_out_16[5]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[1])
      & (~ (z_out_16[4]))) | ((return_add_generic_AC_RND_CONV_false_23_op_smaller_qr_50_1_lpi_3_dfm_mx0[0])
      & (~ (z_out_16[3]))) | (return_add_generic_AC_RND_CONV_false_1_op_bigger_mux_5_cse
      & (~ (z_out_16[2])));
  assign return_add_generic_AC_RND_CONV_false_25_e_dif_qr_lpi_3_dfm_mx0_10_0 = MUX_v_11_2_2((z_out_25[10:0]),
      (z_out_23[10:0]), z_out_25[11]);
  assign return_add_generic_AC_RND_CONV_false_23_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0[11:6]!=6'b000000);
  assign return_add_generic_AC_RND_CONV_false_23_e_dif_sat_sva_1 = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_23_e_dif_qr_lpi_3_dfm_mx0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_23_e_dif_sat_or_1_nl);
  assign return_add_generic_AC_RND_CONV_false_23_return_add_generic_AC_RND_CONV_false_23_if_1_return_add_generic_AC_RND_CONV_false_23_op2_normal_return_extract_59_nor_tmp
      = ~((return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_21_op1_nan_sva_1 = operator_11_true_return_17_sva
      & (~ return_extract_15_m_zero_sva);
  assign return_add_generic_AC_RND_CONV_false_21_op1_inf_sva_1 = operator_11_true_return_17_sva
      & return_extract_15_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_21_if_5_or_nl = return_add_generic_AC_RND_CONV_false_21_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_21_mux_14_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_21_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_21_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_21_exception_sva_1 = return_add_generic_AC_RND_CONV_false_21_op1_inf_sva_1
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_21_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_21_mux_14_nl;
  assign return_add_generic_AC_RND_CONV_false_21_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_21_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_25_res_mant_3_0_sva_1 = return_add_generic_AC_RND_CONV_false_12_sticky_bit_and_54
      | return_add_generic_AC_RND_CONV_false_12_sticky_bit_and_56 | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_2_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_3_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_4_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_5_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_6_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_7_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_8_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_9_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_10_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_11_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_12_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_13_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_14_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_15_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_16_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_17_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_18_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_19_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_20_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_21_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_22_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_23_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_24_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_25_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_26_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_27_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_28_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_29_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_30_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_31_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_32_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_33_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_34_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_35_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_36_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_37_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_38_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_39_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_40_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_41_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_42_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_43_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_44_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_45_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_46_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_47_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_48_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_49_cse | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_50_cse
      | return_add_generic_AC_RND_CONV_false_11_sticky_bit_and_51_cse | return_add_generic_AC_RND_CONV_false_12_sticky_bit_and_58;
  assign return_add_generic_AC_RND_CONV_false_22_if_5_or_nl = return_add_generic_AC_RND_CONV_false_22_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_22_mux_17_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_22_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_22_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_22_exception_sva_1 = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_22_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_22_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_22_mux_17_nl;
  assign return_add_generic_AC_RND_CONV_false_22_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_22_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_22_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_22_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_23_if_5_or_nl = return_add_generic_AC_RND_CONV_false_23_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_23_mux_17_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_23_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_23_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_23_exception_sva_1 = return_add_generic_AC_RND_CONV_false_23_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1 | return_add_generic_AC_RND_CONV_false_23_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | return_add_generic_AC_RND_CONV_false_23_mux_17_nl;
  assign return_add_generic_AC_RND_CONV_false_23_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_23_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_23_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_23_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_24_if_5_or_nl = return_add_generic_AC_RND_CONV_false_24_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_24_mux_10_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_24_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_24_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_24_exception_sva_1 = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_24_mux_10_nl;
  assign return_add_generic_AC_RND_CONV_false_24_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_24_exception_sva_1
      | operator_11_true_return_24_sva;
  assign return_add_generic_AC_RND_CONV_false_24_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_24_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_25_if_5_or_nl = return_add_generic_AC_RND_CONV_false_25_r_inf_lpi_3_dfm_2
      | return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign return_add_generic_AC_RND_CONV_false_25_mux_10_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_25_r_inf_lpi_3_dfm_2,
      return_add_generic_AC_RND_CONV_false_25_if_5_or_nl, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_25_exception_sva_1 = return_add_generic_AC_RND_CONV_false_23_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_inf_sva | return_add_generic_AC_RND_CONV_false_23_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva | return_add_generic_AC_RND_CONV_false_25_mux_10_nl;
  assign return_add_generic_AC_RND_CONV_false_25_or_1_svs_1 = return_add_generic_AC_RND_CONV_false_25_exception_sva_1
      | return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva;
  assign return_add_generic_AC_RND_CONV_false_25_r_inf_lpi_3_dfm_2 = ((operator_33_true_12_acc_psp_sva[11])
      | (~ return_add_generic_AC_RND_CONV_false_25_else_4_unequal_tmp)) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_or_2
      = (~ return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1) | (z_out_18[105]);
  assign return_mult_generic_AC_RND_CONV_false_6_if_if_not_nl = ~ (z_out_29[11]);
  assign return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3 = MUX_v_11_2_2(11'b00000000000,
      (z_out_29[10:0]), return_mult_generic_AC_RND_CONV_false_6_if_if_not_nl);
  assign return_mult_generic_AC_RND_CONV_false_6_e_incr_lpi_2_dfm_2 = ~((~(((z_out_18[104:52]==53'b11111111111111111111111111111111111111111111111111111)
      & ((z_out_18[51]) | return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_or_2))
      | (z_out_18[105]))) | (z_out_27[11]));
  assign return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1
      = ~((out_f_d_rsci_q_d[62:52]==11'b00000000000) & return_extract_3_m_zero_sva_mx1w0);
  assign return_mult_generic_AC_RND_CONV_false_6_lor_lpi_2_dfm_1 = (operator_11_true_24_operator_11_true_24_and_tmp
      & return_extract_3_m_zero_sva_mx1w0) | ((return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3==11'b11111111110)
      & return_mult_generic_AC_RND_CONV_false_6_e_incr_lpi_2_dfm_2) | return_mult_generic_AC_RND_CONV_false_6_op1_nan_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_6_op1_nan_sva_1 = operator_11_true_24_operator_11_true_24_and_tmp
      & (~ return_extract_3_m_zero_sva_mx1w0);
  assign return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1 = (~ return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1)
      | return_mult_generic_AC_RND_CONV_false_6_lor_lpi_2_dfm_1;
  assign return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_nor_nl
      = ~(return_mult_generic_AC_RND_CONV_false_6_if_1_and_1_tmp_1 | (z_out_27[11]));
  assign return_mult_generic_AC_RND_CONV_false_6_and_2_nl = return_mult_generic_AC_RND_CONV_false_6_if_1_and_1_tmp_1
      & (~ (z_out_27[11]));
  assign return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1 =
      MUX1HOT_v_53_3_2((z_out_18[104:52]), (z_out_18[103:51]), (z_out_42[53:1]),
      {return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_nor_nl
      , return_mult_generic_AC_RND_CONV_false_6_and_2_nl , (z_out_27[11])});
  assign return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_mux_1_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1,
      return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva, z_out_27[11]);
  assign return_mult_generic_AC_RND_CONV_false_6_if_1_and_1_tmp_1 = return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_mux_1_nl
      & (~ (z_out_18[105]));
  assign nl_stage_monty_mul_acc_2_psp_sva_1 = operator_32_false_2_acc_psp_1_sva_1
      + conv_u2s_14_15(signext_14_13({(operator_32_false_2_acc_psp_1_sva_1[14]) ,
      11'b00000000000 , (operator_32_false_2_acc_psp_1_sva_1[14])}));
  assign stage_monty_mul_acc_2_psp_sva_1 = nl_stage_monty_mul_acc_2_psp_sva_1[14:0];
  assign nl_operator_32_false_2_acc_psp_1_sva_1 = conv_u2s_14_15(z_out_30[23:10])
      + 15'b100111111111111;
  assign operator_32_false_2_acc_psp_1_sva_1 = nl_operator_32_false_2_acc_psp_1_sva_1[14:0];
  assign return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_9
      = (operator_33_true_12_acc_psp_sva[0]) & return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva;
  assign return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_11
      = MUX_v_10_2_2(10'b0000000000, (operator_33_true_12_acc_psp_sva[10:1]), return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva);
  assign return_add_generic_AC_RND_CONV_false_if_5_or_3 = return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva
      | (~((operator_33_true_12_acc_psp_sva!=13'b0000000000000)));
  assign return_add_generic_AC_RND_CONV_false_mux_28 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva,
      return_add_generic_AC_RND_CONV_false_if_5_or_3, reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_5_sticky_bit_and_54 = return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm
      & (~ (z_out_16[2]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_54 = return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm
      & (~ (z_out_16[54]));
  assign return_add_generic_AC_RND_CONV_false_8_sticky_bit_and_56 = return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm
      & (~ (z_out_16[53]));
  assign nl_return_add_generic_AC_RND_CONV_false_18_acc_3_nl =  -(z_out_37[10:0]);
  assign return_add_generic_AC_RND_CONV_false_18_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_18_acc_3_nl[10:0];
  assign return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1 = readslicef_11_1_10(return_add_generic_AC_RND_CONV_false_18_acc_3_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_20_acc_3_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_20_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_20_acc_3_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_20_acc_3_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_20_acc_3_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_8_acc_3_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_8_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_8_acc_3_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_8_acc_3_nl);
  assign nl_return_add_generic_AC_RND_CONV_false_19_acc_3_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_19_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_19_acc_3_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_19_acc_3_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_19_acc_3_nl);
  assign return_add_generic_AC_RND_CONV_false_6_mux_35 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_9,
      return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_or_2_cse,
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign nl_return_add_generic_AC_RND_CONV_false_15_acc_3_nl =  -(z_out_8[11:0]);
  assign return_add_generic_AC_RND_CONV_false_15_acc_3_nl = nl_return_add_generic_AC_RND_CONV_false_15_acc_3_nl[11:0];
  assign return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1 = readslicef_12_1_11(return_add_generic_AC_RND_CONV_false_15_acc_3_nl);
  assign return_add_generic_AC_RND_CONV_false_19_if_2_return_add_generic_AC_RND_CONV_false_19_if_2_nor_2
      = ~(stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0 | (~ return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm));
  assign return_add_generic_AC_RND_CONV_false_12_sticky_bit_and_54 = return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_52_lpi_3_dfm
      & (~ (z_out_16[54]));
  assign return_add_generic_AC_RND_CONV_false_12_sticky_bit_and_56 = return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_51_lpi_3_dfm
      & (~ (z_out_16[53]));
  assign return_add_generic_AC_RND_CONV_false_12_sticky_bit_and_58 = return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm
      & (~ (z_out_16[2]));
  assign return_add_generic_AC_RND_CONV_false_1_mux_32 = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_9,
      return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_or_2_cse,
      z_out_6[53]);
  assign return_add_generic_AC_RND_CONV_false_15_aif_equal_tmp = ({return_add_generic_AC_RND_CONV_false_13_op1_mu_52_lpi_3_dfm_1
      , return_extract_32_mux_4_cse , return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1})
      == ({drf_qr_lval_13_smx_0_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1});
  assign or_dcpl_11 = (fsm_output[54:53]!=2'b00);
  assign and_dcpl_1 = (~ inverse_lpi_1_dfm_1) & mode_lpi_1_dfm;
  assign or_38_cse = (fsm_output[29]) | (fsm_output[4]);
  assign nor_3_cse = ~(inverse_lpi_1_dfm_1 | mode_lpi_1_dfm);
  assign or_dcpl_48 = ~(nand_12_cse & return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1);
  assign and_dcpl_28 = ~(return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva);
  assign or_dcpl_49 = ~(nand_12_cse & return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1);
  assign and_dcpl_32 = (~ return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva) &
      mode_lpi_1_dfm;
  assign and_dcpl_36 = (~(nand_12_cse & return_add_generic_AC_RND_CONV_false_19_acc_3_itm_11_1))
      & and_dcpl_28;
  assign and_dcpl_63 = ~(return_add_generic_AC_RND_CONV_false_10_op1_nan_sva | return_add_generic_AC_RND_CONV_false_10_op1_inf_sva);
  assign and_2334_cse = BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm & mode_lpi_1_dfm;
  assign nor_158_cse = ~(and_2334_cse | (BUTTERFLY_1_n_9_0_sva_1[9]));
  assign nor_24_cse = ~((fsm_output[52]) | (fsm_output[27]));
  assign and_dcpl_128 = ~((operator_16_false_io_read_mode1_rsc_cse_sva[6:5]!=2'b00));
  assign and_dcpl_129 = and_dcpl_128 & (operator_16_false_io_read_mode1_rsc_cse_sva[4:3]==2'b00);
  assign and_dcpl_135 = ~((operator_16_false_io_read_mode1_rsc_cse_sva[15:14]!=2'b00));
  assign and_dcpl_138 = and_dcpl_135 & (operator_16_false_io_read_mode1_rsc_cse_sva[13:7]==7'b0000000);
  assign or_dcpl_75 = (operator_16_false_io_read_mode1_rsc_cse_sva[3:2]!=2'b00);
  assign or_dcpl_79 = (operator_16_false_io_read_mode1_rsc_cse_sva[7:4]!=4'b0000);
  assign or_dcpl_87 = (operator_16_false_io_read_mode1_rsc_cse_sva[15:8]!=8'b00000000);
  assign and_dcpl_140 = ~((~(or_dcpl_87 | or_dcpl_79 | or_dcpl_75 | (operator_16_false_io_read_mode1_rsc_cse_sva[1:0]!=2'b01)))
      | operator_16_false_operator_16_false_nor_cse_sva);
  assign and_dcpl_146 = ~((~(or_dcpl_87 | or_dcpl_79 | or_dcpl_75 | (~((operator_16_false_io_read_mode1_rsc_cse_sva[1])
      ^ (operator_16_false_io_read_mode1_rsc_cse_sva[0]))))) | operator_16_false_operator_16_false_nor_cse_sva);
  assign or_dcpl_92 = (fsm_output[32:31]!=2'b00);
  assign or_dcpl_95 = (fsm_output[5:4]!=2'b00);
  assign or_dcpl_99 = (fsm_output[34:33]!=2'b00);
  assign or_dcpl_101 = (fsm_output[42:41]!=2'b00);
  assign or_dcpl_102 = (fsm_output[44:43]!=2'b00);
  assign or_dcpl_105 = (fsm_output[49]) | (fsm_output[45]);
  assign or_dcpl_106 = (fsm_output[50]) | (fsm_output[46]);
  assign or_dcpl_108 = (fsm_output[48:47]!=2'b00);
  assign and_dcpl_151 = (operator_16_false_io_read_mode1_rsc_cse_sva[1:0]==2'b01);
  assign and_dcpl_152 = ~((operator_16_false_io_read_mode1_rsc_cse_sva[3:2]!=2'b00));
  assign or_dcpl_115 = (and_dcpl_135 & (operator_16_false_io_read_mode1_rsc_cse_sva[13:4]==10'b0000000000)
      & and_dcpl_152 & and_dcpl_151) | operator_16_false_operator_16_false_nor_cse_sva;
  assign or_dcpl_118 = (fsm_output[30:29]!=2'b00);
  assign or_dcpl_125 = (fsm_output[21:20]!=2'b00);
  assign or_dcpl_126 = (fsm_output[25:24]!=2'b00);
  assign or_dcpl_128 = (fsm_output[23:22]!=2'b00);
  assign or_dcpl_132 = (fsm_output[16]) | (fsm_output[6]);
  assign or_dcpl_133 = (fsm_output[18:17]!=2'b00);
  assign or_dcpl_135 = (fsm_output[9]) | (fsm_output[19]);
  assign or_dcpl_136 = (fsm_output[8:7]!=2'b00);
  assign and_dcpl_165 = ~((fsm_output[56]) | (fsm_output[0]));
  assign or_dcpl_148 = (fsm_output[51]) | (fsm_output[47]);
  assign or_dcpl_159 = (fsm_output[9:8]!=2'b00);
  assign or_dcpl_163 = (fsm_output[7]) | (fsm_output[9]);
  assign or_dcpl_166 = (fsm_output[26]) | (fsm_output[22]);
  assign and_dcpl_166 = reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd
      & return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp;
  assign or_dcpl_185 = ~(inverse_lpi_1_dfm_1 & mode_lpi_1_dfm);
  assign or_dcpl_187 = operator_11_true_return_1_sva | operator_11_true_return_24_sva
      | or_dcpl_185;
  assign and_dcpl_168 = return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp
      & (z_out_6[53]);
  assign or_dcpl_199 = return_add_generic_AC_RND_CONV_false_14_op2_inf_sva | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva;
  assign or_dcpl_201 = return_add_generic_AC_RND_CONV_false_23_op1_inf_sva | return_add_generic_AC_RND_CONV_false_23_op1_nan_sva;
  assign or_dcpl_203 = return_add_generic_AC_RND_CONV_false_2_r_inf_lpi_3_dfm_2 |
      or_dcpl_201;
  assign or_dcpl_207 = or_dcpl_201 | return_add_generic_AC_RND_CONV_false_14_op2_inf_sva;
  assign or_dcpl_211 = ~(return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1 &
      inverse_lpi_1_dfm_1 & mode_lpi_1_dfm);
  assign or_dcpl_214 = return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_10_op2_inf_sva;
  assign or_dcpl_216 = return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2 |
      or_dcpl_214;
  assign or_dcpl_219 = and_dcpl_166 | operator_11_true_return_26_sva | or_dcpl_185;
  assign or_dcpl_224 = ~(return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1 &
      inverse_lpi_1_dfm_1 & mode_lpi_1_dfm);
  assign or_dcpl_225 = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva | return_add_generic_AC_RND_CONV_false_22_op1_inf_sva;
  assign or_dcpl_228 = return_add_generic_AC_RND_CONV_false_6_r_inf_lpi_3_dfm_2 |
      or_dcpl_214;
  assign or_dcpl_231 = and_dcpl_166 | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva;
  assign or_dcpl_234 = ~(return_add_generic_AC_RND_CONV_false_19_acc_3_itm_11_1 &
      mode_lpi_1_dfm);
  assign or_dcpl_235 = and_dcpl_166 | operator_11_true_return_1_sva;
  assign or_dcpl_237 = return_add_generic_AC_RND_CONV_false_7_r_inf_lpi_3_dfm_2 |
      operator_11_true_return_15_sva;
  assign or_dcpl_240 = and_dcpl_166 | operator_11_true_return_1_sva | (~ mode_lpi_1_dfm);
  assign or_dcpl_242 = ~(return_add_generic_AC_RND_CONV_false_20_acc_3_itm_11_1 &
      mode_lpi_1_dfm);
  assign or_dcpl_244 = return_add_generic_AC_RND_CONV_false_10_op2_inf_sva | operator_11_true_return_17_sva
      | and_dcpl_166;
  assign or_dcpl_249 = and_dcpl_166 | operator_11_true_return_17_sva | (~ mode_lpi_1_dfm);
  assign or_dcpl_252 = ~(return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1 &
      mode_lpi_1_dfm);
  assign or_dcpl_261 = operator_11_true_return_15_sva | operator_11_true_return_1_sva;
  assign or_dcpl_275 = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva | return_add_generic_AC_RND_CONV_false_10_op1_inf_sva;
  assign or_dcpl_278 = return_add_generic_AC_RND_CONV_false_15_r_inf_lpi_3_dfm_2
      | or_dcpl_214;
  assign or_dcpl_282 = or_dcpl_214 | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva;
  assign or_dcpl_287 = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva | return_add_generic_AC_RND_CONV_false_14_op2_inf_sva;
  assign or_dcpl_289 = return_add_generic_AC_RND_CONV_false_16_r_inf_lpi_3_dfm_2
      | or_dcpl_287;
  assign or_dcpl_296 = return_add_generic_AC_RND_CONV_false_19_r_inf_lpi_3_dfm_2
      | or_dcpl_214;
  assign or_dcpl_302 = return_add_generic_AC_RND_CONV_false_20_r_inf_lpi_3_dfm_2
      | operator_11_true_return_15_sva;
  assign or_dcpl_395 = (fsm_output[52]) | (fsm_output[27]);
  assign and_dcpl_210 = nor_24_cse & (~ (fsm_output[1]));
  assign and_dcpl_211 = ~((fsm_output[0]) | (fsm_output[53]));
  assign and_dcpl_213 = ~((fsm_output[1]) | (fsm_output[55]));
  assign and_dcpl_214 = and_dcpl_213 & (~ (fsm_output[56]));
  assign and_dcpl_217 = ~((fsm_output[53]) | (fsm_output[54]) | (fsm_output[2]));
  assign or_dcpl_397 = (fsm_output[50]) | (fsm_output[25]);
  assign and_dcpl_233 = nor_24_cse & (~((fsm_output[51]) | (fsm_output[26]))) & and_dcpl_214;
  assign and_dcpl_236 = ~((fsm_output[54]) | (fsm_output[2]));
  assign or_dcpl_401 = (fsm_output[31]) | (fsm_output[6]);
  assign or_dcpl_404 = (fsm_output[37]) | (fsm_output[12]);
  assign or_dcpl_406 = (fsm_output[10]) | (fsm_output[13]);
  assign or_dcpl_407 = or_dcpl_406 | (fsm_output[38]);
  assign or_dcpl_415 = (fsm_output[4]) | (fsm_output[30]);
  assign or_dcpl_417 = (fsm_output[5]) | (fsm_output[29]) | or_dcpl_415;
  assign or_dcpl_418 = (fsm_output[36]) | (fsm_output[11]);
  assign or_dcpl_420 = or_dcpl_418 | or_dcpl_401 | or_dcpl_417;
  assign or_dcpl_421 = (fsm_output[32]) | (fsm_output[8]);
  assign or_dcpl_422 = or_dcpl_421 | or_dcpl_163;
  assign or_dcpl_423 = (fsm_output[13]) | (fsm_output[38]);
  assign or_dcpl_424 = or_dcpl_423 | or_dcpl_99;
  assign or_dcpl_425 = or_dcpl_424 | or_dcpl_422;
  assign and_dcpl_241 = (~ return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva)
      & inverse_lpi_1_dfm_1;
  assign or_dcpl_431 = ~(reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd
      & return_add_generic_AC_RND_CONV_false_9_if_5_return_add_generic_AC_RND_CONV_false_9_if_5_and_tmp);
  assign or_dcpl_438 = or_dcpl_133 | (fsm_output[6]);
  assign or_dcpl_440 = (fsm_output[11]) | (fsm_output[19]);
  assign or_dcpl_444 = (fsm_output[14:13]!=2'b00);
  assign or_dcpl_445 = or_dcpl_444 | (fsm_output[38]);
  assign or_dcpl_447 = (fsm_output[41]) | (fsm_output[39]);
  assign or_dcpl_449 = return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
      | (fsm_output[42]);
  assign or_dcpl_461 = (fsm_output[13]) | (fsm_output[21]);
  assign or_dcpl_462 = or_dcpl_461 | (fsm_output[38]);
  assign or_dcpl_464 = return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
      | (fsm_output[20]);
  assign or_dcpl_465 = (fsm_output[46]) | (fsm_output[44]);
  assign or_dcpl_466 = or_dcpl_465 | (fsm_output[45]);
  assign and_dcpl_257 = ~(and_416_cse | (return_add_generic_AC_RND_CONV_false_4_e_dif_acc_tmp[10]));
  assign and_dcpl_258 = ~(return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_op1_smaller_oelse_and_1_cse
      | (z_out_24[11]));
  assign and_dcpl_259 = ~(return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_and_1_cse
      | (z_out_25[11]));
  assign and_dcpl_260 = ~(return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_7_op1_smaller_oelse_and_cse
      | (z_out_25[11]));
  assign and_dcpl_261 = ~(return_add_generic_AC_RND_CONV_false_9_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_9_op1_smaller_oelse_and_cse
      | (z_out_23[11]));
  assign and_dcpl_262 = ~(return_add_generic_AC_RND_CONV_false_13_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_13_op1_smaller_oelse_and_1_itm
      | (z_out_24[11]));
  assign and_dcpl_263 = ~(return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_and_1_cse
      | (z_out_25[11]));
  assign and_dcpl_264 = ~(return_add_generic_AC_RND_CONV_false_20_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_20_op1_smaller_oelse_and_cse
      | (z_out_26[11]));
  assign and_dcpl_265 = ~(return_add_generic_AC_RND_CONV_false_22_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_22_op1_smaller_oelse_and_cse
      | (z_out_23[11]));
  assign and_dcpl_266 = ~(return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_25_op1_smaller_oelse_and_cse
      | (z_out_25[11]));
  assign or_dcpl_488 = return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
      | (fsm_output[43]);
  assign and_dcpl_267 = ~(return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_8_op1_smaller_oelse_and_cse
      | (z_out_26[11]));
  assign and_dcpl_268 = ~(and_522_cse | (z_out_25[11]));
  assign or_dcpl_493 = (fsm_output[6:5]!=2'b00);
  assign or_dcpl_495 = or_dcpl_493 | (fsm_output[29]) | or_dcpl_415;
  assign or_dcpl_500 = (fsm_output[34]) | (fsm_output[32]);
  assign or_dcpl_501 = or_dcpl_500 | (fsm_output[8]);
  assign or_dcpl_502 = or_dcpl_501 | or_dcpl_163;
  assign or_dcpl_503 = (fsm_output[42]) | (fsm_output[13]);
  assign or_dcpl_511 = or_dcpl_401 | (fsm_output[5]);
  assign or_dcpl_512 = or_dcpl_511 | or_38_cse | (fsm_output[30]);
  assign or_dcpl_513 = or_dcpl_440 | (fsm_output[18]);
  assign or_dcpl_514 = or_dcpl_404 | (fsm_output[36]);
  assign or_dcpl_517 = or_dcpl_163 | (fsm_output[35]);
  assign or_dcpl_518 = or_dcpl_501 | or_dcpl_517;
  assign or_dcpl_519 = or_dcpl_423 | (fsm_output[33]);
  assign and_dcpl_284 = ~((fsm_output[28]) | (fsm_output[3]));
  assign and_dcpl_286 = and_dcpl_211 & and_dcpl_236;
  assign or_dcpl_531 = (fsm_output[45:44]!=2'b00);
  assign or_dcpl_534 = (fsm_output[46]) | (fsm_output[49]);
  assign or_dcpl_542 = or_dcpl_99 | or_dcpl_421;
  assign and_dcpl_326 = ~(return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_12_op1_smaller_oelse_and_cse
      | (z_out_25[11]));
  assign or_dcpl_548 = (fsm_output[10]) | (fsm_output[35]);
  assign or_dcpl_549 = ~(return_add_generic_AC_RND_CONV_false_4_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_17_op1_mu_52_lpi_3_dfm_1 , stage_PE_1_gm_re_d_mux_cse
      , return_add_generic_AC_RND_CONV_false_17_op1_mu_0_lpi_3_dfm_1}) == ({stage_PE_1_gm_im_d_mux_cse
      , stage_PE_1_gm_im_d_mux_2_cse , return_add_generic_AC_RND_CONV_false_17_op2_mu_0_lpi_3_dfm_1})));
  assign or_dcpl_550 = (fsm_output[19:18]!=2'b00);
  assign or_dcpl_551 = or_dcpl_550 | (fsm_output[17]);
  assign or_dcpl_552 = (fsm_output[9]) | (fsm_output[35]);
  assign or_dcpl_553 = or_dcpl_552 | or_dcpl_418;
  assign or_dcpl_556 = or_dcpl_421 | (fsm_output[7]);
  assign or_dcpl_557 = (fsm_output[10]) | (fsm_output[33]);
  assign or_dcpl_558 = or_dcpl_557 | (fsm_output[34]);
  assign or_dcpl_560 = (fsm_output[49]) | (fsm_output[44]);
  assign or_dcpl_561 = or_dcpl_560 | (fsm_output[45]);
  assign or_dcpl_566 = ~(return_add_generic_AC_RND_CONV_false_9_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_22_op1_mu_52_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm
      , return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_9_op2_mu_1_52_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_9_op2_mu_1_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_9_op2_mu_1_0_lpi_3_dfm_1})));
  assign or_dcpl_568 = ~(return_add_generic_AC_RND_CONV_false_23_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm
      , return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm
      , return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1})));
  assign or_dcpl_570 = or_dcpl_557 | or_dcpl_500;
  assign or_dcpl_571 = or_dcpl_570 | or_dcpl_136 | or_dcpl_552;
  assign or_dcpl_573 = (fsm_output[17:16]!=2'b00);
  assign or_dcpl_574 = or_dcpl_550 | or_dcpl_573;
  assign or_dcpl_575 = (fsm_output[21]) | (fsm_output[38]);
  assign or_dcpl_576 = (fsm_output[41]) | (fsm_output[13]);
  assign or_dcpl_579 = (fsm_output[42]) | (fsm_output[20]);
  assign or_dcpl_580 = (fsm_output[15]) | (fsm_output[43]);
  assign or_dcpl_586 = or_dcpl_418 | (fsm_output[31]);
  assign or_dcpl_587 = (fsm_output[35]) | (fsm_output[37]);
  assign or_dcpl_597 = (fsm_output[37:36]!=2'b00);
  assign or_dcpl_607 = (fsm_output[14]) | (fsm_output[38]);
  assign or_dcpl_610 = return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
      | (fsm_output[39]) | or_dcpl_406;
  assign or_dcpl_618 = (fsm_output[12:11]!=2'b00);
  assign or_dcpl_628 = (fsm_output[11]) | (fsm_output[31]);
  assign or_dcpl_631 = or_dcpl_556 | or_dcpl_552;
  assign or_dcpl_660 = (fsm_output[47:46]!=2'b00);
  assign or_dcpl_661 = (fsm_output[23]) | (fsm_output[48]);
  assign or_dcpl_662 = or_dcpl_661 | or_dcpl_660;
  assign or_dcpl_666 = (fsm_output[16]) | (fsm_output[31]);
  assign or_dcpl_682 = (fsm_output[39]) | (fsm_output[13]);
  assign or_dcpl_693 = or_dcpl_493 | (fsm_output[30]);
  assign or_dcpl_694 = (fsm_output[36:35]!=2'b00);
  assign or_dcpl_697 = or_dcpl_136 | (fsm_output[9]);
  assign or_dcpl_704 = (fsm_output[34]) | (fsm_output[8]);
  assign or_dcpl_705 = or_dcpl_575 | (fsm_output[33]);
  assign or_dcpl_707 = (fsm_output[39]) | (fsm_output[10]);
  assign or_dcpl_712 = (fsm_output[11]) | (fsm_output[17]);
  assign or_dcpl_713 = or_dcpl_712 | (fsm_output[16]);
  assign or_dcpl_716 = or_dcpl_99 | (fsm_output[32]);
  assign or_dcpl_719 = or_dcpl_449 | or_dcpl_447 | (fsm_output[10]);
  assign or_dcpl_722 = or_dcpl_401 | return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse;
  assign or_dcpl_736 = (fsm_output[14]) | (fsm_output[21]);
  assign or_dcpl_749 = (fsm_output[20]) | (fsm_output[10]);
  assign or_dcpl_750 = or_dcpl_749 | (fsm_output[21]);
  assign or_dcpl_751 = (fsm_output[45]) | (fsm_output[22]);
  assign or_dcpl_769 = (fsm_output[23]) | (fsm_output[46]);
  assign or_dcpl_776 = (fsm_output[38]) | (fsm_output[33]);
  assign or_dcpl_780 = (fsm_output[34]) | (fsm_output[9]);
  assign or_dcpl_788 = (fsm_output[43:42]!=2'b00);
  assign or_dcpl_789 = or_dcpl_788 | (fsm_output[20]);
  assign or_dcpl_790 = or_dcpl_660 | or_dcpl_531;
  assign or_dcpl_793 = or_dcpl_628 | (fsm_output[6]);
  assign or_dcpl_799 = or_dcpl_406 | (fsm_output[14]);
  assign or_dcpl_803 = (fsm_output[44]) | (fsm_output[40]) | (fsm_output[15]);
  assign or_dcpl_840 = (fsm_output[12]) | (fsm_output[36]) | (fsm_output[11]);
  assign and_dcpl_348 = ~(and_470_cse | (z_out_24[11]));
  assign and_dcpl_349 = ~(and_468_cse | (z_out_24[11]));
  assign or_dcpl_863 = ~((({return_add_generic_AC_RND_CONV_false_op2_mu_52_lpi_3_dfm_1
      , return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx1 , return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1})
      == ({drf_qr_lval_13_smx_0_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1})) & return_add_generic_AC_RND_CONV_false_e1_eq_e2_equal_tmp);
  assign or_dcpl_870 = (fsm_output[22]) | (fsm_output[40]);
  assign or_dcpl_876 = ~(return_add_generic_AC_RND_CONV_false_15_aif_equal_tmp &
      return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp);
  assign or_dcpl_882 = or_dcpl_803 | or_dcpl_789;
  assign or_dcpl_906 = or_dcpl_736 | (fsm_output[38]);
  assign or_dcpl_911 = ~((({drf_qr_lval_13_smx_0_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_op2_mu_52_lpi_3_dfm_1
      , return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx1 , return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1}))
      & return_add_generic_AC_RND_CONV_false_1_e1_eq_e2_equal_tmp);
  assign or_dcpl_912 = ~(return_add_generic_AC_RND_CONV_false_10_e1_eq_e2_equal_tmp
      & (({drf_qr_lval_13_smx_0_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_10_op2_mu_1_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_10_op2_mu_1_50_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1})));
  assign or_dcpl_913 = ~((({drf_qr_lval_13_smx_0_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_13_op1_mu_52_lpi_3_dfm_1
      , return_extract_32_mux_4_cse , return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1}))
      & return_add_generic_AC_RND_CONV_false_14_e1_eq_e2_equal_tmp);
  assign or_dcpl_914 = ~(return_add_generic_AC_RND_CONV_false_22_e1_eq_e2_equal_tmp
      & (({return_add_generic_AC_RND_CONV_false_22_op1_mu_52_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm
      , return_add_generic_AC_RND_CONV_false_9_op1_mu_0_lpi_3_dfm_1}) == ({return_add_generic_AC_RND_CONV_false_22_op2_mu_1_52_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_22_op2_mu_1_51_lpi_3_dfm_mx0 , return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0
      , return_add_generic_AC_RND_CONV_false_22_op2_mu_1_0_lpi_3_dfm_1})));
  assign or_dcpl_919 = or_dcpl_719 | or_dcpl_445 | or_dcpl_99;
  assign or_dcpl_928 = or_dcpl_870 | (fsm_output[15]);
  assign or_dcpl_929 = or_dcpl_661 | (fsm_output[47]);
  assign or_dcpl_937 = or_dcpl_929 | or_dcpl_106;
  assign or_dcpl_940 = (fsm_output[36]) | (fsm_output[19]);
  assign or_dcpl_949 = or_dcpl_661 | (fsm_output[50]);
  assign or_dcpl_953 = or_dcpl_552 | (fsm_output[36]);
  assign or_dcpl_961 = (fsm_output[49]) | (fsm_output[22]);
  assign or_dcpl_976 = or_dcpl_531 | (fsm_output[22]);
  assign or_dcpl_985 = (fsm_output[43]) | (fsm_output[20]);
  assign or_dcpl_999 = (fsm_output[22]) | (fsm_output[25]) | (fsm_output[24]);
  assign or_dcpl_1001 = or_dcpl_929 | or_dcpl_466;
  assign or_dcpl_1015 = (fsm_output[32]) | (fsm_output[9]);
  assign or_dcpl_1069 = operator_11_true_return_26_sva | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva;
  assign and_dcpl_385 = (~ return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva)
      & inverse_lpi_1_dfm_1;
  assign and_dcpl_399 = and_dcpl_28 & (~ return_add_generic_AC_RND_CONV_false_10_op1_nan_sva);
  assign and_dcpl_408 = ~(operator_11_true_return_15_sva | operator_11_true_return_1_sva
      | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva);
  assign and_dcpl_413 = and_dcpl_28 & (~(operator_11_true_return_17_sva | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva));
  assign or_tmp_61 = operator_16_false_operator_16_false_nor_cse_sva & (fsm_output[54]);
  assign and_571_cse = and_dcpl_146 & (fsm_output[54]);
  assign and_592_cse = and_dcpl_140 & or_dcpl_11;
  assign or_tmp_82 = inverse_lpi_1_dfm_1 & (fsm_output[3]);
  assign or_tmp_83 = (~ inverse_lpi_1_dfm_1) & (fsm_output[3]);
  assign and_666_cse = and_dcpl_140 & (fsm_output[53]);
  assign or_tmp_112 = inverse_lpi_1_dfm_1 & (fsm_output[28]);
  assign or_tmp_113 = (~ inverse_lpi_1_dfm_1) & (fsm_output[28]);
  assign or_tmp_208 = (~ inverse_lpi_1_dfm_1) & (fsm_output[2]);
  assign or_tmp_234 = (fsm_output[46]) | (fsm_output[21]);
  assign or_tmp_261 = (fsm_output[31:30]!=2'b00);
  assign and_1013_cse = (fsm_output[44]) | (fsm_output[13]) | (fsm_output[38]) |
      or_dcpl_404 | or_dcpl_418 | or_dcpl_133;
  assign or_tmp_348 = return_add_generic_AC_RND_CONV_false_9_op1_smaller_return_add_generic_AC_RND_CONV_false_9_op1_smaller_or_cse
      & (fsm_output[16]);
  assign and_1163_cse = return_add_generic_AC_RND_CONV_false_25_op1_smaller_return_add_generic_AC_RND_CONV_false_25_op1_smaller_or_cse
      & (fsm_output[43]);
  assign or_tmp_403 = or_dcpl_423 | or_dcpl_597;
  assign or_tmp_440 = (fsm_output[6]) | (fsm_output[4]);
  assign and_1583_cse = return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse
      & (fsm_output[5]);
  assign and_1584_cse = return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse
      & (fsm_output[30]);
  assign or_tmp_561 = and_1583_cse | and_1584_cse;
  assign or_tmp_564 = inverse_lpi_1_dfm_1 & (fsm_output[10]);
  assign and_1598_cse = return_add_generic_AC_RND_CONV_false_7_op1_smaller_return_add_generic_AC_RND_CONV_false_7_op1_smaller_or_cse
      & (fsm_output[14]);
  assign or_tmp_570 = inverse_lpi_1_dfm_1 & (fsm_output[35]);
  assign and_1608_cse = return_add_generic_AC_RND_CONV_false_20_op1_smaller_return_add_generic_AC_RND_CONV_false_20_op1_smaller_or_cse
      & (fsm_output[39]);
  assign or_tmp_771 = (fsm_output[22]) | (fsm_output[16]) | (fsm_output[31]);
  assign or_tmp_823 = return_add_generic_AC_RND_CONV_false_22_op1_smaller_return_add_generic_AC_RND_CONV_false_22_op1_smaller_or_cse
      & (fsm_output[41]);
  assign or_tmp_852 = (fsm_output[44]) | (fsm_output[18]) | (fsm_output[17]);
  assign or_tmp_857 = or_dcpl_488 | (fsm_output[42]) | (fsm_output[19]);
  assign and_2281_cse = return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse
      & (fsm_output[18]);
  assign out1_rsci_idat_63_0_mx0c1 = and_dcpl_138 & and_dcpl_129 & (operator_16_false_io_read_mode1_rsc_cse_sva[2:0]==3'b001)
      & (~ operator_16_false_operator_16_false_nor_cse_sva) & (fsm_output[54]);
  assign out1_rsci_idat_63_0_mx0c2 = and_dcpl_140 & (fsm_output[54]);
  assign out1_rsci_idat_79_64_mx0c1 = and_dcpl_138 & and_dcpl_129 & (operator_16_false_io_read_mode1_rsc_cse_sva[2:1]==2'b01)
      & (~((operator_16_false_io_read_mode1_rsc_cse_sva[0]) | operator_16_false_operator_16_false_nor_cse_sva))
      & (fsm_output[54]);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx6c1 = ~(return_add_generic_AC_RND_CONV_false_13_return_add_generic_AC_RND_CONV_false_13_or_1_tmp
      | inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx6c2 = return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse
      & inverse_lpi_1_dfm_1;
  assign stage_PE_1_tmp_im_d_1_sva_1_mx0c3 = or_dcpl_790 | or_dcpl_789 | (fsm_output[41])
      | (fsm_output[37]) | (fsm_output[12]) | or_dcpl_550 | (fsm_output[16]);
  assign stage_PE_1_tmp_re_d_1_sva_1_mx0c0 = or_dcpl_976 | or_dcpl_985 | (fsm_output[21])
      | or_dcpl_551 | or_dcpl_401;
  assign stage_PE_1_tmp_re_d_1_sva_1_mx0c4 = or_dcpl_548 | or_dcpl_418;
  assign not_tmp_302 = return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm
      ^ stage_PE_tmp_im_d_1_lpi_3_dfm_63_mx0;
  assign BUTTERFLY_1_i_mux1h_1_nl = MUX1HOT_s_1_7_2((BUTTERFLY_1_i_9_0_sva[9]), (~
      (BUTTERFLY_1_i_9_0_sva[9])), (BUTTERFLY_1_fry_9_0_sva[9]), (~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm),
      (z_out_2[9]), (~ (z_out_2[9])), (~ (BUTTERFLY_1_fry_9_0_sva[9])), {or_1231_ssc
      , or_1232_ssc , or_1233_ssc , or_1234_ssc , or_tmp_112 , or_tmp_113 , and_720_ssc});
  assign or_2472_nl = or_1231_ssc | or_1232_ssc;
  assign or_2473_nl = and_720_ssc | or_1233_ssc;
  assign mux1h_6_nl = MUX1HOT_v_9_4_2((BUTTERFLY_1_i_9_0_sva[8:0]), BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2,
      (BUTTERFLY_1_fry_9_0_sva[8:0]), (z_out_2[8:0]), {or_2472_nl , or_1234_ssc ,
      or_2473_nl , BUTTERFLY_1_i_or_cse});
  assign in_f_d_rsci_adr_d = {BUTTERFLY_1_i_mux1h_1_nl , mux1h_6_nl};
  assign nor_160_m1c = ~(or_tmp | or_tmp_916 | or_tmp_917);
  assign nor_161_m1c = ~(BUTTERFLY_if_1_if_or_1_cse | or_tmp_919);
  assign BUTTERFLY_if_1_if_and_9_cse = return_add_generic_AC_RND_CONV_false_10_or_1_svs_1
      & (fsm_output[22]);
  assign BUTTERFLY_if_1_if_and_5_cse = return_add_generic_AC_RND_CONV_false_or_1_svs_1
      & (fsm_output[6]);
  assign BUTTERFLY_if_1_if_and_11_cse = return_add_generic_AC_RND_CONV_false_12_or_1_svs_1
      & (fsm_output[26]);
  assign BUTTERFLY_if_1_if_and_8_cse = return_add_generic_AC_RND_CONV_false_9_or_1_svs_1
      & (fsm_output[20]);
  assign BUTTERFLY_if_1_if_and_10_cse = return_add_generic_AC_RND_CONV_false_11_or_1_svs_1
      & (fsm_output[24]);
  assign BUTTERFLY_if_1_if_and_6_cse = return_add_generic_AC_RND_CONV_false_1_or_1_svs_1
      & (fsm_output[8]);
  assign BUTTERFLY_if_1_if_or_1_cse = ((~ return_add_generic_AC_RND_CONV_false_or_1_svs_1)
      & (fsm_output[6])) | ((~ return_add_generic_AC_RND_CONV_false_9_or_1_svs_1)
      & (fsm_output[20])) | ((~ return_add_generic_AC_RND_CONV_false_10_or_1_svs_1)
      & (fsm_output[22])) | ((~ return_add_generic_AC_RND_CONV_false_11_or_1_svs_1)
      & (fsm_output[24])) | ((~ return_add_generic_AC_RND_CONV_false_12_or_1_svs_1)
      & (fsm_output[26]));
  assign BUTTERFLY_if_1_if_or_nl = (fsm_output[6]) | (fsm_output[8]) | (fsm_output[22]);
  assign BUTTERFLY_if_1_if_mux1h_nl = MUX1HOT_s_1_6_2(operator_11_true_return_26_sva,
      return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva,
      return_add_generic_AC_RND_CONV_false_17_mux_6_itm, return_add_generic_AC_RND_CONV_false_11_mux_itm,
      return_add_generic_AC_RND_CONV_false_12_mux_itm, {BUTTERFLY_if_1_if_or_nl ,
      (fsm_output[16]) , (fsm_output[18]) , (fsm_output[20]) , (fsm_output[24]) ,
      (fsm_output[26])});
  assign and_2423_nl = (fsm_output[6]) & nor_160_m1c;
  assign and_2424_nl = (fsm_output[8]) & nor_160_m1c;
  assign and_2425_nl = (fsm_output[16]) & nor_160_m1c;
  assign and_2426_nl = (fsm_output[18]) & nor_160_m1c;
  assign or_2461_nl = ((fsm_output[20]) & nor_160_m1c) | ((fsm_output[22]) & nor_160_m1c)
      | ((fsm_output[24]) & nor_160_m1c) | ((fsm_output[26]) & nor_160_m1c);
  assign mux1h_nl = MUX1HOT_v_10_6_2(return_add_generic_AC_RND_CONV_false_e_r_return_add_generic_AC_RND_CONV_false_e_r_or_cse,
      return_add_generic_AC_RND_CONV_false_1_e_r_return_add_generic_AC_RND_CONV_false_1_e_r_or_cse,
      return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1,
      (return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_5_cse[9:0]),
      return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_11,
      {and_2423_nl , and_2424_nl , and_2425_nl , and_2426_nl , or_2461_nl , or_tmp_916});
  assign not_760_nl = ~ or_tmp_917;
  assign and_2431_nl = MUX_v_10_2_2(10'b0000000000, mux1h_nl, not_760_nl);
  assign or_2035_nl = MUX_v_10_2_2(and_2431_nl, 10'b1111111111, or_tmp);
  assign or_245_nl = return_add_generic_AC_RND_CONV_false_r_inf_lpi_3_dfm_2 | operator_11_true_return_1_sva
      | and_dcpl_166 | operator_11_true_return_24_sva;
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs, or_245_nl);
  assign return_add_generic_AC_RND_CONV_false_e_r_return_add_generic_AC_RND_CONV_false_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_6_mux_35 & (~ return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_nl))
      | return_add_generic_AC_RND_CONV_false_exception_sva_1;
  assign or_257_nl = return_add_generic_AC_RND_CONV_false_1_r_inf_lpi_3_dfm_2 | operator_11_true_return_1_sva
      | and_dcpl_168 | operator_11_true_return_24_sva;
  assign return_add_generic_AC_RND_CONV_false_14_e_r_qelse_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs, or_257_nl);
  assign return_add_generic_AC_RND_CONV_false_1_e_r_return_add_generic_AC_RND_CONV_false_1_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_32 & (~ return_add_generic_AC_RND_CONV_false_14_e_r_qelse_mux_nl))
      | return_add_generic_AC_RND_CONV_false_1_exception_sva_1;
  assign or_375_nl = return_add_generic_AC_RND_CONV_false_9_r_inf_lpi_3_dfm_2 | return_add_generic_AC_RND_CONV_false_23_op1_inf_sva
      | return_add_generic_AC_RND_CONV_false_23_op1_nan_sva | operator_11_true_return_1_sva
      | and_dcpl_166;
  assign return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs, or_375_nl);
  assign return_add_generic_AC_RND_CONV_false_9_e_r_return_add_generic_AC_RND_CONV_false_9_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_6_mux_35 & (~ return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_nl))
      | return_add_generic_AC_RND_CONV_false_9_exception_sva_1;
  assign or_386_nl = return_add_generic_AC_RND_CONV_false_10_r_inf_lpi_3_dfm_2 |
      operator_11_true_return_15_sva | or_dcpl_275 | and_dcpl_166;
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_21_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs, or_386_nl);
  assign return_add_generic_AC_RND_CONV_false_10_e_r_return_add_generic_AC_RND_CONV_false_10_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_6_mux_35 & (~ return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_21_nl))
      | return_add_generic_AC_RND_CONV_false_10_exception_sva_1;
  assign or_397_nl = return_add_generic_AC_RND_CONV_false_11_r_inf_lpi_3_dfm_2 |
      or_dcpl_201 | or_dcpl_199 | and_dcpl_166;
  assign return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_5_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs, or_397_nl);
  assign return_add_generic_AC_RND_CONV_false_11_e_r_return_add_generic_AC_RND_CONV_false_11_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_6_mux_35 & (~ return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_5_nl))
      | return_add_generic_AC_RND_CONV_false_11_exception_sva_1;
  assign or_407_nl = return_add_generic_AC_RND_CONV_false_12_r_inf_lpi_3_dfm_2 |
      or_dcpl_214 | or_dcpl_275 | and_dcpl_166;
  assign return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_3_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs, or_407_nl);
  assign return_add_generic_AC_RND_CONV_false_12_e_r_return_add_generic_AC_RND_CONV_false_12_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_6_mux_35 & (~ return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_3_nl))
      | return_add_generic_AC_RND_CONV_false_12_exception_sva_1;
  assign BUTTERFLY_if_1_if_mux1h_2_nl = MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_e_r_return_add_generic_AC_RND_CONV_false_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_1_e_r_return_add_generic_AC_RND_CONV_false_1_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_9_e_r_return_add_generic_AC_RND_CONV_false_9_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_10_e_r_return_add_generic_AC_RND_CONV_false_10_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_11_e_r_return_add_generic_AC_RND_CONV_false_11_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_12_e_r_return_add_generic_AC_RND_CONV_false_12_e_r_or_1_nl,
      {(fsm_output[6]) , (fsm_output[8]) , (fsm_output[16]) , (fsm_output[18]) ,
      (fsm_output[20]) , (fsm_output[22]) , (fsm_output[24]) , (fsm_output[26])});
  assign return_add_generic_AC_RND_CONV_false_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_9_op1_nan_sva_1
      | return_add_generic_AC_RND_CONV_false_1_op1_nan_sva_mx3w0 | (return_add_generic_AC_RND_CONV_false_9_op1_inf_sva_1
      & return_extract_2_and_1_tmp & return_add_generic_AC_RND_CONV_false_12_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_9_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_23_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_9_op2_nan_sva_mx7w0 | (return_add_generic_AC_RND_CONV_false_23_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_9_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_14_op2_nan_sva);
  assign return_add_generic_AC_RND_CONV_false_10_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_11_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_23_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva | return_add_generic_AC_RND_CONV_false_10_unequal_tmp;
  assign return_add_generic_AC_RND_CONV_false_12_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | operator_11_true_return_1_sva;
  assign BUTTERFLY_if_1_if_or_2_nl = BUTTERFLY_if_1_if_and_5_cse | BUTTERFLY_if_1_if_and_6_cse;
  assign BUTTERFLY_if_1_if_and_7_nl = (~ return_add_generic_AC_RND_CONV_false_1_or_1_svs_1)
      & (fsm_output[8]);
  assign BUTTERFLY_if_1_if_mux1h_3_nl = MUX1HOT_s_1_9_2(return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_r_nan_or_nl, (return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_and_5_cse[51]),
      return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_8_m_r_51_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_9_r_nan_or_nl, return_add_generic_AC_RND_CONV_false_10_r_nan_or_nl,
      return_add_generic_AC_RND_CONV_false_11_r_nan_or_nl, return_add_generic_AC_RND_CONV_false_12_r_nan_or_nl,
      {BUTTERFLY_if_1_if_or_1_cse , BUTTERFLY_if_1_if_or_2_nl , BUTTERFLY_if_1_if_and_7_nl
      , (fsm_output[16]) , (fsm_output[18]) , BUTTERFLY_if_1_if_and_8_cse , BUTTERFLY_if_1_if_and_9_cse
      , BUTTERFLY_if_1_if_and_10_cse , BUTTERFLY_if_1_if_and_11_cse});
  assign and_2433_nl = (fsm_output[8]) & nor_161_m1c;
  assign and_2434_nl = (fsm_output[16]) & nor_161_m1c;
  assign and_2435_nl = (fsm_output[18]) & nor_161_m1c;
  assign mux1h_1_nl = MUX1HOT_v_51_4_2((return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_and_5_cse[50:0]),
      return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm,
      {and_2433_nl , and_2434_nl , and_2435_nl , BUTTERFLY_if_1_if_or_1_cse});
  assign and_2432_nl = ((fsm_output[6]) | (fsm_output[20]) | (fsm_output[22]) | (fsm_output[24])
      | (fsm_output[26])) & nor_161_m1c;
  assign nor_183_nl = ~(MUX_v_51_2_2(mux1h_1_nl, 51'b111111111111111111111111111111111111111111111111111,
      and_2432_nl));
  assign nor_182_nl = ~(MUX_v_51_2_2(nor_183_nl, 51'b111111111111111111111111111111111111111111111111111,
      or_tmp_919));
  assign in_f_d_rsci_d_d = {BUTTERFLY_if_1_if_mux1h_nl , or_2035_nl , BUTTERFLY_if_1_if_mux1h_2_nl
      , BUTTERFLY_if_1_if_mux1h_3_nl , nor_182_nl};
  assign in_f_d_rsci_we_d_pff = (and_dcpl_1 & (or_dcpl_166 | (fsm_output[24]) | (fsm_output[20])))
      | (stage_PE_1_and_1_tmp & ((fsm_output[8]) | (fsm_output[18]) | or_dcpl_132));
  assign in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = (mode_lpi_1_dfm & ((fsm_output[28])
      | (fsm_output[31]) | or_dcpl_118)) | and_666_cse;
  assign BUTTERFLY_1_i_or_cse = or_tmp_112 | or_tmp_113;
  assign or_1217_nl = (fsm_output[8]) | (fsm_output[5]) | (fsm_output[29]);
  assign or_1218_nl = or_dcpl_11 | or_dcpl_163;
  assign in_u_rsci_adr_d = MUX1HOT_v_10_3_2(BUTTERFLY_1_i_9_0_sva, BUTTERFLY_1_fry_9_0_sva,
      z_out_2, {or_1217_nl , or_1218_nl , BUTTERFLY_1_i_or_cse});
  assign mux1h_7_nl = MUX1HOT_v_2_4_2((z_out_45[15:14]), BUTTERFLY_1_else_3_else_acc_4_itm_15_14,
      (signext_2_1(stage_monty_mul_acc_2_psp_sva_1[14])), (z_out_38[15:14]), {(fsm_output[7])
      , (fsm_output[9]) , (fsm_output[54]) , or_dcpl_1189});
  assign mux1h_8_nl = MUX1HOT_v_3_4_2((z_out_45[13:11]), BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_0,
      (stage_monty_mul_acc_2_psp_sva_1[13:11]), (z_out_38[13:11]), {(fsm_output[7])
      , (fsm_output[9]) , (fsm_output[54]) , or_dcpl_1189});
  assign mux1h_12_nl = MUX1HOT_s_1_4_2((z_out_45[10]), BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1,
      (stage_monty_mul_acc_2_psp_sva_1[10]), (z_out_38[10]), {(fsm_output[7]) , (fsm_output[9])
      , (fsm_output[54]) , or_dcpl_1189});
  assign mux1h_13_nl = MUX1HOT_v_5_4_2((z_out_45[9:5]), reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd,
      (stage_monty_mul_acc_2_psp_sva_1[9:5]), (z_out_38[9:5]), {(fsm_output[7]) ,
      (fsm_output[9]) , (fsm_output[54]) , or_dcpl_1189});
  assign mux1h_14_nl = MUX1HOT_v_5_4_2((z_out_45[4:0]), reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1,
      (stage_monty_mul_acc_2_psp_sva_1[4:0]), (z_out_38[4:0]), {(fsm_output[7]) ,
      (fsm_output[9]) , (fsm_output[54]) , or_dcpl_1189});
  assign in_u_rsci_d_d = {mux1h_7_nl , mux1h_8_nl , mux1h_12_nl , mux1h_13_nl , mux1h_14_nl};
  assign in_u_rsci_we_d_pff = (stage_PE_1_and_cse & or_219_cse) | (nor_3_cse & or_dcpl_159)
      | and_571_cse;
  assign in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = (~(mode_lpi_1_dfm | (~((fsm_output[29:28]!=2'b00)))))
      | and_666_cse;
  assign BUTTERFLY_if_1_mux1h_2_nl = MUX1HOT_s_1_7_2((z_out_2[9]), (~ (z_out_2[9])),
      (BUTTERFLY_1_i_9_0_sva[9]), (~ (BUTTERFLY_1_i_9_0_sva[9])), (~ (BUTTERFLY_1_fry_9_0_sva[9])),
      (BUTTERFLY_1_fry_9_0_sva[9]), (~ BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm),
      {or_tmp_82 , or_tmp_83 , or_1205_ssc , or_1206_ssc , and_654_ssc , or_1208_ssc
      , or_1209_ssc});
  assign or_2474_nl = or_1205_ssc | or_1206_ssc;
  assign or_2475_nl = or_1208_ssc | and_654_ssc;
  assign mux1h_9_nl = MUX1HOT_v_9_4_2((BUTTERFLY_1_i_9_0_sva[8:0]), BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2,
      (BUTTERFLY_1_fry_9_0_sva[8:0]), (z_out_2[8:0]), {or_2474_nl , or_1209_ssc ,
      or_2475_nl , BUTTERFLY_else_1_or_cse});
  assign out_f_d_rsci_adr_d = {BUTTERFLY_if_1_mux1h_2_nl , mux1h_9_nl};
  assign nor_162_m1c = ~(or_tmp_920 | or_tmp_921 | or_tmp_922);
  assign nor_163_m1c = ~(BUTTERFLY_if_1_or_1_cse | or_tmp_924);
  assign BUTTERFLY_if_1_and_7_cse = return_add_generic_AC_RND_CONV_false_13_or_1_svs_1
      & (fsm_output[31]);
  assign BUTTERFLY_if_1_and_11_cse = return_add_generic_AC_RND_CONV_false_23_or_1_svs_1
      & (fsm_output[47]);
  assign BUTTERFLY_if_1_and_13_cse = return_add_generic_AC_RND_CONV_false_25_or_1_svs_1
      & (fsm_output[51]);
  assign BUTTERFLY_if_1_and_10_cse = return_add_generic_AC_RND_CONV_false_22_or_1_svs_1
      & (fsm_output[45]);
  assign BUTTERFLY_if_1_and_12_cse = return_add_generic_AC_RND_CONV_false_24_or_1_svs_1
      & (fsm_output[49]);
  assign BUTTERFLY_if_1_and_8_cse = return_add_generic_AC_RND_CONV_false_14_or_1_svs_1
      & (fsm_output[33]);
  assign BUTTERFLY_if_1_or_1_cse = ((~ return_add_generic_AC_RND_CONV_false_13_or_1_svs_1)
      & (fsm_output[31])) | ((~ return_add_generic_AC_RND_CONV_false_22_or_1_svs_1)
      & (fsm_output[45])) | ((~ return_add_generic_AC_RND_CONV_false_23_or_1_svs_1)
      & (fsm_output[47])) | ((~ return_add_generic_AC_RND_CONV_false_24_or_1_svs_1)
      & (fsm_output[49])) | ((~ return_add_generic_AC_RND_CONV_false_25_or_1_svs_1)
      & (fsm_output[51]));
  assign BUTTERFLY_if_1_or_nl = (fsm_output[31]) | (fsm_output[33]) | (fsm_output[45]);
  assign BUTTERFLY_if_1_mux1h_1_nl = MUX1HOT_s_1_6_2(operator_11_true_return_26_sva,
      return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva,
      return_add_generic_AC_RND_CONV_false_11_mux_itm, return_add_generic_AC_RND_CONV_false_12_mux_itm,
      return_add_generic_AC_RND_CONV_false_17_mux_6_itm, {BUTTERFLY_if_1_or_nl ,
      (fsm_output[41]) , (fsm_output[43]) , (fsm_output[47]) , (fsm_output[49]) ,
      (fsm_output[51])});
  assign and_2441_nl = (fsm_output[31]) & nor_162_m1c;
  assign and_2442_nl = (fsm_output[33]) & nor_162_m1c;
  assign and_2443_nl = (fsm_output[41]) & nor_162_m1c;
  assign and_2444_nl = (fsm_output[43]) & nor_162_m1c;
  assign or_2460_nl = ((fsm_output[45]) & nor_162_m1c) | ((fsm_output[47]) & nor_162_m1c)
      | ((fsm_output[49]) & nor_162_m1c) | ((fsm_output[51]) & nor_162_m1c);
  assign mux1h_2_nl = MUX1HOT_v_10_6_2(return_add_generic_AC_RND_CONV_false_e_r_return_add_generic_AC_RND_CONV_false_e_r_or_cse,
      return_add_generic_AC_RND_CONV_false_1_e_r_return_add_generic_AC_RND_CONV_false_1_e_r_or_cse,
      return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1,
      (return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_5_cse[9:0]),
      return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_11,
      {and_2441_nl , and_2442_nl , and_2443_nl , and_2444_nl , or_2460_nl , or_tmp_921});
  assign not_763_nl = ~ or_tmp_922;
  assign and_2449_nl = MUX_v_10_2_2(10'b0000000000, mux1h_2_nl, not_763_nl);
  assign or_2036_nl = MUX_v_10_2_2(and_2449_nl, 10'b1111111111, or_tmp_920);
  assign or_320_nl = return_add_generic_AC_RND_CONV_false_13_r_inf_lpi_3_dfm_2 |
      operator_11_true_return_15_sva | and_dcpl_166 | operator_11_true_return_1_sva;
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_11_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs, or_320_nl);
  assign return_add_generic_AC_RND_CONV_false_13_e_r_return_add_generic_AC_RND_CONV_false_13_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_6_mux_35 & (~ return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_11_nl))
      | return_add_generic_AC_RND_CONV_false_13_exception_sva_1;
  assign or_332_nl = return_add_generic_AC_RND_CONV_false_14_r_inf_lpi_3_dfm_2 |
      operator_11_true_return_15_sva | and_dcpl_168 | operator_11_true_return_1_sva;
  assign return_add_generic_AC_RND_CONV_false_14_e_r_qelse_mux_3_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs, or_332_nl);
  assign return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_1_mux_32 & (~ return_add_generic_AC_RND_CONV_false_14_e_r_qelse_mux_3_nl))
      | return_add_generic_AC_RND_CONV_false_14_exception_sva_1;
  assign or_417_nl = return_add_generic_AC_RND_CONV_false_22_r_inf_lpi_3_dfm_2 |
      operator_11_true_return_1_sva | or_dcpl_225 | and_dcpl_166;
  assign return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_7_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs, or_417_nl);
  assign return_add_generic_AC_RND_CONV_false_22_e_r_return_add_generic_AC_RND_CONV_false_22_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_6_mux_35 & (~ return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_7_nl))
      | return_add_generic_AC_RND_CONV_false_22_exception_sva_1;
  assign or_429_nl = return_add_generic_AC_RND_CONV_false_23_r_inf_lpi_3_dfm_2 |
      return_add_generic_AC_RND_CONV_false_23_op1_inf_sva | return_add_generic_AC_RND_CONV_false_23_op1_nan_sva
      | operator_11_true_return_15_sva | and_dcpl_166;
  assign return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_23_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs, or_429_nl);
  assign return_add_generic_AC_RND_CONV_false_23_e_r_return_add_generic_AC_RND_CONV_false_23_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_6_mux_35 & (~ return_add_generic_AC_RND_CONV_false_6_e_r_qelse_mux_23_nl))
      | return_add_generic_AC_RND_CONV_false_23_exception_sva_1;
  assign or_439_nl = return_add_generic_AC_RND_CONV_false_24_r_inf_lpi_3_dfm_2 |
      or_dcpl_214 | or_dcpl_225 | and_dcpl_166;
  assign return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_5_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs, or_439_nl);
  assign return_add_generic_AC_RND_CONV_false_24_e_r_return_add_generic_AC_RND_CONV_false_24_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_6_mux_35 & (~ return_add_generic_AC_RND_CONV_false_12_e_r_qelse_mux_5_nl))
      | return_add_generic_AC_RND_CONV_false_24_exception_sva_1;
  assign or_449_nl = return_add_generic_AC_RND_CONV_false_25_r_inf_lpi_3_dfm_2 |
      or_dcpl_201 | or_dcpl_199 | and_dcpl_166;
  assign return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_9_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0,
      return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs, or_449_nl);
  assign return_add_generic_AC_RND_CONV_false_25_e_r_return_add_generic_AC_RND_CONV_false_25_e_r_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_6_mux_35 & (~ return_add_generic_AC_RND_CONV_false_11_e_r_qelse_mux_9_nl))
      | return_add_generic_AC_RND_CONV_false_25_exception_sva_1;
  assign BUTTERFLY_if_1_mux1h_6_nl = MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_13_e_r_return_add_generic_AC_RND_CONV_false_13_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_14_e_r_return_add_generic_AC_RND_CONV_false_14_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_22_e_r_return_add_generic_AC_RND_CONV_false_22_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_23_e_r_return_add_generic_AC_RND_CONV_false_23_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_24_e_r_return_add_generic_AC_RND_CONV_false_24_e_r_or_1_nl,
      return_add_generic_AC_RND_CONV_false_25_e_r_return_add_generic_AC_RND_CONV_false_25_e_r_or_1_nl,
      {(fsm_output[31]) , (fsm_output[33]) , (fsm_output[41]) , (fsm_output[43])
      , (fsm_output[45]) , (fsm_output[47]) , (fsm_output[49]) , (fsm_output[51])});
  assign return_add_generic_AC_RND_CONV_false_13_r_nan_or_1_nl = return_add_generic_AC_RND_CONV_false_9_op2_nan_sva_mx7w0
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_9_op2_inf_sva_1
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_12_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_22_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_22_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_22_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_11_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_23_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_23_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1 | (return_add_generic_AC_RND_CONV_false_23_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1 & return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_24_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | return_add_generic_AC_RND_CONV_false_10_unequal_tmp;
  assign return_add_generic_AC_RND_CONV_false_25_r_nan_or_nl = return_add_generic_AC_RND_CONV_false_23_op1_nan_sva
      | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva | operator_11_true_return_1_sva;
  assign BUTTERFLY_if_1_or_2_nl = BUTTERFLY_if_1_and_7_cse | BUTTERFLY_if_1_and_8_cse;
  assign BUTTERFLY_if_1_and_9_nl = (~ return_add_generic_AC_RND_CONV_false_14_or_1_svs_1)
      & (fsm_output[33]);
  assign BUTTERFLY_if_1_mux1h_7_nl = MUX1HOT_s_1_9_2(return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_13_r_nan_or_1_nl, (return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_and_5_cse[51]),
      return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_21_m_r_51_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_22_r_nan_or_nl, return_add_generic_AC_RND_CONV_false_23_r_nan_or_nl,
      return_add_generic_AC_RND_CONV_false_24_r_nan_or_nl, return_add_generic_AC_RND_CONV_false_25_r_nan_or_nl,
      {BUTTERFLY_if_1_or_1_cse , BUTTERFLY_if_1_or_2_nl , BUTTERFLY_if_1_and_9_nl
      , (fsm_output[41]) , (fsm_output[43]) , BUTTERFLY_if_1_and_10_cse , BUTTERFLY_if_1_and_11_cse
      , BUTTERFLY_if_1_and_12_cse , BUTTERFLY_if_1_and_13_cse});
  assign and_2451_nl = (fsm_output[33]) & nor_163_m1c;
  assign and_2452_nl = (fsm_output[41]) & nor_163_m1c;
  assign and_2453_nl = (fsm_output[43]) & nor_163_m1c;
  assign mux1h_3_nl = MUX1HOT_v_51_4_2((return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_and_5_cse[50:0]),
      return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm,
      {and_2451_nl , and_2452_nl , and_2453_nl , BUTTERFLY_if_1_or_1_cse});
  assign and_2450_nl = ((fsm_output[31]) | (fsm_output[45]) | (fsm_output[47]) |
      (fsm_output[49]) | (fsm_output[51])) & nor_163_m1c;
  assign nor_187_nl = ~(MUX_v_51_2_2(mux1h_3_nl, 51'b111111111111111111111111111111111111111111111111111,
      and_2450_nl));
  assign nor_186_nl = ~(MUX_v_51_2_2(nor_187_nl, 51'b111111111111111111111111111111111111111111111111111,
      or_tmp_924));
  assign out_f_d_rsci_d_d = {BUTTERFLY_if_1_mux1h_1_nl , or_2036_nl , BUTTERFLY_if_1_mux1h_6_nl
      , BUTTERFLY_if_1_mux1h_7_nl , nor_186_nl};
  assign out_f_d_rsci_we_d_pff = (stage_PE_1_and_1_tmp & ((fsm_output[43]) | (fsm_output[41])
      | (fsm_output[33]) | (fsm_output[31]))) | (and_dcpl_1 & (or_dcpl_148 | or_dcpl_105));
  assign out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = (mode_lpi_1_dfm & ((fsm_output[3])
      | (fsm_output[6]) | or_dcpl_95)) | (or_dcpl_115 & (fsm_output[53]));
  assign BUTTERFLY_else_1_or_cse = or_tmp_82 | or_tmp_83;
  assign or_1191_nl = (fsm_output[33]) | (fsm_output[4]) | (fsm_output[30]);
  assign or_1192_nl = (fsm_output[53]) | (fsm_output[34]) | (fsm_output[32]);
  assign out_u_rsci_adr_d = MUX1HOT_v_10_3_2(z_out_2, BUTTERFLY_1_i_9_0_sva, BUTTERFLY_1_fry_9_0_sva,
      {BUTTERFLY_else_1_or_cse , or_1191_nl , or_1192_nl});
  assign nor_204_cse = ~((fsm_output[34]) | or_dcpl_1191);
  assign mux1h_10_nl = MUX1HOT_v_2_3_2((z_out_45[15:14]), BUTTERFLY_1_else_3_else_acc_4_itm_15_14,
      (z_out_38[15:14]), {nor_204_cse , (fsm_output[34]) , or_dcpl_1191});
  assign mux1h_11_nl = MUX1HOT_v_3_3_2((z_out_45[13:11]), BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_0,
      (z_out_38[13:11]), {nor_204_cse , (fsm_output[34]) , or_dcpl_1191});
  assign mux1h_15_nl = MUX1HOT_s_1_3_2((z_out_45[10]), BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1,
      (z_out_38[10]), {nor_204_cse , (fsm_output[34]) , or_dcpl_1191});
  assign mux1h_16_nl = MUX1HOT_v_5_3_2((z_out_45[9:5]), reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd,
      (z_out_38[9:5]), {nor_204_cse , (fsm_output[34]) , or_dcpl_1191});
  assign mux1h_17_nl = MUX1HOT_v_5_3_2((z_out_45[4:0]), reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1,
      (z_out_38[4:0]), {nor_204_cse , (fsm_output[34]) , or_dcpl_1191});
  assign out_u_rsci_d_d = {mux1h_10_nl , mux1h_11_nl , mux1h_15_nl , mux1h_16_nl
      , mux1h_17_nl};
  assign out_u_rsci_we_d_pff = (nor_3_cse & or_dcpl_99) | (stage_PE_1_and_cse & or_200_cse);
  assign out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = (~(mode_lpi_1_dfm | (~((fsm_output[4:3]!=2'b00)))))
      | (operator_16_false_operator_16_false_nor_cse_sva & (fsm_output[53]));
  assign or_tmp = (return_add_generic_AC_RND_CONV_false_10_exception_sva_1 & (fsm_output[22]))
      | (return_add_generic_AC_RND_CONV_false_exception_sva_1 & (fsm_output[6]))
      | (return_add_generic_AC_RND_CONV_false_12_exception_sva_1 & (fsm_output[26]))
      | (return_add_generic_AC_RND_CONV_false_9_exception_sva_1 & (fsm_output[20]))
      | (return_add_generic_AC_RND_CONV_false_11_exception_sva_1 & (fsm_output[24]))
      | (return_add_generic_AC_RND_CONV_false_1_exception_sva_1 & (fsm_output[8]));
  assign or_tmp_916 = ((~(return_add_generic_AC_RND_CONV_false_10_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0))
      & (fsm_output[22])) | ((~(return_add_generic_AC_RND_CONV_false_12_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx1w0))
      & (fsm_output[26])) | ((~(return_add_generic_AC_RND_CONV_false_9_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx1w0))
      & (fsm_output[20])) | ((~(return_add_generic_AC_RND_CONV_false_11_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0))
      & (fsm_output[24]));
  assign or_tmp_917 = ((~ return_add_generic_AC_RND_CONV_false_10_exception_sva_1)
      & return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0 & (fsm_output[22]))
      | ((~ return_add_generic_AC_RND_CONV_false_12_exception_sva_1) & return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx1w0
      & (fsm_output[26])) | ((~ return_add_generic_AC_RND_CONV_false_9_exception_sva_1)
      & return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx1w0 & (fsm_output[20]))
      | ((~ return_add_generic_AC_RND_CONV_false_11_exception_sva_1) & return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0
      & (fsm_output[24]));
  assign or_tmp_919 = BUTTERFLY_if_1_if_and_9_cse | BUTTERFLY_if_1_if_and_5_cse |
      BUTTERFLY_if_1_if_and_11_cse | BUTTERFLY_if_1_if_and_8_cse | BUTTERFLY_if_1_if_and_10_cse
      | BUTTERFLY_if_1_if_and_6_cse;
  assign or_tmp_920 = (return_add_generic_AC_RND_CONV_false_13_exception_sva_1 &
      (fsm_output[31])) | (return_add_generic_AC_RND_CONV_false_23_exception_sva_1
      & (fsm_output[47])) | (return_add_generic_AC_RND_CONV_false_25_exception_sva_1
      & (fsm_output[51])) | (return_add_generic_AC_RND_CONV_false_22_exception_sva_1
      & (fsm_output[45])) | (return_add_generic_AC_RND_CONV_false_24_exception_sva_1
      & (fsm_output[49])) | (return_add_generic_AC_RND_CONV_false_14_exception_sva_1
      & (fsm_output[33]));
  assign or_tmp_921 = ((~(return_add_generic_AC_RND_CONV_false_23_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0))
      & (fsm_output[47])) | ((~(return_add_generic_AC_RND_CONV_false_25_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0))
      & (fsm_output[51])) | ((~(return_add_generic_AC_RND_CONV_false_22_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0))
      & (fsm_output[45])) | ((~(return_add_generic_AC_RND_CONV_false_24_exception_sva_1
      | reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd | return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx1w0))
      & (fsm_output[49]));
  assign or_tmp_922 = ((~ return_add_generic_AC_RND_CONV_false_23_exception_sva_1)
      & return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0 & (fsm_output[47]))
      | ((~ return_add_generic_AC_RND_CONV_false_25_exception_sva_1) & return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0
      & (fsm_output[51])) | ((~ return_add_generic_AC_RND_CONV_false_22_exception_sva_1)
      & return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0 & (fsm_output[45]))
      | ((~ return_add_generic_AC_RND_CONV_false_24_exception_sva_1) & return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx1w0
      & (fsm_output[49]));
  assign or_tmp_924 = BUTTERFLY_if_1_and_7_cse | BUTTERFLY_if_1_and_11_cse | BUTTERFLY_if_1_and_13_cse
      | BUTTERFLY_if_1_and_10_cse | BUTTERFLY_if_1_and_12_cse | BUTTERFLY_if_1_and_8_cse;
  assign return_add_generic_AC_RND_CONV_false_e_r_qelse_not_5_nl = ~ return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
  assign return_add_generic_AC_RND_CONV_false_e_r_return_add_generic_AC_RND_CONV_false_e_r_or_cse
      = MUX_v_10_2_2(10'b0000000000, z_out_10, return_add_generic_AC_RND_CONV_false_e_r_qelse_not_5_nl);
  assign return_add_generic_AC_RND_CONV_false_1_e_r_qelse_not_3_nl = ~ return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs_mx1w0;
  assign return_add_generic_AC_RND_CONV_false_1_e_r_return_add_generic_AC_RND_CONV_false_1_e_r_or_cse
      = MUX_v_10_2_2(10'b0000000000, z_out_10, return_add_generic_AC_RND_CONV_false_1_e_r_qelse_not_3_nl);
  assign or_tmp_927 = (fsm_output[6]) | (fsm_output[8]) | (fsm_output[31]) | (fsm_output[33]);
  assign or_tmp_929 = (fsm_output[12]) | (fsm_output[18]) | (fsm_output[37]) | (fsm_output[43]);
  assign or_tmp_930 = (fsm_output[14]) | (fsm_output[16]) | (fsm_output[39]) | (fsm_output[41]);
  assign or_tmp_940 = inverse_lpi_1_dfm_1 & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  assign or_tmp_979 = ~(inverse_lpi_1_dfm_1 | and_dcpl_284);
  assign or_tmp_983 = (fsm_output[42]) | (fsm_output[36]) | (fsm_output[17]) | (fsm_output[11]);
  assign or_tmp_1248 = (fsm_output[31]) | (fsm_output[6]) | (fsm_output[8]) | (fsm_output[33])
      | (fsm_output[29]) | (fsm_output[4]);
  assign or_tmp_1249 = (fsm_output[44]) | (fsm_output[16]) | (fsm_output[41]);
  assign or_tmp_1250 = (fsm_output[20]) | (fsm_output[17]);
  assign or_tmp_1251 = (fsm_output[40]) | (fsm_output[42]) | (fsm_output[45]) | (fsm_output[15]);
  assign BUTTERFLY_1_else_1_if_and_ssc = run_wen & (~(return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse
      | or_dcpl_401));
  assign BUTTERFLY_1_else_1_if_and_3_cse = ~((fsm_output[37]) | (~(or_dcpl_407 |
      or_dcpl_404 | (fsm_output[11]))));
  assign BUTTERFLY_1_else_1_if_and_1_cse = BUTTERFLY_1_else_1_if_and_ssc & (~(or_dcpl_423
      | or_dcpl_618));
  assign return_add_generic_AC_RND_CONV_false_15_op_bigger_and_ssc = run_wen & (~
      or_tmp_403);
  assign return_add_generic_AC_RND_CONV_false_17_m_r_and_ssc = run_wen & (~(or_dcpl_425
      | or_dcpl_618 | or_dcpl_401 | or_dcpl_417));
  assign BUTTERFLY_1_else_2_or_cse = or_38_cse | ((~ mode_lpi_1_dfm) & or_dcpl_401);
  assign BUTTERFLY_1_else_2_and_27_cse = (~ inverse_lpi_1_dfm_1) & return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse;
  assign and_1153_rgt = or_590_cse & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  assign BUTTERFLY_1_else_2_and_46_cse = run_wen & (~(or_dcpl_108 | (fsm_output[50])
      | or_dcpl_534 | or_dcpl_531 | (fsm_output[19]) | or_dcpl_133)) & ((~ or_1670_ssc)
      | or_tmp_561 | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
      | or_tmp_564 | return_add_generic_AC_RND_CONV_false_17_e_r_and_cse | or_1673_ssc
      | and_1598_cse | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_34_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse | or_tmp_570
      | or_1678_ssc | and_1608_cse | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse
      | and_1153_rgt | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_6_cse
      | or_tmp_348 | return_add_generic_AC_RND_CONV_false_11_exp_and_3_cse | and_1163_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_16_cse | BUTTERFLY_1_else_2_or_cse
      | BUTTERFLY_1_else_2_and_27_cse);
  assign BUTTERFLY_1_else_3_else_and_1_ssc = BUTTERFLY_1_else_3_else_and_ssc & (~
      or_38_cse);
  assign BUTTERFLY_1_else_3_else_and_11_cse = (~ mode_lpi_1_dfm) & return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse;
  assign BUTTERFLY_1_else_3_else_or_rgt = (mode_lpi_1_dfm & return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse)
      | (inverse_lpi_1_dfm_1 & return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse)
      | or_dcpl_423 | (fsm_output[35]) | or_dcpl_514;
  assign BUTTERFLY_1_else_3_else_and_26_cse = or_tmp_561 & BUTTERFLY_1_else_3_else_or_rgt;
  assign BUTTERFLY_1_else_3_else_and_27_cse = (and_1615_cse | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse)
      & BUTTERFLY_1_else_3_else_or_rgt;
  assign BUTTERFLY_1_else_3_else_and_28_cse = (return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse) & BUTTERFLY_1_else_3_else_or_rgt;
  assign BUTTERFLY_1_else_3_else_and_30_cse = (return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse
      | and_1626_cse) & BUTTERFLY_1_else_3_else_or_rgt;
  assign BUTTERFLY_1_else_3_else_and_24_cse = BUTTERFLY_1_else_3_else_and_1_ssc &
      (~(or_dcpl_662 | or_dcpl_976 | or_dcpl_126 | or_dcpl_788 | or_dcpl_125 | (fsm_output[19])))
      & (~ or_tmp_403);
  assign stage_PE_1_tmp_im_d_and_ssc = run_wen & ((inverse_lpi_1_dfm_1 & (~(or_dcpl_586
      | or_dcpl_693))) | (fsm_output[4]) | stage_PE_1_tmp_im_d_1_sva_1_mx0c3 | (fsm_output[29]));
  assign stage_PE_1_tmp_re_d_or_4_rgt = stage_PE_1_tmp_re_d_1_sva_1_mx0c0 | return_extract_26_exception_or_3_cse
      | (inverse_lpi_1_dfm_1 & (fsm_output[7])) | (inverse_lpi_1_dfm_1 & (fsm_output[32]));
  assign stage_PE_1_tmp_re_d_and_5_rgt = (~ inverse_lpi_1_dfm_1) & (fsm_output[7]);
  assign stage_PE_1_tmp_re_d_and_7_rgt = (~ inverse_lpi_1_dfm_1) & (fsm_output[32]);
  assign stage_PE_1_tmp_re_d_or_6_cse = (~(or_dcpl_976 | or_dcpl_125 | (fsm_output[33])
      | (fsm_output[32]) | (fsm_output[8]) | (fsm_output[7]) | (fsm_output[18])))
      | stage_PE_1_tmp_re_d_and_5_rgt | stage_PE_1_tmp_re_d_and_7_rgt;
  assign return_add_generic_AC_RND_CONV_false_4_mux_24_cse = MUX_v_56_2_2((z_out_43[56:1]),
      (~ (z_out_43[56:1])), return_add_generic_AC_RND_CONV_false_17_do_sub_sva_1);
  assign return_add_generic_AC_RND_CONV_false_5_mux_18_cse = MUX_v_56_2_2((z_out_43[56:1]),
      (~ (z_out_43[56:1])), return_add_generic_AC_RND_CONV_false_10_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_res_mant_conc_2_itm_56_1 = MUX_v_56_2_2((z_out_43[56:1]),
      (~ (z_out_43[56:1])), xor_cse);
  assign return_add_generic_AC_RND_CONV_false_conc_6_itm_54_4 = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx1,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse);
  assign BUTTERFLY_else_1_BUTTERFLY_else_1_and_cse = MUX_v_2_2_2(2'b00, (z_out_3[17:16]),
      inverse_lpi_1_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_5_mux_19_cse = MUX_v_56_2_2((z_out_43[56:1]),
      (~ (z_out_43[56:1])), return_add_generic_AC_RND_CONV_false_11_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_12_mux_19_cse = MUX_v_56_2_2((z_out_43[56:1]),
      (~ (z_out_43[56:1])), return_add_generic_AC_RND_CONV_false_14_op2_nan_sva);
  assign return_add_generic_AC_RND_CONV_false_23_conc_6_itm_53_4 = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[49:0]),
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_25_op1_smaller_return_add_generic_AC_RND_CONV_false_25_op1_smaller_or_cse);
  assign return_add_generic_AC_RND_CONV_false_1_res_mant_conc_2_itm_56_1 = MUX_v_56_2_2((z_out_43[56:1]),
      (~ (z_out_43[56:1])), xor_2_cse);
  assign return_add_generic_AC_RND_CONV_false_1_conc_6_itm_54_4 = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx1, return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse);
  assign return_add_generic_AC_RND_CONV_false_5_mux_20_cse = MUX_v_56_2_2((z_out_43[56:1]),
      (~ (z_out_43[56:1])), return_add_generic_AC_RND_CONV_false_16_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_6_mux_33_cse = MUX_v_56_2_2((~ (z_out_43[56:1])),
      (z_out_43[56:1]), not_tmp_302);
  assign return_add_generic_AC_RND_CONV_false_6_conc_6_itm_53_4 = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm,
      return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_49_0_mx0, or_918_cse);
  assign return_add_generic_AC_RND_CONV_false_8_res_mant_conc_7_itm_56_1 = MUX_v_56_2_2((z_out_43[56:1]),
      (~ (z_out_43[56:1])), return_add_generic_AC_RND_CONV_false_14_op2_inf_sva);
  assign return_add_generic_AC_RND_CONV_false_10_conc_6_itm_53_4 = MUX_v_50_2_2((return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49:0]),
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse);
  assign return_add_generic_AC_RND_CONV_false_14_res_mant_conc_2_itm_56_1 = MUX_v_56_2_2((z_out_43[56:1]),
      (~ (z_out_43[56:1])), xor_4_cse);
  assign return_add_generic_AC_RND_CONV_false_14_conc_6_itm_54_4 = MUX_v_51_2_2(return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm,
      return_extract_32_mux_4_cse, return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse);
  assign return_add_generic_AC_RND_CONV_false_19_conc_6_itm_53_4 = MUX_v_50_2_2(return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm,
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_49_0_mx0, or_920_cse);
  assign return_add_generic_AC_RND_CONV_false_12_mux_21_cse = MUX_v_56_2_2((z_out_43[56:1]),
      (~ (z_out_43[56:1])), return_add_generic_AC_RND_CONV_false_12_do_sub_sva);
  assign return_add_generic_AC_RND_CONV_false_13_res_mant_conc_2_itm_56_1 = MUX_v_56_2_2((z_out_43[56:1]),
      (~ (z_out_43[56:1])), xor_3_cse);
  assign return_add_generic_AC_RND_CONV_false_13_conc_6_itm_54_4 = MUX_v_51_2_2(return_extract_32_mux_4_cse,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse);
  assign return_mult_generic_AC_RND_CONV_false_6_op1_normal_not_5_nl = ~ return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp;
  assign return_mult_generic_AC_RND_CONV_false_6_if_conc_itm_51_0 = MUX_v_52_2_2(52'b0000000000000000000000000000000000000000000000000000,
      (out_f_d_rsci_q_d[51:0]), return_mult_generic_AC_RND_CONV_false_6_op1_normal_not_5_nl);
  assign operator_6_false_1_or_1_ssc = or_dcpl_548 | or_tmp_930;
  assign operator_6_false_1_or_8_cse = (fsm_output[20]) | (fsm_output[51]);
  assign operator_6_false_1_or_4_cse = (fsm_output[24]) | (fsm_output[47]);
  assign operator_6_false_1_or_6_cse = (fsm_output[26]) | (fsm_output[49]);
  assign operator_6_false_or_3_ssc = or_dcpl_780 | or_dcpl_423 | return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse;
  assign operator_6_false_or_15_cse = (fsm_output[19]) | (fsm_output[50]);
  assign operator_6_false_or_6_cse = (fsm_output[21]) | (fsm_output[44]);
  assign operator_6_false_or_12_cse = (fsm_output[25]) | (fsm_output[48]);
  assign operator_6_false_or_ssc = or_dcpl_780 | (fsm_output[23]) | (fsm_output[44])
      | (fsm_output[50]);
  assign operator_6_false_or_1_ssc = or_tmp_983 | or_dcpl_423 | (fsm_output[21])
      | (fsm_output[46]);
  assign return_add_generic_AC_RND_CONV_false_4_or_ssc = (fsm_output[9]) | (fsm_output[19])
      | (fsm_output[23]) | (fsm_output[34]) | (fsm_output[46]);
  assign return_add_generic_AC_RND_CONV_false_4_or_20_ssc = (fsm_output[3]) | or_38_cse
      | (fsm_output[5]) | return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
      | (fsm_output[28]) | (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_4_or_18_ssc = return_extract_26_exception_or_3_cse
      | (fsm_output[11]) | (fsm_output[13]) | (fsm_output[17]) | (fsm_output[21])
      | (fsm_output[36]) | (fsm_output[38]) | (fsm_output[42]) | (fsm_output[44])
      | (fsm_output[48]);
  assign BUTTERFLY_i_nor_2_cse_1 = ~(return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      | (fsm_output[5]) | (fsm_output[30]));
  assign BUTTERFLY_i_or_4_cse = (fsm_output[14]) | (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_or_6_cse = (fsm_output[7])
      | (fsm_output[18]) | (fsm_output[32]) | (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_4_or_35_cse = or_38_cse | (fsm_output[43])
      | (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_4_or_33_cse = or_dcpl_401 | (fsm_output[19])
      | (fsm_output[42]);
  assign return_add_generic_AC_RND_CONV_false_4_or_43_cse = (fsm_output[17]) | (fsm_output[44]);
  assign return_add_generic_AC_RND_CONV_false_4_or_47_cse = return_extract_26_exception_or_3_cse
      | return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_27_cse = (fsm_output[17]) | return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse
      | (fsm_output[44]) | (fsm_output[20]);
  assign return_add_generic_AC_RND_CONV_false_4_or_31_cse = (fsm_output[19]) | (fsm_output[42])
      | (fsm_output[45]) | return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse;
  assign return_add_generic_AC_RND_CONV_false_e_dif1_or_1_ssc = (fsm_output[7]) |
      (fsm_output[18]) | (fsm_output[32]);
  assign return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_or_cse
      = ((z_out_21[105]) & (~ (z_out_17[52]))) | ((z_out_21[104]) & (~ (z_out_17[51])))
      | ((z_out_21[103]) & (~ (z_out_17[50]))) | ((z_out_21[102]) & (~ (z_out_17[49])))
      | ((z_out_21[101]) & (~ (z_out_17[48]))) | ((z_out_21[100]) & (~ (z_out_17[47])))
      | ((z_out_21[99]) & (~ (z_out_17[46]))) | ((z_out_21[98]) & (~ (z_out_17[45])))
      | ((z_out_21[97]) & (~ (z_out_17[44]))) | ((z_out_21[96]) & (~ (z_out_17[43])))
      | ((z_out_21[95]) & (~ (z_out_17[42]))) | ((z_out_21[94]) & (~ (z_out_17[41])))
      | ((z_out_21[93]) & (~ (z_out_17[40]))) | ((z_out_21[92]) & (~ (z_out_17[39])))
      | ((z_out_21[91]) & (~ (z_out_17[38]))) | ((z_out_21[90]) & (~ (z_out_17[37])))
      | ((z_out_21[89]) & (~ (z_out_17[36]))) | ((z_out_21[88]) & (~ (z_out_17[35])))
      | ((z_out_21[87]) & (~ (z_out_17[34]))) | ((z_out_21[86]) & (~ (z_out_17[33])))
      | ((z_out_21[85]) & (~ (z_out_17[32]))) | ((z_out_21[84]) & (~ (z_out_17[31])))
      | ((z_out_21[83]) & (~ (z_out_17[30]))) | ((z_out_21[82]) & (~ (z_out_17[29])))
      | ((z_out_21[81]) & (~ (z_out_17[28]))) | ((z_out_21[80]) & (~ (z_out_17[27])))
      | ((z_out_21[79]) & (~ (z_out_17[26]))) | ((z_out_21[78]) & (~ (z_out_17[25])))
      | ((z_out_21[77]) & (~ (z_out_17[24]))) | ((z_out_21[76]) & (~ (z_out_17[23])))
      | ((z_out_21[75]) & (~ (z_out_17[22]))) | ((z_out_21[74]) & (~ (z_out_17[21])))
      | ((z_out_21[73]) & (~ (z_out_17[20]))) | ((z_out_21[72]) & (~ (z_out_17[19])))
      | ((z_out_21[71]) & (~ (z_out_17[18]))) | ((z_out_21[70]) & (~ (z_out_17[17])))
      | ((z_out_21[69]) & (~ (z_out_17[16]))) | ((z_out_21[68]) & (~ (z_out_17[15])))
      | ((z_out_21[67]) & (~ (z_out_17[14]))) | ((z_out_21[66]) & (~ (z_out_17[13])))
      | ((z_out_21[65]) & (~ (z_out_17[12]))) | ((z_out_21[64]) & (~ (z_out_17[11])))
      | ((z_out_21[63]) & (~ (z_out_17[10]))) | ((z_out_21[62]) & (~ (z_out_17[9])))
      | ((z_out_21[61]) & (~ (z_out_17[8]))) | ((z_out_21[60]) & (~ (z_out_17[7])))
      | ((z_out_21[59]) & (~ (z_out_17[6]))) | ((z_out_21[58]) & (~ (z_out_17[5])))
      | ((z_out_21[57]) & (~ (z_out_17[4]))) | ((z_out_21[56]) & (~ (z_out_17[3])))
      | ((z_out_21[55]) & (~ (z_out_17[2]))) | ((z_out_21[54]) & (~ (z_out_17[1])))
      | ((z_out_21[53]) & (~ (z_out_17[0]))) | (z_out_21[52:0]!=53'b00000000000000000000000000000000000000000000000000000);
  assign operator_6_false_8_nor_1_cse = ~((fsm_output[3]) | or_38_cse | (fsm_output[28]));
  assign operator_6_false_or_20_cse = (fsm_output[19]) | (fsm_output[25]) | (fsm_output[48]);
  assign return_add_generic_AC_RND_CONV_false_20_ma1_lt_ma2_mux_1_cse = MUX_s_1_2_2((~
      return_mult_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_mx1), (~ return_mult_generic_AC_RND_CONV_false_2_m_r_51_lpi_3_dfm_mx1),
      fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_20_ma1_lt_ma2_mux_4_cse = MUX_v_51_2_2((~
      return_mult_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1), (~ return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1),
      fsm_output[14]);
  assign BUTTERFLY_1_else_1_if_BUTTERFLY_1_else_1_if_mux_2_cse = MUX_s_1_2_2((z_out_37[17]),
      (z_out_45[17]), return_extract_26_exception_or_3_cse);
  assign return_add_generic_AC_RND_CONV_false_4_or_86_cse = (fsm_output[19]) | or_tmp_1249;
  assign return_add_generic_AC_RND_CONV_false_4_or_87_cse = or_tmp_1250 | or_tmp_1251;
  assign return_add_generic_AC_RND_CONV_false_4_res_rounded_or_1_cse = (fsm_output[3])
      | or_38_cse | (fsm_output[5]) | (fsm_output[9]) | (fsm_output[11]) | (fsm_output[13])
      | (fsm_output[15]) | (fsm_output[17]) | (fsm_output[19]) | (fsm_output[21])
      | (fsm_output[23]) | (fsm_output[25]) | (fsm_output[30]) | (fsm_output[34])
      | (fsm_output[36]) | (fsm_output[38]) | (fsm_output[40]) | (fsm_output[42])
      | (fsm_output[44]) | (fsm_output[46]) | (fsm_output[48]) | (fsm_output[50])
      | return_extract_26_exception_or_3_cse | (fsm_output[28]);
  assign return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_or_1_cse
      = (fsm_output[10]) | (fsm_output[12]) | (fsm_output[14]) | (fsm_output[35])
      | (fsm_output[37]) | (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_4_or_99_cse = or_38_cse | or_dcpl_401
      | return_extract_26_exception_or_3_cse;
  assign return_add_generic_AC_RND_CONV_false_4_and_105_cse = (~ or_590_cse) & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_97_cse = (fsm_output[5]) | (fsm_output[30])
      | (fsm_output[37]);
  assign return_add_generic_AC_RND_CONV_false_4_or_95_cse = (fsm_output[19]) | or_tmp_1248
      | or_tmp_1249;
  assign return_add_generic_AC_RND_CONV_false_4_and_5_cse = (~ return_add_generic_AC_RND_CONV_false_9_acc_2_itm_11_1)
      & (fsm_output[19]);
  assign return_add_generic_AC_RND_CONV_false_4_and_13_cse = (~ return_add_generic_AC_RND_CONV_false_22_acc_2_itm_11_1)
      & (fsm_output[44]);
  assign return_add_generic_AC_RND_CONV_false_4_or_52_cse = (return_add_generic_AC_RND_CONV_false_9_acc_2_itm_11_1
      & (fsm_output[19])) | (return_add_generic_AC_RND_CONV_false_12_acc_2_itm_11_1
      & (fsm_output[25])) | (return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11_1
      & (fsm_output[48]));
  assign return_add_generic_AC_RND_CONV_false_4_and_7_cse = (~ return_add_generic_AC_RND_CONV_false_10_acc_2_itm_11_1)
      & (fsm_output[21]);
  assign return_add_generic_AC_RND_CONV_false_4_and_15_cse = (~ return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1)
      & (fsm_output[46]);
  assign return_add_generic_AC_RND_CONV_false_4_or_54_cse = (return_add_generic_AC_RND_CONV_false_10_acc_2_itm_11_1
      & (fsm_output[21])) | (return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1
      & (fsm_output[46]));
  assign return_add_generic_AC_RND_CONV_false_4_and_9_cse = (~ return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1)
      & (fsm_output[23]);
  assign return_add_generic_AC_RND_CONV_false_4_and_17_cse = (~ return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11_1)
      & (fsm_output[48]);
  assign return_add_generic_AC_RND_CONV_false_4_or_56_cse = (return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1
      & (fsm_output[23])) | (return_add_generic_AC_RND_CONV_false_22_acc_2_itm_11_1
      & (fsm_output[44])) | (return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11_1
      & (fsm_output[50]));
  assign return_add_generic_AC_RND_CONV_false_4_and_11_cse = (~ return_add_generic_AC_RND_CONV_false_12_acc_2_itm_11_1)
      & (fsm_output[25]);
  assign return_add_generic_AC_RND_CONV_false_4_and_19_cse = (~ return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11_1)
      & (fsm_output[50]);
  assign return_add_generic_AC_RND_CONV_false_4_and_67_cse = (~ return_add_generic_AC_RND_CONV_false_25_op1_smaller_return_add_generic_AC_RND_CONV_false_25_op1_smaller_or_cse)
      & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_4_and_71_cse = (~ or_918_cse) & (fsm_output[12]);
  assign return_add_generic_AC_RND_CONV_false_4_and_77_cse = (~ or_920_cse) & (fsm_output[37]);
  assign return_add_generic_AC_RND_CONV_false_4_and_73_cse = (~ return_add_generic_AC_RND_CONV_false_12_op1_smaller_return_add_generic_AC_RND_CONV_false_12_op1_smaller_or_cse)
      & (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_4_or_70_cse = ((~ return_add_generic_AC_RND_CONV_false_2_op1_smaller_return_add_generic_AC_RND_CONV_false_2_op1_smaller_or_cse)
      & (fsm_output[5])) | and_1615_cse;
  assign return_add_generic_AC_RND_CONV_false_4_and_69_cse = (~ return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse)
      & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_4_and_75_cse = (~ return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse)
      & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_4_or_73_cse = and_1626_cse | ((~ return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse)
      & (fsm_output[30]));
  assign or_dcpl_1189 = (fsm_output[5]) | (fsm_output[8]);
  assign or_dcpl_1191 = (fsm_output[30]) | (fsm_output[33]);
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_or_cse = return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      | ((~ inverse_lpi_1_dfm_1) & (fsm_output[37]));
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_and_1_cse = inverse_lpi_1_dfm_1
      & (fsm_output[37]);
  assign return_add_generic_AC_RND_CONV_false_5_conc_itm_3_0 = MUX_v_4_2_2(reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2,
      (rtn_out[4:1]), return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1);
  assign return_add_generic_AC_RND_CONV_false_2_conc_68_itm_3_0 = MUX_v_4_2_2(reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2,
      (return_add_generic_AC_RND_CONV_false_11_ls_sva[4:1]), return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_2_conc_69_itm_3_0 = MUX_v_4_2_2(reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2,
      (return_add_generic_AC_RND_CONV_false_10_ls_sva[4:1]), return_add_generic_AC_RND_CONV_false_19_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_2_conc_70_itm_3_0 = MUX_v_4_2_2(reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2,
      (rtn_out[4:1]), return_add_generic_AC_RND_CONV_false_20_acc_3_itm_11_1);
  assign return_add_generic_AC_RND_CONV_false_4_or_51_itm = return_add_generic_AC_RND_CONV_false_4_and_5_cse
      | return_add_generic_AC_RND_CONV_false_4_and_19_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_53_itm = return_add_generic_AC_RND_CONV_false_4_and_7_cse
      | return_add_generic_AC_RND_CONV_false_4_and_13_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_55_itm = return_add_generic_AC_RND_CONV_false_4_and_9_cse
      | return_add_generic_AC_RND_CONV_false_4_and_15_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_57_itm = return_add_generic_AC_RND_CONV_false_4_and_11_cse
      | return_add_generic_AC_RND_CONV_false_4_and_17_cse;
  assign return_add_generic_AC_RND_CONV_false_2_or_2_seb = (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[16]) | (fsm_output[30]) | (fsm_output[32]) | (fsm_output[41]);
  assign BUTTERFLY_1_nor_1_seb = ~((fsm_output[5]) | (fsm_output[30]));
  assign BUTTERFLY_i_conc_3_itm_10_9 = MUX_v_2_2_2(BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1,
      (z_out_3[10:9]), inverse_lpi_1_dfm_1);
  assign BUTTERFLY_i_conc_3_itm_8_0 = MUX_v_9_2_2(BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2,
      (z_out_3[8:0]), inverse_lpi_1_dfm_1);
  assign return_mult_generic_AC_RND_CONV_false_exp_or_4_itm = (fsm_output[10]) |
      (fsm_output[12]) | (fsm_output[35]) | (fsm_output[37]);
  assign nl_operator_6_false_8_acc_itm = ({1'b1 , (~ (rtn_out[5:1]))}) + 6'b000001;
  assign operator_6_false_8_acc_itm = nl_operator_6_false_8_acc_itm[5:0];
  assign nl_exs_26_itm_5_0 = ({1'b1 , (~ (rtn_out[5:1]))}) + 6'b000001;
  assign exs_26_itm_5_0 = nl_exs_26_itm_5_0[5:0];
  assign nl_exs_27_itm_5_0 = ({1'b1 , (~ (rtn_out[5:1]))}) + 6'b000001;
  assign exs_27_itm_5_0 = nl_exs_27_itm_5_0[5:0];
  assign return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_and_cse
      = (z_out_21[105]) & (~ (fsm_output[54]));
  assign return_mult_generic_AC_RND_CONV_false_if_1_return_mult_generic_AC_RND_CONV_false_if_1_mux_2_cse
      = MUX_s_1_2_2((z_out_21[104]), return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp,
      fsm_output[54]);
  assign return_add_generic_AC_RND_CONV_false_4_or_112_cse = ((~ return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1)
      & or_38_cse) | ((~ return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1)
      & or_dcpl_780) | ((~ return_add_generic_AC_RND_CONV_false_19_acc_3_itm_11_1)
      & or_dcpl_423) | ((~ return_add_generic_AC_RND_CONV_false_20_acc_3_itm_11_1)
      & return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse);
  assign return_add_generic_AC_RND_CONV_false_4_or_113_cse = (return_add_generic_AC_RND_CONV_false_18_acc_3_itm_10_1
      & or_38_cse) | (return_add_generic_AC_RND_CONV_false_20_acc_3_itm_11_1 & return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse);
  assign return_add_generic_AC_RND_CONV_false_4_or_116_cse = (return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1
      & or_dcpl_780) | return_add_generic_AC_RND_CONV_false_4_or_56_cse;
  assign return_add_generic_AC_RND_CONV_false_4_and_132_cse = return_add_generic_AC_RND_CONV_false_19_acc_3_itm_11_1
      & or_dcpl_423;
  assign return_mult_generic_AC_RND_CONV_false_1_if_mux_6_tmp = MUX_s_1_2_2(return_extract_13_return_extract_13_or_1_cse_sva_1,
      return_extract_45_return_extract_45_or_1_cse_sva_1, fsm_output[37]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      out1_rsci_idat_63 <= 1'b0;
      out1_rsci_idat_62_52 <= 11'b00000000000;
      out1_rsci_idat_51 <= 1'b0;
      out1_rsci_idat_50_0 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      out1_rsci_idat_63 <= 1'b0;
      out1_rsci_idat_62_52 <= 11'b00000000000;
      out1_rsci_idat_51 <= 1'b0;
      out1_rsci_idat_50_0 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( for_1_if_and_ssc ) begin
      out1_rsci_idat_63 <= MUX_s_1_2_2((out_f_d_rsci_q_d[63]), (in_f_d_rsci_q_d[63]),
          out1_rsci_idat_63_0_mx0c2);
      out1_rsci_idat_62_52 <= MUX1HOT_v_11_3_2((out_f_d_rsci_q_d[62:52]), return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_or_nl,
          (in_f_d_rsci_q_d[62:52]), {or_tmp_61 , out1_rsci_idat_63_0_mx0c1 , out1_rsci_idat_63_0_mx0c2});
      out1_rsci_idat_51 <= MUX1HOT_s_1_4_2((out_f_d_rsci_q_d[51]), (z_out_6[51]),
          return_mult_generic_AC_RND_CONV_false_6_op1_nan_sva_1, (in_f_d_rsci_q_d[51]),
          {or_tmp_61 , BUTTERFLY_if_1_and_nl , BUTTERFLY_if_1_and_1_nl , out1_rsci_idat_63_0_mx0c2});
      out1_rsci_idat_50_0 <= MUX1HOT_v_51_3_2((out_f_d_rsci_q_d[50:0]), return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_and_1_nl,
          (in_f_d_rsci_q_d[50:0]), {or_tmp_61 , out1_rsci_idat_63_0_mx0c1 , out1_rsci_idat_63_0_mx0c2});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      out1_rsci_idat_79_64 <= 16'b0000000000000000;
    end
    else if ( rst ) begin
      out1_rsci_idat_79_64 <= 16'b0000000000000000;
    end
    else if ( run_wen & (or_tmp_61 | out1_rsci_idat_79_64_mx0c1 | and_571_cse) )
        begin
      out1_rsci_idat_79_64 <= MUX1HOT_v_16_3_2(out_u_rsci_q_d, in_u_rsci_q_d, ({{1{stage_monty_mul_acc_2_psp_sva_1[14]}},
          stage_monty_mul_acc_2_psp_sva_1}), {or_tmp_61 , out1_rsci_idat_79_64_mx0c1
          , and_571_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_out_u_triosy_obj_iswt0_cse <= 1'b0;
      reg_out1_rsci_iswt0_cse <= 1'b0;
      reg_out_u_rsci_cgo_ir_cse <= 1'b0;
      reg_out_f_d_rsci_cgo_ir_cse <= 1'b0;
      reg_in_u_rsci_cgo_ir_cse <= 1'b0;
      reg_in_f_d_rsci_cgo_ir_cse <= 1'b0;
      reg_ap_start_rsci_iswt0_cse <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva
          <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd <= 1'b0;
      BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_0 <= 6'b000000;
    end
    else if ( rst ) begin
      reg_out_u_triosy_obj_iswt0_cse <= 1'b0;
      reg_out1_rsci_iswt0_cse <= 1'b0;
      reg_out_u_rsci_cgo_ir_cse <= 1'b0;
      reg_out_f_d_rsci_cgo_ir_cse <= 1'b0;
      reg_in_u_rsci_cgo_ir_cse <= 1'b0;
      reg_in_f_d_rsci_cgo_ir_cse <= 1'b0;
      reg_ap_start_rsci_iswt0_cse <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva
          <= 1'b0;
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd <= 1'b0;
      BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_0 <= 6'b000000;
    end
    else if ( run_wen ) begin
      reg_out_u_triosy_obj_iswt0_cse <= (z_out_19[10]) & (fsm_output[55]);
      reg_out1_rsci_iswt0_cse <= fsm_output[54];
      reg_out_u_rsci_cgo_ir_cse <= or_1178_rmff;
      reg_out_f_d_rsci_cgo_ir_cse <= or_1179_rmff;
      reg_in_u_rsci_cgo_ir_cse <= or_1180_rmff;
      reg_in_f_d_rsci_cgo_ir_cse <= or_1181_rmff;
      reg_ap_start_rsci_iswt0_cse <= ~ and_dcpl_165;
      return_add_generic_AC_RND_CONV_false_10_if_4_slc_return_add_generic_AC_RND_CONV_false_10_acc_2_11_mdf_sva
          <= MUX1HOT_s_1_18_2(return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp,
          return_add_generic_AC_RND_CONV_false_acc_2_itm_11_1, return_add_generic_AC_RND_CONV_false_1_acc_2_itm_11_1,
          return_add_generic_AC_RND_CONV_false_15_acc_3_itm_11_1, return_add_generic_AC_RND_CONV_false_8_acc_3_itm_11_1,
          return_add_generic_AC_RND_CONV_false_19_acc_3_itm_11_1, return_add_generic_AC_RND_CONV_false_20_acc_3_itm_11_1,
          return_add_generic_AC_RND_CONV_false_9_acc_2_itm_11_1, return_add_generic_AC_RND_CONV_false_10_acc_2_itm_11_1,
          return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1, return_add_generic_AC_RND_CONV_false_12_acc_2_itm_11_1,
          return_add_generic_AC_RND_CONV_false_13_return_add_generic_AC_RND_CONV_false_13_or_1_tmp,
          return_add_generic_AC_RND_CONV_false_13_acc_2_itm_11_1, return_add_generic_AC_RND_CONV_false_14_acc_2_itm_11_1,
          return_add_generic_AC_RND_CONV_false_22_acc_2_itm_11_1, return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1,
          return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11_1, return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11_1,
          {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , or_dcpl_780 , or_1606_nl
          , or_dcpl_423 , return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
          , (fsm_output[19]) , (fsm_output[21]) , (fsm_output[23]) , (fsm_output[25])
          , (fsm_output[29]) , (fsm_output[30]) , (fsm_output[32]) , (fsm_output[44])
          , (fsm_output[46]) , (fsm_output[48]) , (fsm_output[50])});
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd <= z_out_6[53];
      BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_0 <= MUX_v_6_2_2((z_out_40[16:11]),
          (z_out_45[16:11]), return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_nor_cse
        & (fsm_output[14]) ) begin
      return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_2_if_acc_1_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_nor_cse
        & (fsm_output[10]) ) begin
      return_mult_generic_AC_RND_CONV_false_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_if_acc_1_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_nor_cse
        & (fsm_output[12]) ) begin
      return_mult_generic_AC_RND_CONV_false_1_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_1_if_acc_1_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_r_inf_lpi_3_dfm_2
        | and_dcpl_166 | or_dcpl_187)) & (fsm_output[6]) ) begin
      return_add_generic_AC_RND_CONV_false_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & return_add_generic_AC_RND_CONV_false_acc_2_itm_11_1 & inverse_lpi_1_dfm_1
        & mode_lpi_1_dfm & (fsm_output[5]) ) begin
      return_add_generic_AC_RND_CONV_false_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_1_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_1_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_185 | (~ return_add_generic_AC_RND_CONV_false_1_acc_2_itm_11_1)))
        & (fsm_output[7]) ) begin
      return_add_generic_AC_RND_CONV_false_1_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_1_r_inf_lpi_3_dfm_2
        | and_dcpl_168 | or_dcpl_187)) & (fsm_output[8]) ) begin
      return_add_generic_AC_RND_CONV_false_1_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_207 | return_add_generic_AC_RND_CONV_false_2_r_inf_lpi_3_dfm_2
        | and_dcpl_166 | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva | or_dcpl_185))
        & (fsm_output[10]) ) begin
      return_add_generic_AC_RND_CONV_false_2_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_2_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_2_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_211) & (fsm_output[9]) ) begin
      return_add_generic_AC_RND_CONV_false_2_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_214 | return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
        | return_add_generic_AC_RND_CONV_false_3_r_inf_lpi_3_dfm_2 | or_dcpl_219))
        & (fsm_output[12]) ) begin
      return_add_generic_AC_RND_CONV_false_3_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_3_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_3_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_224) & (fsm_output[11]) ) begin
      return_add_generic_AC_RND_CONV_false_3_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_228 | or_dcpl_231 | return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
        | (~ mode_lpi_1_dfm))) & (fsm_output[14]) ) begin
      return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_234) & (fsm_output[13]) ) begin
      return_add_generic_AC_RND_CONV_false_6_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_237 | or_dcpl_240)) & (fsm_output[16]) ) begin
      return_add_generic_AC_RND_CONV_false_7_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_7_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_7_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_242) & (fsm_output[15]) ) begin
      return_add_generic_AC_RND_CONV_false_7_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_8_r_inf_lpi_3_dfm_2
        | or_dcpl_214 | or_dcpl_249)) & (fsm_output[18]) ) begin
      return_add_generic_AC_RND_CONV_false_8_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_8_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_8_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_252) & (fsm_output[17]) ) begin
      return_add_generic_AC_RND_CONV_false_8_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_nor_cse
        & (fsm_output[39]) ) begin
      return_mult_generic_AC_RND_CONV_false_5_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_5_if_acc_1_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_nor_cse
        & (fsm_output[35]) ) begin
      return_mult_generic_AC_RND_CONV_false_3_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_3_if_acc_1_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_return_mult_generic_AC_RND_CONV_false_2_do_shift_left_1_nor_cse
        & (fsm_output[37]) ) begin
      return_mult_generic_AC_RND_CONV_false_4_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_4_if_acc_1_itm_12_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_13_r_inf_lpi_3_dfm_2
        | or_dcpl_261 | and_dcpl_166 | or_dcpl_185)) & (fsm_output[31]) ) begin
      return_add_generic_AC_RND_CONV_false_13_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_13_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_13_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & return_add_generic_AC_RND_CONV_false_13_acc_2_itm_11_1 &
        inverse_lpi_1_dfm_1 & mode_lpi_1_dfm & (fsm_output[30]) ) begin
      return_add_generic_AC_RND_CONV_false_13_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_14_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_14_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & return_add_generic_AC_RND_CONV_false_14_acc_2_itm_11_1 &
        inverse_lpi_1_dfm_1 & mode_lpi_1_dfm & (fsm_output[32]) ) begin
      return_add_generic_AC_RND_CONV_false_14_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_14_r_inf_lpi_3_dfm_2
        | or_dcpl_261 | and_dcpl_168 | or_dcpl_185)) & (fsm_output[33]) ) begin
      return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_14_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_282 | return_add_generic_AC_RND_CONV_false_15_r_inf_lpi_3_dfm_2
        | and_dcpl_166 | return_add_generic_AC_RND_CONV_false_10_op1_inf_sva | or_dcpl_185))
        & (fsm_output[35]) ) begin
      return_add_generic_AC_RND_CONV_false_15_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_15_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_15_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_211) & (fsm_output[34]) ) begin
      return_add_generic_AC_RND_CONV_false_15_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_287 | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva
        | return_add_generic_AC_RND_CONV_false_16_r_inf_lpi_3_dfm_2 | or_dcpl_219))
        & (fsm_output[37]) ) begin
      return_add_generic_AC_RND_CONV_false_16_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_16_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_16_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_224) & (fsm_output[36]) ) begin
      return_add_generic_AC_RND_CONV_false_16_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_296 | or_dcpl_231 | return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
        | (~ mode_lpi_1_dfm))) & (fsm_output[39]) ) begin
      return_add_generic_AC_RND_CONV_false_19_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_234) & (fsm_output[38]) ) begin
      return_add_generic_AC_RND_CONV_false_19_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_302 | or_dcpl_240)) & (fsm_output[41]) ) begin
      return_add_generic_AC_RND_CONV_false_20_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_20_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_20_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_242) & (fsm_output[40]) ) begin
      return_add_generic_AC_RND_CONV_false_20_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_21_r_inf_lpi_3_dfm_2
        | or_dcpl_214 | or_dcpl_249)) & (fsm_output[43]) ) begin
      return_add_generic_AC_RND_CONV_false_21_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_21_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_21_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_252) & (fsm_output[42]) ) begin
      return_add_generic_AC_RND_CONV_false_21_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva <= 1'b0;
    end
    else if ( run_wen & and_dcpl_138 & and_dcpl_128 & (~ (operator_16_false_io_read_mode1_rsc_cse_sva[4]))
        & and_dcpl_152 & and_dcpl_151 & (~(operator_16_false_operator_16_false_nor_cse_sva
        | (z_out_27[11]))) & (fsm_output[54]) ) begin
      return_mult_generic_AC_RND_CONV_false_6_do_shift_left_1_sva <= return_mult_generic_AC_RND_CONV_false_6_if_acc_1_itm_11_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_9_r_inf_lpi_3_dfm_2
        | or_dcpl_201 | and_dcpl_166 | operator_11_true_return_1_sva | or_46_cse))
        & (fsm_output[20]) ) begin
      return_add_generic_AC_RND_CONV_false_9_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_9_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_9_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ return_add_generic_AC_RND_CONV_false_9_acc_2_itm_11_1)
        | inverse_lpi_1_dfm_1 | (~ mode_lpi_1_dfm))) & (fsm_output[19]) ) begin
      return_add_generic_AC_RND_CONV_false_9_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_10_r_inf_lpi_3_dfm_2
        | operator_11_true_return_15_sva | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
        | and_dcpl_166 | return_add_generic_AC_RND_CONV_false_10_op1_inf_sva | or_46_cse))
        & (fsm_output[22]) ) begin
      return_add_generic_AC_RND_CONV_false_10_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ return_add_generic_AC_RND_CONV_false_10_acc_2_itm_11_1)
        | inverse_lpi_1_dfm_1 | (~ mode_lpi_1_dfm))) & (fsm_output[21]) ) begin
      return_add_generic_AC_RND_CONV_false_10_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_207 | return_add_generic_AC_RND_CONV_false_11_r_inf_lpi_3_dfm_2
        | and_dcpl_166 | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva | or_46_cse))
        & (fsm_output[24]) ) begin
      return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ return_add_generic_AC_RND_CONV_false_11_acc_2_itm_11_1)
        | inverse_lpi_1_dfm_1 | (~ mode_lpi_1_dfm))) & (fsm_output[23]) ) begin
      return_add_generic_AC_RND_CONV_false_11_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_282 | return_add_generic_AC_RND_CONV_false_12_r_inf_lpi_3_dfm_2
        | and_dcpl_166 | return_add_generic_AC_RND_CONV_false_10_op1_inf_sva | or_46_cse))
        & (fsm_output[26]) ) begin
      return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ return_add_generic_AC_RND_CONV_false_12_acc_2_itm_11_1)
        | inverse_lpi_1_dfm_1 | (~ mode_lpi_1_dfm))) & (fsm_output[25]) ) begin
      return_add_generic_AC_RND_CONV_false_12_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_22_r_inf_lpi_3_dfm_2
        | operator_11_true_return_1_sva | return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
        | and_dcpl_166 | return_add_generic_AC_RND_CONV_false_22_op1_inf_sva | or_46_cse))
        & (fsm_output[45]) ) begin
      return_add_generic_AC_RND_CONV_false_22_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_22_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_22_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ return_add_generic_AC_RND_CONV_false_22_acc_2_itm_11_1)
        | inverse_lpi_1_dfm_1 | (~ mode_lpi_1_dfm))) & (fsm_output[44]) ) begin
      return_add_generic_AC_RND_CONV_false_22_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_23_r_inf_lpi_3_dfm_2
        | or_dcpl_201 | and_dcpl_166 | operator_11_true_return_15_sva | or_46_cse))
        & (fsm_output[47]) ) begin
      return_add_generic_AC_RND_CONV_false_23_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_6_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_23_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_23_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ return_add_generic_AC_RND_CONV_false_23_acc_2_itm_11_1)
        | inverse_lpi_1_dfm_1 | (~ mode_lpi_1_dfm))) & (fsm_output[46]) ) begin
      return_add_generic_AC_RND_CONV_false_23_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_282 | return_add_generic_AC_RND_CONV_false_24_r_inf_lpi_3_dfm_2
        | and_dcpl_166 | return_add_generic_AC_RND_CONV_false_22_op1_inf_sva | or_46_cse))
        & (fsm_output[49]) ) begin
      return_add_generic_AC_RND_CONV_false_24_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_12_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_24_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_24_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ return_add_generic_AC_RND_CONV_false_24_acc_2_itm_11_1)
        | inverse_lpi_1_dfm_1 | (~ mode_lpi_1_dfm))) & (fsm_output[48]) ) begin
      return_add_generic_AC_RND_CONV_false_24_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_207 | return_add_generic_AC_RND_CONV_false_25_r_inf_lpi_3_dfm_2
        | and_dcpl_166 | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva | or_46_cse))
        & (fsm_output[51]) ) begin
      return_add_generic_AC_RND_CONV_false_25_e_r_qelse_or_svs <= return_add_generic_AC_RND_CONV_false_11_e_r_qelse_or_svs_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_25_else_4_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_25_else_4_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~((~ return_add_generic_AC_RND_CONV_false_25_acc_2_itm_11_1)
        | inverse_lpi_1_dfm_1 | (~ mode_lpi_1_dfm))) & (fsm_output[50]) ) begin
      return_add_generic_AC_RND_CONV_false_25_else_4_unequal_tmp <= return_add_generic_AC_RND_CONV_false_1_else_4_return_add_generic_AC_RND_CONV_false_1_else_4_nand_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_16_false_io_read_mode1_rsc_cse_sva <= 16'b0000000000000000;
    end
    else if ( rst ) begin
      operator_16_false_io_read_mode1_rsc_cse_sva <= 16'b0000000000000000;
    end
    else if ( operator_16_false_and_cse & (~ operator_16_false_operator_16_false_nor_tmp)
        ) begin
      operator_16_false_io_read_mode1_rsc_cse_sva <= mode1_rsci_idat;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_16_false_operator_16_false_nor_cse_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_16_false_operator_16_false_nor_cse_sva <= 1'b0;
    end
    else if ( operator_16_false_and_cse ) begin
      operator_16_false_operator_16_false_nor_cse_sva <= operator_16_false_operator_16_false_nor_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      t_in_10_0_lpi_1_dfm_1_8 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_7 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_6 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_5 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_4 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_3 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_2 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_1 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_0 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_10 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_9 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_14 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_13 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_12 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_11 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_10 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_9 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_8 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_7 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_6 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_5 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_4 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_3 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_2 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_1 <= 1'b0;
      for_i_0_sva <= 1'b0;
    end
    else if ( rst ) begin
      t_in_10_0_lpi_1_dfm_1_8 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_7 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_6 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_5 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_4 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_3 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_2 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_1 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_0 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_10 <= 1'b0;
      t_in_10_0_lpi_1_dfm_1_9 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_14 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_13 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_12 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_11 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_10 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_9 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_8 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_7 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_6 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_5 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_4 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_3 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_2 <= 1'b0;
      m_in_15_1_lpi_1_dfm_1_1 <= 1'b0;
      for_i_0_sva <= 1'b0;
    end
    else if ( t_in_and_cse ) begin
      t_in_10_0_lpi_1_dfm_1_8 <= t_in_10_0_lpi_1_dfm_1_9 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_7 <= t_in_10_0_lpi_1_dfm_1_8 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_6 <= t_in_10_0_lpi_1_dfm_1_7 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_5 <= t_in_10_0_lpi_1_dfm_1_6 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_4 <= t_in_10_0_lpi_1_dfm_1_5 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_3 <= t_in_10_0_lpi_1_dfm_1_4 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_2 <= t_in_10_0_lpi_1_dfm_1_3 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_1 <= t_in_10_0_lpi_1_dfm_1_2 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_0 <= t_in_10_0_lpi_1_dfm_1_1 & (~ (fsm_output[1]));
      t_in_10_0_lpi_1_dfm_1_10 <= ~(operator_16_false_1_operator_16_false_1_and_mdf_sva_1
          | operator_16_false_operator_16_false_nor_tmp | or_dcpl_395);
      t_in_10_0_lpi_1_dfm_1_9 <= MUX_s_1_2_2(mode_lpi_1_dfm_mx0w0, t_in_10_0_lpi_1_dfm_1_10,
          or_dcpl_395);
      m_in_15_1_lpi_1_dfm_1_14 <= m_in_15_1_lpi_1_dfm_1_13 & or_dcpl_395;
      m_in_15_1_lpi_1_dfm_1_13 <= m_in_15_1_lpi_1_dfm_1_12 & or_dcpl_395;
      m_in_15_1_lpi_1_dfm_1_12 <= m_in_15_1_lpi_1_dfm_1_11 & or_dcpl_395;
      m_in_15_1_lpi_1_dfm_1_11 <= m_in_15_1_lpi_1_dfm_1_10 & or_dcpl_395;
      m_in_15_1_lpi_1_dfm_1_10 <= m_in_15_1_lpi_1_dfm_1_9 & or_dcpl_395;
      m_in_15_1_lpi_1_dfm_1_9 <= m_in_15_1_lpi_1_dfm_1_8 & or_dcpl_395;
      m_in_15_1_lpi_1_dfm_1_8 <= m_in_15_1_lpi_1_dfm_1_7 & or_dcpl_395;
      m_in_15_1_lpi_1_dfm_1_7 <= m_in_15_1_lpi_1_dfm_1_6 & or_dcpl_395;
      m_in_15_1_lpi_1_dfm_1_6 <= m_in_15_1_lpi_1_dfm_1_5 & or_dcpl_395;
      m_in_15_1_lpi_1_dfm_1_5 <= m_in_15_1_lpi_1_dfm_1_4 & or_dcpl_395;
      m_in_15_1_lpi_1_dfm_1_4 <= m_in_15_1_lpi_1_dfm_1_3 & or_dcpl_395;
      m_in_15_1_lpi_1_dfm_1_3 <= m_in_15_1_lpi_1_dfm_1_2 & or_dcpl_395;
      m_in_15_1_lpi_1_dfm_1_2 <= m_in_15_1_lpi_1_dfm_1_1 & or_dcpl_395;
      m_in_15_1_lpi_1_dfm_1_1 <= t_in_10_0_lpi_1_dfm_1_9 & or_dcpl_395;
      for_i_0_sva <= (~ for_i_0_sva) & or_dcpl_395;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      mode_lpi_1_dfm <= 1'b0;
      inverse_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( rst ) begin
      mode_lpi_1_dfm <= 1'b0;
      inverse_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( mode_and_cse ) begin
      mode_lpi_1_dfm <= mode_lpi_1_dfm_mx0w0;
      inverse_lpi_1_dfm_1 <= ~(((mode1_rsci_idat==16'b0000000000000010)) | operator_16_false_operator_16_false_nor_tmp);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_qr_1_10_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_qr_1_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_8 <= 1'b0;
      reg_stage_PE_1_qr_10_1_lpi_2_dfm_7_0_ftd <= 1'b0;
      reg_stage_PE_1_qr_10_1_lpi_2_dfm_7_0_ftd_1 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_qr_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_index_const_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_15_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_index_const_10_lpi_2_dfm <= 1'b0;
    end
    else if ( rst ) begin
      stage_PE_1_qr_1_10_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_qr_1_10_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_qr_1_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_8 <= 1'b0;
      reg_stage_PE_1_qr_10_1_lpi_2_dfm_7_0_ftd <= 1'b0;
      reg_stage_PE_1_qr_10_1_lpi_2_dfm_7_0_ftd_1 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_qr_10_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_qr_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_8 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_7 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_6 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_5 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_4 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_index_const_9_1_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_index_const_0_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_15_lpi_2_dfm <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_3 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_2 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_1 <= 1'b0;
      stage_PE_1_index_const_14_11_lpi_2_dfm_0 <= 1'b0;
      stage_PE_1_index_const_10_lpi_2_dfm <= 1'b0;
    end
    else if ( stage_PE_1_and_2_cse ) begin
      stage_PE_1_qr_1_10_1_lpi_2_dfm_8 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_8,
          t_in_10_0_lpi_1_dfm_1_9, t_in_10_0_lpi_1_dfm_1_8, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_7 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_7,
          t_in_10_0_lpi_1_dfm_1_8, t_in_10_0_lpi_1_dfm_1_7, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_6 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_6,
          t_in_10_0_lpi_1_dfm_1_7, t_in_10_0_lpi_1_dfm_1_6, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_5 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_5,
          t_in_10_0_lpi_1_dfm_1_6, t_in_10_0_lpi_1_dfm_1_5, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_4 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_4,
          t_in_10_0_lpi_1_dfm_1_5, t_in_10_0_lpi_1_dfm_1_4, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_3 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_3,
          t_in_10_0_lpi_1_dfm_1_4, t_in_10_0_lpi_1_dfm_1_3, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_2 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_2,
          t_in_10_0_lpi_1_dfm_1_3, t_in_10_0_lpi_1_dfm_1_2, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_1 <= MUX1HOT_s_1_3_2(m_in_15_1_lpi_1_dfm_1_1,
          t_in_10_0_lpi_1_dfm_1_2, t_in_10_0_lpi_1_dfm_1_1, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_10_1_lpi_2_dfm_0 <= MUX1HOT_s_1_3_2(t_in_10_0_lpi_1_dfm_1_9,
          t_in_10_0_lpi_1_dfm_1_1, t_in_10_0_lpi_1_dfm_1_0, {(~ inverse_lpi_1_dfm_1)
          , stage_PE_1_and_cse , stage_PE_1_and_1_tmp});
      stage_PE_1_qr_1_0_lpi_2_dfm <= t_in_10_0_lpi_1_dfm_1_10;
      stage_PE_1_qr_10_1_lpi_2_dfm_8 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_8,
          t_in_10_0_lpi_1_dfm_1_9, or_tmp_208);
      reg_stage_PE_1_qr_10_1_lpi_2_dfm_7_0_ftd <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_7,
          t_in_10_0_lpi_1_dfm_1_8, or_tmp_208);
      reg_stage_PE_1_qr_10_1_lpi_2_dfm_7_0_ftd_1 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_6,
          t_in_10_0_lpi_1_dfm_1_7, or_tmp_208);
      stage_PE_1_qr_10_1_lpi_2_dfm_5 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_5,
          t_in_10_0_lpi_1_dfm_1_6, or_tmp_208);
      stage_PE_1_qr_10_1_lpi_2_dfm_4 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_4,
          t_in_10_0_lpi_1_dfm_1_5, or_tmp_208);
      stage_PE_1_qr_10_1_lpi_2_dfm_3 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_3,
          t_in_10_0_lpi_1_dfm_1_4, or_tmp_208);
      stage_PE_1_qr_10_1_lpi_2_dfm_2 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_2,
          t_in_10_0_lpi_1_dfm_1_3, or_tmp_208);
      stage_PE_1_qr_10_1_lpi_2_dfm_1 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_1,
          t_in_10_0_lpi_1_dfm_1_2, or_tmp_208);
      stage_PE_1_qr_10_1_lpi_2_dfm_0 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_0,
          t_in_10_0_lpi_1_dfm_1_1, or_tmp_208);
      stage_PE_1_qr_0_lpi_2_dfm <= MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_9, t_in_10_0_lpi_1_dfm_1_10,
          stage_PE_qif_qelse_or_nl);
      stage_PE_1_index_const_9_1_lpi_2_dfm_8 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_8,
          t_in_10_0_lpi_1_dfm_1_10, or_tmp_208);
      stage_PE_1_index_const_9_1_lpi_2_dfm_7 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_7,
          t_in_10_0_lpi_1_dfm_1_9, or_tmp_208);
      stage_PE_1_index_const_9_1_lpi_2_dfm_6 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_6,
          t_in_10_0_lpi_1_dfm_1_8, or_tmp_208);
      stage_PE_1_index_const_9_1_lpi_2_dfm_5 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_5,
          t_in_10_0_lpi_1_dfm_1_7, or_tmp_208);
      stage_PE_1_index_const_9_1_lpi_2_dfm_4 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_4,
          t_in_10_0_lpi_1_dfm_1_6, or_tmp_208);
      stage_PE_1_index_const_9_1_lpi_2_dfm_3 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_3,
          t_in_10_0_lpi_1_dfm_1_5, or_tmp_208);
      stage_PE_1_index_const_9_1_lpi_2_dfm_2 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_2,
          t_in_10_0_lpi_1_dfm_1_4, or_tmp_208);
      stage_PE_1_index_const_9_1_lpi_2_dfm_1 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_1,
          t_in_10_0_lpi_1_dfm_1_3, or_tmp_208);
      stage_PE_1_index_const_9_1_lpi_2_dfm_0 <= MUX_s_1_2_2(stage_PE_qif_qr_15_1_lpi_2_dfm_mx0_0,
          t_in_10_0_lpi_1_dfm_1_2, or_tmp_208);
      stage_PE_1_index_const_0_lpi_2_dfm <= MUX_s_1_2_2(stage_PE_qif_qelse_mux_nl,
          t_in_10_0_lpi_1_dfm_1_1, or_tmp_208);
      stage_PE_1_index_const_15_lpi_2_dfm <= m_in_15_1_lpi_1_dfm_1_14 & (~ mode_lpi_1_dfm)
          & inverse_lpi_1_dfm_1;
      stage_PE_1_index_const_14_11_lpi_2_dfm_3 <= stage_PE_qif_qelse_mux_1_nl & inverse_lpi_1_dfm_1;
      stage_PE_1_index_const_14_11_lpi_2_dfm_2 <= stage_PE_qif_qelse_mux_14_nl &
          inverse_lpi_1_dfm_1;
      stage_PE_1_index_const_14_11_lpi_2_dfm_1 <= stage_PE_qif_qelse_mux_13_nl &
          inverse_lpi_1_dfm_1;
      stage_PE_1_index_const_14_11_lpi_2_dfm_0 <= stage_PE_qif_qelse_mux_12_nl &
          inverse_lpi_1_dfm_1;
      stage_PE_1_index_const_10_lpi_2_dfm <= stage_PE_qif_qelse_mux_11_nl & inverse_lpi_1_dfm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_fry_9_0_sva <= 10'b0000000000;
    end
    else if ( rst ) begin
      BUTTERFLY_1_fry_9_0_sva <= 10'b0000000000;
    end
    else if ( run_wen & (~(and_dcpl_233 & (~((fsm_output[0]) | (fsm_output[2]) |
        (fsm_output[28]))) & (~((fsm_output[3]) | (fsm_output[50]) | (fsm_output[25])))))
        ) begin
      BUTTERFLY_1_fry_9_0_sva <= MUX_v_10_2_2(10'b0000000000, BUTTERFLY_fry_BUTTERFLY_fry_mux_nl,
          not_709_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_26_m_zero_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_26_m_zero_sva <= 1'b0;
    end
    else if ( run_wen & ((~(inverse_lpi_1_dfm_1 | (and_dcpl_214 & and_dcpl_211 &
        and_dcpl_236 & (~((fsm_output[31]) | (fsm_output[6])))))) | (fsm_output[2]))
        ) begin
      return_extract_26_m_zero_sva <= MUX1HOT_s_1_3_2(stage_PE_1_and_1_tmp, return_extract_3_m_zero_sva_mx1w0,
          return_extract_26_m_zero_sva_2, {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[31])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_15_return_extract_15_nor_cse_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_15_return_extract_15_nor_cse_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm <= 1'b0;
    end
    else if ( return_extract_15_and_3_cse ) begin
      return_extract_15_return_extract_15_nor_cse_sva <= MUX1HOT_s_1_6_2(return_extract_15_return_extract_15_nor_nl,
          return_extract_15_return_extract_15_nor_cse_sva_mx1, stage_d_mul_return_d_2_63_sva_1,
          return_extract_47_return_extract_47_nor_nl, return_extract_15_return_extract_15_nor_cse_sva_mx2,
          stage_d_mul_return_d_5_63_sva_1, {(fsm_output[3]) , (fsm_output[10]) ,
          (fsm_output[12]) , (fsm_output[28]) , (fsm_output[35]) , (fsm_output[37])});
      return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm <= MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1,
          (stage_PE_1_tmp_re_d_1_sva_1_63_57[6]), return_add_generic_AC_RND_CONV_false_11_mux_itm,
          stage_d_mul_return_d_4_63_sva_1, return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm_1,
          stage_d_mul_return_d_63_sva_1, {(fsm_output[3]) , return_add_generic_AC_RND_CONV_false_17_e_r_and_cse
          , return_add_generic_AC_RND_CONV_false_17_e_r_and_1_nl , (fsm_output[12])
          , (fsm_output[28]) , (fsm_output[37])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_15_m_zero_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_15_m_zero_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_449 | or_dcpl_447 | or_dcpl_445 | or_dcpl_421
        | or_dcpl_163 | (fsm_output[12]) | or_dcpl_440 | or_dcpl_438 | or_dcpl_95))
        ) begin
      return_extract_15_m_zero_sva <= MUX1HOT_s_1_5_2(return_extract_15_m_zero_mux1h_cse,
          return_extract_20_m_zero_return_extract_20_m_zero_nor_nl, return_extract_25_m_zero_return_extract_25_m_zero_nor_nl,
          return_extract_26_m_zero_sva_2, return_extract_54_m_zero_return_extract_54_m_zero_nor_nl,
          {(fsm_output[3]) , (fsm_output[10]) , (fsm_output[16]) , or_tmp_261 , (fsm_output[37])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_15_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_15_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_466 | or_dcpl_464 | or_dcpl_462 | or_dcpl_136
        | (fsm_output[9]) | (fsm_output[37]) | (fsm_output[12]) | or_dcpl_418 | (fsm_output[19])
        | (fsm_output[6]) | (fsm_output[5]) | or_dcpl_415)) ) begin
      operator_11_true_return_15_sva <= MUX1HOT_s_1_8_2(operator_11_true_15_operator_11_true_15_and_nl,
          return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_tmp,
          operator_11_true_21_operator_11_true_21_and_nl, operator_11_true_27_operator_11_true_27_and_nl,
          operator_11_true_33_operator_11_true_33_and_tmp, return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp,
          operator_11_true_53_operator_11_true_53_and_nl, operator_11_true_59_operator_11_true_59_and_nl,
          {(fsm_output[3]) , (fsm_output[10]) , (fsm_output[14]) , (fsm_output[18])
          , or_1375_cse , (fsm_output[35]) , (fsm_output[39]) , (fsm_output[43])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_11_op_bigger_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm <= MUX1HOT_s_1_13_2(return_add_generic_AC_RND_CONV_false_17_op2_mu_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_17_op1_mu_0_lpi_3_dfm_1, drf_qr_lval_13_smx_0_lpi_3_dfm,
          return_add_generic_AC_RND_CONV_false_op2_mu_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_3_nl,
          return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_6_cse,
          return_add_generic_AC_RND_CONV_false_13_op1_mu_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_3_nl,
          return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_12_cse,
          return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[50]),
          {return_add_generic_AC_RND_CONV_false_11_op_bigger_and_5_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_6_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_5_nl , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse
          , (fsm_output[10]) , (fsm_output[14]) , (fsm_output[16]) , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_7_cse
          , (fsm_output[35]) , (fsm_output[39]) , (fsm_output[41]) , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_16_cse});
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm <= MUX1HOT_s_1_15_2(stage_PE_1_gm_im_d_mux_cse,
          return_add_generic_AC_RND_CONV_false_17_op1_mu_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1,
          (return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1[50]), return_add_generic_AC_RND_CONV_false_11_mux_2_itm_mx3,
          return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_21_cse,
          return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1, (return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1[50]),
          drf_qr_lval_14_smx_0_lpi_3_dfm_mx3, return_add_generic_AC_RND_CONV_false_20_op2_mu_1_51_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_27_cse, return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1,
          {return_add_generic_AC_RND_CONV_false_11_op_bigger_and_5_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_6_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_8_nl , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_6_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_10_nl , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_23_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_24_cse , (fsm_output[14])
          , (fsm_output[16]) , return_add_generic_AC_RND_CONV_false_11_op_bigger_or_7_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_29_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_30_cse
          , (fsm_output[39]) , (fsm_output[41]) , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_15_e_dif_sat_sva <= 6'b000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_15_e_dif_sat_sva <= 6'b000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_11_op_smaller_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm <= MUX1HOT_s_1_11_2(return_add_generic_AC_RND_CONV_false_4_op_smaller_qr_0_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx1,
          return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx2,
          return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_2_cse, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx5,
          return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_0_lpi_3_dfm_mx6,
          return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_20_op2_mu_1_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_3_cse, {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
          , (fsm_output[5]) , (fsm_output[7]) , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_4_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse , (fsm_output[16])
          , (fsm_output[30]) , (fsm_output[32]) , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_cse , (fsm_output[41])});
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_51_lpi_3_dfm <= MUX1HOT_s_1_9_2(return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_6_cse,
          return_add_generic_AC_RND_CONV_false_op2_mu_52_lpi_3_dfm_1, drf_qr_lval_13_smx_0_lpi_3_dfm,
          return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm, return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_cse, return_add_generic_AC_RND_CONV_false_13_op1_mu_52_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_20_op2_mu_1_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_5_op_smaller_mux_cse,
          {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_or_nl
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_or_5_nl , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_4_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse , (fsm_output[16])
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_or_6_nl , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_cse
          , (fsm_output[41])});
      return_add_generic_AC_RND_CONV_false_15_e_dif_sat_sva <= MUX1HOT_v_6_6_2(return_add_generic_AC_RND_CONV_false_4_e_dif_sat_sva_1,
          return_add_generic_AC_RND_CONV_false_2_e_dif_sat_sva_1, return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_cse,
          return_add_generic_AC_RND_CONV_false_8_e_dif_sat_or_cse, return_add_generic_AC_RND_CONV_false_11_e_dif_sat_or_nl,
          return_add_generic_AC_RND_CONV_false_21_e_dif_sat_or_cse, {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
          , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse
          , (fsm_output[14]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse
          , (fsm_output[39])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & ((~(return_add_generic_AC_RND_CONV_false_8_op1_smaller_return_add_generic_AC_RND_CONV_false_8_op1_smaller_or_cse
        | or_dcpl_488 | or_dcpl_503 | (fsm_output[33]) | or_dcpl_502 | or_dcpl_418
        | (fsm_output[18]) | (fsm_output[17]) | (fsm_output[31]) | or_dcpl_495))
        | (fsm_output[3]) | (fsm_output[10]) | (fsm_output[12]) | (fsm_output[16])
        | (fsm_output[28]) | (fsm_output[35]) | (fsm_output[39]) | (fsm_output[41]))
        ) begin
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm <= MUX1HOT_s_1_12_2(return_extract_15_return_extract_15_or_1_nl,
          return_extract_15_return_extract_15_nor_cse_sva_mx1, stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx1_50,
          return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_2_nl,
          return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_22_op1_mu_mux_cse,
          return_extract_47_return_extract_47_or_1_nl, return_extract_44_return_extract_44_or_1_cse_sva_1,
          return_extract_15_return_extract_15_nor_cse_sva_mx2, return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm,
          return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_22_op1_mu_mux_1_cse,
          {(fsm_output[3]) , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_12_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_13_cse , (fsm_output[12])
          , (fsm_output[14]) , (fsm_output[16]) , (fsm_output[28]) , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_14_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_15_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_cse , (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm <= 1'b0;
    end
    else if ( rst ) begin
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm <= 1'b0;
    end
    else if ( run_wen & ((inverse_lpi_1_dfm_1 & (~(or_dcpl_102 | (fsm_output[10])
        | or_dcpl_519 | or_dcpl_518 | or_dcpl_514 | or_dcpl_513 | or_dcpl_512)))
        | return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse | (fsm_output[16])
        | or_tmp_234 | or_dcpl_397 | (fsm_output[41])) ) begin
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm <= MUX1HOT_s_1_5_2(return_extract_9_return_extract_9_or_1_cse_sva_1,
          BUTTERFLY_1_fiy_mux1h_2_cse, (BUTTERFLY_1_fry_9_0_sva[9]), (BUTTERFLY_1_i_9_0_sva[9]),
          BUTTERFLY_1_fiy_mux1h_6_cse, {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
          , (fsm_output[16]) , BUTTERFLY_1_fiy_or_1_cse , or_tmp_234 , (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_14_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      drf_qr_lval_14_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & ((~(and_dcpl_233 & and_dcpl_286 & and_dcpl_284 & (~ (fsm_output[50]))
        & (~((fsm_output[49]) | (fsm_output[25]))) & (~((fsm_output[40]) | (fsm_output[15])))
        & (~((fsm_output[24]) | (fsm_output[39]))) & (~((fsm_output[10]) | (fsm_output[14])))
        & (~ (fsm_output[11])))) | (fsm_output[12]) | (fsm_output[16]) | (fsm_output[35])
        | (fsm_output[41])) ) begin
      drf_qr_lval_14_smx_0_lpi_3_dfm <= MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_4_m_r_51_lpi_3_dfm_1,
          drf_qr_lval_14_smx_0_lpi_3_dfm_mx1, BUTTERFLY_1_fiy_mux1h_2_cse, drf_qr_lval_14_smx_0_lpi_3_dfm_mx3,
          BUTTERFLY_1_fiy_mux1h_6_cse, {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
          , (fsm_output[12]) , (fsm_output[16]) , (fsm_output[35]) , (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_i_9_0_sva <= 10'b0000000000;
    end
    else if ( rst ) begin
      BUTTERFLY_1_i_9_0_sva <= 10'b0000000000;
    end
    else if ( run_wen & (~(nor_24_cse & (~ (fsm_output[51])) & (~((fsm_output[26])
        | (fsm_output[1]) | (fsm_output[55]))) & and_dcpl_165 & (~ (fsm_output[53]))
        & (~((fsm_output[54]) | (fsm_output[23]) | (fsm_output[48]))) & (~((fsm_output[2])
        | (fsm_output[28]) | (fsm_output[3]))) & (~((fsm_output[47]) | (fsm_output[50])
        | (fsm_output[46]))) & (~((fsm_output[49]) | (fsm_output[22]) | (fsm_output[25])))
        & (~((fsm_output[24]) | (fsm_output[21]))))) ) begin
      BUTTERFLY_1_i_9_0_sva <= BUTTERFLY_i_9_0_sva_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_n_9_0_sva_1 <= 10'b0000000000;
    end
    else if ( rst ) begin
      BUTTERFLY_1_n_9_0_sva_1 <= 10'b0000000000;
    end
    else if ( BUTTERFLY_1_n_and_cse & (~(BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_tmp
        & mode_lpi_1_dfm)) ) begin
      BUTTERFLY_1_n_9_0_sva_1 <= z_out_19[9:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_13_smx_10_1_lpi_3_dfm <= 10'b0000000000;
    end
    else if ( rst ) begin
      drf_qr_lval_13_smx_10_1_lpi_3_dfm <= 10'b0000000000;
    end
    else if ( run_wen & (~(or_dcpl_102 | (fsm_output[42]) | or_dcpl_125 | or_dcpl_542
        | or_dcpl_163 | (fsm_output[19]) | or_dcpl_401 | or_dcpl_417)) ) begin
      drf_qr_lval_13_smx_10_1_lpi_3_dfm <= MUX1HOT_v_10_6_2(return_add_generic_AC_RND_CONV_false_4_e_r_qelse_qr_10_1_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1, (stage_PE_1_x_im_d_sva[62:53]),
          return_add_generic_AC_RND_CONV_false_17_e_r_qelse_qr_10_1_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1, (stage_PE_1_x_re_d_sva[62:53]),
          {(fsm_output[3]) , return_add_generic_AC_RND_CONV_false_10_exp_and_2_cse
          , return_add_generic_AC_RND_CONV_false_10_exp_and_3_cse , (fsm_output[28])
          , return_add_generic_AC_RND_CONV_false_10_exp_and_4_cse , return_add_generic_AC_RND_CONV_false_10_exp_and_5_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm <= 1'b0;
    end
    else if ( rst ) begin
      BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm <= 1'b0;
    end
    else if ( BUTTERFLY_1_n_and_cse & mode_lpi_1_dfm ) begin
      BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_itm <= BUTTERFLY_1_if_3_BUTTERFLY_1_if_3_if_1_and_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_17_mux_6_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_17_mux_6_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_108 | or_dcpl_106 | or_dcpl_561 | or_dcpl_558
        | or_dcpl_556 | or_dcpl_553 | or_dcpl_551 | or_dcpl_512)) ) begin
      return_add_generic_AC_RND_CONV_false_17_mux_6_itm <= MUX1HOT_s_1_9_2(return_add_generic_AC_RND_CONV_false_17_if_2_return_add_generic_AC_RND_CONV_false_17_if_2_nor_1_nl,
          (O_1_out[63]), (~ inverse_lpi_1_dfm_1), return_add_generic_AC_RND_CONV_false_9_if_2_return_add_generic_AC_RND_CONV_false_9_if_2_and_1_mx2w0,
          (stage_PE_1_x_re_d_sva[63]), return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_12_if_2_return_add_generic_AC_RND_CONV_false_12_if_2_nor_mx4w0,
          (stage_PE_1_x_im_d_sva[63]), (~ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva),
          {return_add_generic_AC_RND_CONV_false_17_and_1_nl , return_add_generic_AC_RND_CONV_false_17_and_7_nl
          , return_add_generic_AC_RND_CONV_false_17_and_8_nl , return_add_generic_AC_RND_CONV_false_17_and_3_cse
          , return_add_generic_AC_RND_CONV_false_17_and_9_cse , return_add_generic_AC_RND_CONV_false_17_and_10_cse
          , return_add_generic_AC_RND_CONV_false_17_and_5_cse , return_add_generic_AC_RND_CONV_false_17_and_11_cse
          , return_add_generic_AC_RND_CONV_false_17_and_12_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_571 | or_dcpl_420)) & mode_lpi_1_dfm ) begin
      return_add_generic_AC_RND_CONV_false_18_mux_itm <= MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_18_if_2_return_add_generic_AC_RND_CONV_false_18_if_2_and_2_nl,
          return_add_generic_AC_RND_CONV_false_18_r_sign_mux_1_nl, or_dcpl_549);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_do_sub_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_do_sub_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_465 | (fsm_output[45]) | (fsm_output[40]) | or_dcpl_580
        | or_dcpl_579 | or_dcpl_576 | or_dcpl_575 | or_dcpl_574)) ) begin
      return_add_generic_AC_RND_CONV_false_10_do_sub_sva <= MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_5_do_sub_return_add_generic_AC_RND_CONV_false_5_do_sub_xor_nl,
          return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_tmp,
          return_add_generic_AC_RND_CONV_false_10_do_sub_return_add_generic_AC_RND_CONV_false_10_do_sub_xor_nl,
          return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp,
          return_add_generic_AC_RND_CONV_false_23_do_sub_return_add_generic_AC_RND_CONV_false_23_do_sub_xor_nl,
          {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , (fsm_output[12])
          , (fsm_output[14]) , (fsm_output[37]) , (fsm_output[39])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
        | (fsm_output[10]) | or_dcpl_519 | or_dcpl_502 | or_dcpl_587 | (fsm_output[12])
        | or_dcpl_586 | or_dcpl_495)) ) begin
      return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1 <= MUX1HOT_s_1_3_2(return_extract_18_and_nl,
          return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1, return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2,
          {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , (fsm_output[14])
          , (fsm_output[39])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & ((reg_return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_rgt_nl
        & (~(or_dcpl_610 | or_dcpl_607 | or_dcpl_99 | or_dcpl_159 | (fsm_output[35])
        | or_dcpl_404 | or_dcpl_418 | or_dcpl_573))) | (fsm_output[3]) | (fsm_output[4])
        | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[28]) | (fsm_output[29]))
        & ((~ and_dcpl_258) | return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
        | return_add_generic_AC_RND_CONV_false_13_op2_mu_or_3_rgt | or_1375_cse |
        return_add_generic_AC_RND_CONV_false_13_op2_mu_or_8_rgt | return_add_generic_AC_RND_CONV_false_13_op2_mu_or_9_rgt)
        ) begin
      return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm <= MUX1HOT_v_51_5_2(return_add_generic_AC_RND_CONV_false_17_op_bigger_mux_8_cse,
          return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx1, return_extract_32_mux_4_cse,
          (in_f_d_rsci_q_d[51:1]), (in_f_d_rsci_q_d[50:0]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
          , return_add_generic_AC_RND_CONV_false_13_op2_mu_or_10_nl , or_1375_cse
          , return_add_generic_AC_RND_CONV_false_13_op2_mu_or_8_rgt , return_add_generic_AC_RND_CONV_false_13_op2_mu_or_9_rgt});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_gm_im_d_61_0_lpi_3_dfm <= 62'b00000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      stage_PE_1_gm_im_d_61_0_lpi_3_dfm <= 62'b00000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_407 | or_dcpl_99 | or_dcpl_631 | or_dcpl_514 |
        or_dcpl_628 | or_dcpl_495)) & mode_lpi_1_dfm ) begin
      stage_PE_1_gm_im_d_61_0_lpi_3_dfm <= O_1_out_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_else_3_else_acc_4_itm_15_14 <= 2'b00;
    end
    else if ( rst ) begin
      BUTTERFLY_1_else_3_else_acc_4_itm_15_14 <= 2'b00;
    end
    else if ( BUTTERFLY_1_else_3_else_and_ssc ) begin
      BUTTERFLY_1_else_3_else_acc_4_itm_15_14 <= MUX_v_2_2_2((z_out_4_31_16[15:14]),
          (z_out_38[15:14]), return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_1_m_zero_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_1_m_zero_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_466 | return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
        | or_dcpl_444 | or_dcpl_99 | return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse
        | (fsm_output[35]) | (fsm_output[36]) | (fsm_output[17]) | or_dcpl_666 |
        return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse)) ) begin
      return_extract_1_m_zero_sva <= MUX1HOT_s_1_5_2(return_extract_3_m_zero_sva_mx1w0,
          return_extract_22_m_zero_return_extract_22_m_zero_nor_nl, return_extract_15_m_zero_mux1h_cse,
          return_extract_53_m_zero_return_extract_53_m_zero_nor_nl, return_extract_59_m_zero_return_extract_59_m_zero_nor_nl,
          {or_tmp_440 , (fsm_output[12]) , (fsm_output[29]) , (fsm_output[39]) ,
          (fsm_output[43])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_1_sva <= 1'b0;
    end
    else if ( run_wen & (~((fsm_output[50]) | (fsm_output[49]) | (fsm_output[44])
        | (fsm_output[25]) | (fsm_output[40]) | (fsm_output[15]) | (fsm_output[24])
        | (fsm_output[43]) | (fsm_output[42]) | or_dcpl_682 | (fsm_output[14]) |
        (fsm_output[38]) | (fsm_output[32]) | (fsm_output[7]) | or_dcpl_514 | or_dcpl_513
        | (fsm_output[17]) | (fsm_output[5]))) ) begin
      operator_11_true_return_1_sva <= MUX1HOT_s_1_8_2(operator_11_true_24_operator_11_true_24_and_tmp,
          operator_11_true_20_operator_11_true_20_and_nl, operator_11_true_25_operator_11_true_25_and_nl,
          return_add_generic_AC_RND_CONV_false_12_r_nan_and_nl, operator_11_true_33_operator_11_true_33_and_tmp,
          operator_11_true_52_operator_11_true_52_and_nl, operator_11_true_57_operator_11_true_57_and_nl,
          return_add_generic_AC_RND_CONV_false_25_r_nan_and_nl, {or_tmp_440 , (fsm_output[10])
          , (fsm_output[16]) , (fsm_output[23]) , or_tmp_261 , (fsm_output[35]) ,
          (fsm_output[41]) , (fsm_output[48])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_17_return_extract_17_nor_cse_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_17_return_extract_17_nor_cse_sva <= 1'b0;
    end
    else if ( return_extract_17_and_3_cse & mode_lpi_1_dfm ) begin
      return_extract_17_return_extract_17_nor_cse_sva <= ~((return_add_generic_AC_RND_CONV_false_5_e_r_qelse_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
          | return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_17_m_zero_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_17_m_zero_sva <= 1'b0;
    end
    else if ( run_wen & ((return_extract_17_m_zero_mux_nl & (~(or_dcpl_464 | or_dcpl_707
        | or_dcpl_705 | or_dcpl_704 | or_dcpl_517 | or_dcpl_597 | or_dcpl_440 | (fsm_output[31])
        | or_dcpl_493))) | (fsm_output[4]) | (fsm_output[14]) | (fsm_output[18])
        | (fsm_output[29])) ) begin
      return_extract_17_m_zero_sva <= MUX1HOT_s_1_4_2(return_extract_15_m_zero_mux1h_cse,
          return_extract_21_m_zero_return_extract_21_m_zero_nor_nl, return_extract_27_m_zero_return_extract_27_m_zero_nor_nl,
          return_extract_26_m_zero_sva_2, {(fsm_output[4]) , (fsm_output[14]) , (fsm_output[18])
          , return_extract_17_m_zero_or_2_nl});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_17_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_17_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_719 | or_dcpl_445 | or_dcpl_716 | or_dcpl_697
        | or_dcpl_713 | or_dcpl_511 | or_dcpl_118)) ) begin
      operator_11_true_return_17_sva <= MUX1HOT_s_1_4_2(operator_11_true_return_17_sva_mx0w0,
          operator_11_true_22_operator_11_true_22_and_nl, operator_11_true_47_operator_11_true_47_and_nl,
          operator_11_true_54_operator_11_true_54_and_nl, {(fsm_output[4]) , (fsm_output[12])
          , (fsm_output[28]) , (fsm_output[37])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & (~((fsm_output[44]) | (fsm_output[10]) | or_dcpl_99 | or_dcpl_422
        | or_dcpl_694 | or_dcpl_440 | or_dcpl_722)) ) begin
      return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm <= MUX1HOT_s_1_7_2(return_extract_17_return_extract_17_or_1_nl,
          return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm_mx1,
          return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_2_cse, return_add_generic_AC_RND_CONV_false_1_op_bigger_mux_4_cse,
          return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm_mx4,
          return_add_generic_AC_RND_CONV_false_9_op_bigger_mux_3_cse, return_add_generic_AC_RND_CONV_false_1_op_bigger_mux_5_cse,
          {or_38_cse , (fsm_output[14]) , (fsm_output[16]) , (fsm_output[18]) , (fsm_output[39])
          , (fsm_output[41]) , (fsm_output[43])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_13_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      drf_qr_lval_13_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_466 | (fsm_output[15]) | (fsm_output[20]) | or_dcpl_406
        | or_dcpl_736 | (fsm_output[38]) | (fsm_output[8]) | (fsm_output[7]) | (fsm_output[9])
        | (fsm_output[12]) | or_dcpl_440 | or_dcpl_573)) ) begin
      drf_qr_lval_13_smx_0_lpi_3_dfm <= MUX1HOT_s_1_7_2(return_add_generic_AC_RND_CONV_false_op2_mu_52_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_10_exp_mux1h_8_cse, return_add_generic_AC_RND_CONV_false_13_op1_mu_52_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm_mx0w4, (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[50]),
          return_add_generic_AC_RND_CONV_false_11_mux_2_itm_mx9, return_add_generic_AC_RND_CONV_false_10_exp_mux1h_11_cse,
          {or_tmp_440 , (fsm_output[18]) , or_1586_nl , (fsm_output[36]) , return_add_generic_AC_RND_CONV_false_10_exp_and_6_cse
          , return_add_generic_AC_RND_CONV_false_10_exp_and_7_cse , (fsm_output[43])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_15_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      drf_qr_lval_15_smx_0_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_661 | (fsm_output[47]) | (fsm_output[50]) | or_dcpl_534
        | (fsm_output[44]) | or_dcpl_751 | or_dcpl_126 | or_dcpl_750 | or_dcpl_542
        | or_dcpl_517 | or_dcpl_418 | (fsm_output[19]) | (fsm_output[31]) | or_dcpl_693))
        ) begin
      drf_qr_lval_15_smx_0_lpi_3_dfm <= MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_4_m_r_51_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_10_exp_mux1h_8_cse, return_add_generic_AC_RND_CONV_false_10_exp_mux1h_11_cse,
          {or_38_cse , (fsm_output[18]) , (fsm_output[43])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_14_smx_10_1_lpi_3_dfm <= 10'b0000000000;
    end
    else if ( rst ) begin
      drf_qr_lval_14_smx_10_1_lpi_3_dfm <= 10'b0000000000;
    end
    else if ( run_wen & (~(or_dcpl_769 | (fsm_output[44]) | or_dcpl_751 | (fsm_output[20])
        | (fsm_output[10]) | (fsm_output[21]) | (fsm_output[33]) | or_dcpl_501 |
        or_dcpl_517 | or_dcpl_418 | (fsm_output[19]) | or_dcpl_133 | (fsm_output[31])
        | or_dcpl_693)) ) begin
      drf_qr_lval_14_smx_10_1_lpi_3_dfm <= MUX1HOT_v_10_5_2(return_add_generic_AC_RND_CONV_false_5_e_r_qelse_qr_10_1_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1, (stage_PE_1_x_re_d_sva[62:53]),
          return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1, (stage_PE_1_x_im_d_sva[62:53]),
          {or_38_cse , return_add_generic_AC_RND_CONV_false_11_exp_and_2_cse , return_add_generic_AC_RND_CONV_false_11_exp_and_3_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_16_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_18_e_r_qr_0_lpi_3_dfm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_18_e_r_qr_0_lpi_3_dfm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_406 | or_dcpl_776 | or_dcpl_500 | or_dcpl_136
        | or_dcpl_553 | or_dcpl_722)) ) begin
      return_add_generic_AC_RND_CONV_false_18_e_r_qr_0_lpi_3_dfm <= MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1,
          stage_d_mul_return_d_63_sva_1, stage_d_mul_return_d_4_63_sva_1, {or_38_cse
          , (fsm_output[12]) , (fsm_output[37])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( return_extract_17_and_3_cse ) begin
      return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm <= return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_extract_24_m_zero_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_extract_24_m_zero_sva <= 1'b0;
    end
    else if ( run_wen & ((inverse_lpi_1_dfm_1 & (~(or_dcpl_803 | or_dcpl_788 | (fsm_output[39])
        | or_dcpl_799 | or_dcpl_776 | (fsm_output[34]) | or_dcpl_421 | (fsm_output[9])
        | or_dcpl_514 | or_dcpl_793 | or_dcpl_118))) | (fsm_output[5]) | (fsm_output[28])
        | (fsm_output[35]) | (fsm_output[41])) ) begin
      return_extract_24_m_zero_sva <= MUX1HOT_s_1_4_2(return_extract_3_m_zero_sva_mx1w0,
          return_extract_15_m_zero_mux1h_cse, return_extract_52_m_zero_return_extract_52_m_zero_nor_nl,
          return_extract_57_m_zero_return_extract_57_m_zero_nor_nl, {or_219_cse ,
          (fsm_output[28]) , (fsm_output[35]) , (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_24_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_24_sva <= 1'b0;
    end
    else if ( run_wen & ((inverse_lpi_1_dfm_1 & (~(or_dcpl_662 | or_dcpl_751 | (fsm_output[25])
        | (fsm_output[15]) | (fsm_output[24]) | or_dcpl_406 | or_dcpl_736 | (fsm_output[33])
        | or_dcpl_500 | or_dcpl_159 | (fsm_output[35]) | (fsm_output[12]) | (fsm_output[36])
        | or_dcpl_513 | or_dcpl_401 | (fsm_output[30])))) | (fsm_output[5]) | (fsm_output[17])
        | (fsm_output[20]) | (fsm_output[29]) | (fsm_output[44])) ) begin
      operator_11_true_return_24_sva <= MUX1HOT_s_1_3_2(operator_11_true_24_operator_11_true_24_and_tmp,
          all_same_out, operator_11_true_return_17_sva_mx0w0, {or_219_cse , return_extract_1_exception_or_cse
          , (fsm_output[29])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_mux_2_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_mux_2_itm <= 1'b0;
    end
    else if ( run_wen & (~((fsm_output[43]) | (fsm_output[13]) | (fsm_output[38])
        | or_dcpl_618 | (fsm_output[18]))) ) begin
      return_add_generic_AC_RND_CONV_false_11_mux_2_itm <= MUX1HOT_s_1_22_2((~ return_add_generic_AC_RND_CONV_false_2_res_mant_3_0_sva_1),
          return_add_generic_AC_RND_CONV_false_2_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_3_res_mant_3_0_sva_1),
          return_add_generic_AC_RND_CONV_false_3_res_mant_3_0_sva_1, return_add_generic_AC_RND_CONV_false_11_mux_2_itm_mx3,
          return_add_generic_AC_RND_CONV_false_7_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_7_res_mant_3_0_sva_1),
          return_add_generic_AC_RND_CONV_false_9_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_9_res_mant_3_0_sva_1),
          return_add_generic_AC_RND_CONV_false_11_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_11_res_mant_3_0_sva_1),
          (~ return_add_generic_AC_RND_CONV_false_15_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_15_res_mant_3_0_sva_1,
          (~ return_add_generic_AC_RND_CONV_false_16_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_16_res_mant_3_0_sva_1,
          return_add_generic_AC_RND_CONV_false_11_mux_2_itm_mx9, return_add_generic_AC_RND_CONV_false_20_res_mant_3_0_sva_1,
          (~ return_add_generic_AC_RND_CONV_false_20_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_22_res_mant_3_0_sva_1,
          (~ return_add_generic_AC_RND_CONV_false_22_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_8_res_mant_3_0_sva_1,
          (~ return_add_generic_AC_RND_CONV_false_8_res_mant_3_0_sva_1), {return_add_generic_AC_RND_CONV_false_11_and_3_cse
          , return_add_generic_AC_RND_CONV_false_11_and_4_cse , return_add_generic_AC_RND_CONV_false_11_and_5_cse
          , return_add_generic_AC_RND_CONV_false_11_and_6_cse , (fsm_output[10])
          , return_add_generic_AC_RND_CONV_false_11_and_7_nl , return_add_generic_AC_RND_CONV_false_11_and_8_nl
          , return_add_generic_AC_RND_CONV_false_11_and_9_nl , return_add_generic_AC_RND_CONV_false_11_and_10_nl
          , return_add_generic_AC_RND_CONV_false_11_and_11_nl , return_add_generic_AC_RND_CONV_false_11_and_12_nl
          , return_add_generic_AC_RND_CONV_false_11_and_13_cse , return_add_generic_AC_RND_CONV_false_11_and_14_cse
          , return_add_generic_AC_RND_CONV_false_11_and_15_cse , return_add_generic_AC_RND_CONV_false_11_and_16_cse
          , (fsm_output[37]) , return_add_generic_AC_RND_CONV_false_11_and_17_nl
          , return_add_generic_AC_RND_CONV_false_11_and_18_nl , return_add_generic_AC_RND_CONV_false_11_and_19_nl
          , return_add_generic_AC_RND_CONV_false_11_and_20_nl , return_add_generic_AC_RND_CONV_false_11_and_21_nl
          , return_add_generic_AC_RND_CONV_false_11_and_22_nl});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm
          <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm
          <= 1'b0;
    end
    else if ( run_wen & (~((fsm_output[40]) | (fsm_output[42]) | (fsm_output[41])
        | (fsm_output[39]) | (fsm_output[38]) | (fsm_output[33]) | or_dcpl_500 |
        (fsm_output[35]) | or_dcpl_597 | (fsm_output[11]))) ) begin
      return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm
          <= MUX1HOT_s_1_4_2((return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_and_5_cse[51]),
          return_extract_12_return_extract_12_or_1_cse_sva_1, return_extract_15_return_extract_15_nor_cse_sva_mx1,
          return_add_generic_AC_RND_CONV_false_13_op1_mu_52_lpi_3_dfm_1, {return_add_generic_AC_RND_CONV_false_13_or_nl
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_12_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_13_cse
          , (fsm_output[31])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_22_op1_mu_52_lpi_3_dfm <= 1'b0;
      stage_PE_1_x_re_d_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_22_op1_mu_52_lpi_3_dfm <= 1'b0;
      stage_PE_1_x_re_d_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_22_op1_mu_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_22_op1_mu_52_lpi_3_dfm <= MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_op2_mu_52_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_13_op1_mu_52_lpi_3_dfm_1, fsm_output[30]);
      stage_PE_1_x_re_d_sva <= MUX_v_64_2_2(out_f_d_rsci_q_d, in_f_d_rsci_q_d, fsm_output[30]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_mux_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_mux_itm <= 1'b0;
    end
    else if ( run_wen & ((~(inverse_lpi_1_dfm_1 | or_dcpl_769 | or_dcpl_531 | or_dcpl_870
        | (fsm_output[42]) | (fsm_output[20]) | (fsm_output[41]) | (fsm_output[39])
        | or_dcpl_705 | or_dcpl_518 | or_dcpl_597 | (fsm_output[19]) | or_dcpl_438))
        | (fsm_output[5]) | (fsm_output[16]) | (fsm_output[30]) | (fsm_output[43]))
        ) begin
      return_add_generic_AC_RND_CONV_false_11_mux_itm <= MUX1HOT_s_1_12_2(return_add_generic_AC_RND_CONV_false_2_if_2_return_add_generic_AC_RND_CONV_false_2_if_2_nor_1_nl,
          (out_f_d_rsci_q_d[63]), (~ (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[6])), return_add_generic_AC_RND_CONV_false_11_if_2_return_add_generic_AC_RND_CONV_false_11_if_2_nor_mx2w0,
          (stage_PE_1_x_re_d_sva[63]), (~ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1),
          return_add_generic_AC_RND_CONV_false_15_if_2_return_add_generic_AC_RND_CONV_false_15_if_2_nor_1_nl,
          (in_f_d_rsci_q_d[63]), operator_11_true_33_operator_11_true_33_and_tmp,
          return_add_generic_AC_RND_CONV_false_10_if_2_return_add_generic_AC_RND_CONV_false_10_if_2_and_1_mx5w0,
          (stage_PE_1_x_im_d_sva[63]), return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva,
          {return_add_generic_AC_RND_CONV_false_11_and_23_cse , return_add_generic_AC_RND_CONV_false_11_and_31_cse
          , return_add_generic_AC_RND_CONV_false_11_or_nl , return_add_generic_AC_RND_CONV_false_17_and_3_cse
          , return_add_generic_AC_RND_CONV_false_17_and_9_cse , return_add_generic_AC_RND_CONV_false_17_and_10_cse
          , return_add_generic_AC_RND_CONV_false_11_and_27_nl , return_add_generic_AC_RND_CONV_false_11_and_35_nl
          , (fsm_output[31]) , return_add_generic_AC_RND_CONV_false_17_and_5_cse
          , return_add_generic_AC_RND_CONV_false_17_and_11_cse , return_add_generic_AC_RND_CONV_false_17_and_12_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_do_sub_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_do_sub_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_882 | or_dcpl_576 | (fsm_output[38]) | or_dcpl_99
        | or_dcpl_556 | or_dcpl_135 | or_dcpl_133 | (fsm_output[16]) | or_dcpl_401))
        ) begin
      return_add_generic_AC_RND_CONV_false_11_do_sub_sva <= MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_2_do_sub_return_add_generic_AC_RND_CONV_false_2_do_sub_return_add_generic_AC_RND_CONV_false_2_do_sub_xnor_nl,
          return_add_generic_AC_RND_CONV_false_6_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_xnor_nl,
          return_add_generic_AC_RND_CONV_false_15_do_sub_return_add_generic_AC_RND_CONV_false_15_do_sub_return_add_generic_AC_RND_CONV_false_15_do_sub_xnor_nl,
          return_add_generic_AC_RND_CONV_false_22_do_sub_return_add_generic_AC_RND_CONV_false_22_do_sub_xor_nl,
          {(fsm_output[5]) , or_dcpl_404 , (fsm_output[14]) , (fsm_output[30]) ,
          (fsm_output[39])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_do_sub_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_do_sub_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_790 | or_dcpl_870 | or_dcpl_580 | or_dcpl_579
        | (fsm_output[41]) | (fsm_output[21]) | or_dcpl_574)) ) begin
      return_add_generic_AC_RND_CONV_false_12_do_sub_sva <= MUX1HOT_s_1_6_2(xor_cse,
          xor_2_cse, return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_xnor_nl,
          xor_3_cse, xor_4_cse, return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_xnor_nl,
          {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[14]) , (fsm_output[30])
          , (fsm_output[32]) , (fsm_output[39])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_ls_sva <= 6'b000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_ls_sva <= 6'b000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_10_r_zero_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva <= all_same_out;
      return_add_generic_AC_RND_CONV_false_10_ls_sva <= rtn_out;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva <= 1'b0;
    end
    else if ( run_wen & ((inverse_lpi_1_dfm_1 & (~(and_dcpl_233 & and_dcpl_286 &
        and_dcpl_284 & (~((fsm_output[25:24]!=2'b00))) & (~ (fsm_output[41])) & (~((fsm_output[18:17]!=2'b00)))
        & (~((fsm_output[16]) | (fsm_output[31]))) & (~ (fsm_output[6])) & (~((fsm_output[29])
        | (fsm_output[4])))))) | (fsm_output[5]) | (fsm_output[19]) | (fsm_output[30])
        | (fsm_output[42]) | (fsm_output[45])) ) begin
      return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva <= MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp,
          all_same_out, return_add_generic_AC_RND_CONV_false_13_return_add_generic_AC_RND_CONV_false_13_or_1_tmp,
          {(fsm_output[5]) , return_add_generic_AC_RND_CONV_false_10_or_3_nl , (fsm_output[30])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_11_true_return_26_sva <= 1'b0;
    end
    else if ( rst ) begin
      operator_11_true_return_26_sva <= 1'b0;
    end
    else if ( run_wen & ((inverse_lpi_1_dfm_1 & (~(or_dcpl_882 | or_dcpl_707 | (fsm_output[13])
        | or_dcpl_906 | or_dcpl_780 | (fsm_output[35]) | or_dcpl_514 | or_dcpl_440
        | (fsm_output[17]) | or_dcpl_666))) | (fsm_output[5]) | (fsm_output[6]) |
        (fsm_output[18]) | (fsm_output[30]) | (fsm_output[41])) ) begin
      operator_11_true_return_26_sva <= MUX1HOT_s_1_17_2(return_add_generic_AC_RND_CONV_false_if_2_return_add_generic_AC_RND_CONV_false_if_2_and_2_nl,
          (out_f_d_rsci_q_d[63]), (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[6]), operator_11_true_24_operator_11_true_24_and_tmp,
          return_add_generic_AC_RND_CONV_false_1_if_2_return_add_generic_AC_RND_CONV_false_1_if_2_and_2_nl,
          (stage_PE_1_x_im_d_sva[63]), return_add_generic_AC_RND_CONV_false_1_op1_nan_sva_mx3w0,
          return_add_generic_AC_RND_CONV_false_10_if_2_return_add_generic_AC_RND_CONV_false_10_if_2_and_1_mx5w0,
          return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva,
          operator_11_true_33_operator_11_true_33_and_tmp, return_add_generic_AC_RND_CONV_false_13_if_2_return_add_generic_AC_RND_CONV_false_13_if_2_and_2_nl,
          (in_f_d_rsci_q_d[63]), return_add_generic_AC_RND_CONV_false_14_if_2_return_add_generic_AC_RND_CONV_false_14_if_2_and_2_nl,
          return_add_generic_AC_RND_CONV_false_9_op2_nan_sva_mx7w0, return_add_generic_AC_RND_CONV_false_9_if_2_return_add_generic_AC_RND_CONV_false_9_if_2_and_1_mx2w0,
          (stage_PE_1_x_re_d_sva[63]), return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1,
          {return_add_generic_AC_RND_CONV_false_11_and_23_cse , return_extract_26_exception_or_nl
          , return_extract_26_exception_or_4_nl , (fsm_output[6]) , return_extract_26_exception_and_4_nl
          , return_extract_26_exception_or_5_nl , (fsm_output[8]) , return_extract_26_exception_and_6_cse
          , return_extract_26_exception_and_18_cse , return_extract_26_exception_and_8_nl
          , and_493_nl , return_extract_26_exception_or_6_nl , return_extract_26_exception_and_9_nl
          , (fsm_output[33]) , return_extract_26_exception_and_11_cse , return_extract_26_exception_and_21_cse
          , return_extract_26_exception_and_22_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_33_true_12_acc_psp_sva <= 13'b0000000000000;
    end
    else if ( rst ) begin
      operator_33_true_12_acc_psp_sva <= 13'b0000000000000;
    end
    else if ( run_wen & mode_lpi_1_dfm ) begin
      operator_33_true_12_acc_psp_sva <= z_out_8;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm
          <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm
          <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_919 | or_dcpl_631 | or_dcpl_514 | (fsm_output[11])
        | (fsm_output[6]))) ) begin
      return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm
          <= MUX1HOT_v_51_4_2((return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_and_5_cse[50:0]),
          (out_f_d_rsci_q_d[51:1]), (out_f_d_rsci_q_d[50:0]), return_extract_32_mux_4_cse,
          {return_add_generic_AC_RND_CONV_false_10_or_4_nl , and_498_nl , return_add_generic_AC_RND_CONV_false_10_and_4_nl
          , (fsm_output[31])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_unequal_tmp <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & ((inverse_lpi_1_dfm_1 & (~(or_dcpl_929 | or_dcpl_928 | or_dcpl_101
        | (fsm_output[39]) | or_dcpl_799 | or_dcpl_776 | (fsm_output[32]) | or_dcpl_136
        | (fsm_output[35]) | or_dcpl_514 | or_dcpl_713))) | (fsm_output[6]) | (fsm_output[21])
        | (fsm_output[31]) | (fsm_output[46])) ) begin
      return_add_generic_AC_RND_CONV_false_10_unequal_tmp <= MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp,
          return_add_generic_AC_RND_CONV_false_3_r_nan_and_nl, return_add_generic_AC_RND_CONV_false_2_r_nan_and_2,
          return_add_generic_AC_RND_CONV_false_13_return_add_generic_AC_RND_CONV_false_13_or_1_tmp,
          return_add_generic_AC_RND_CONV_false_16_r_nan_and_nl, return_add_generic_AC_RND_CONV_false_24_r_nan_and_nl,
          {(fsm_output[6]) , (fsm_output[9]) , (fsm_output[21]) , (fsm_output[31])
          , (fsm_output[34]) , (fsm_output[46])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_23_op1_nan_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_23_op1_inf_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_23_op1_nan_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_23_op1_inf_sva <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_23_op1_nan_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_23_op1_nan_sva <= MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_op1_nan_sva_1,
          return_extract_58_and_2_nl, fsm_output[43]);
      return_add_generic_AC_RND_CONV_false_23_op1_inf_sva <= MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_9_op1_inf_sva_1,
          return_extract_58_and_1_nl, fsm_output[43]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_14_op2_nan_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_14_op2_nan_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_949 | or_dcpl_561 | or_dcpl_928 | or_dcpl_788
        | (fsm_output[41]) | (fsm_output[21]) | (fsm_output[34]) | (fsm_output[8])
        | or_dcpl_517 | or_dcpl_940 | (fsm_output[18]) | or_dcpl_573)) ) begin
      return_add_generic_AC_RND_CONV_false_14_op2_nan_sva <= MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_1_op1_nan_sva_mx3w0,
          return_add_generic_AC_RND_CONV_false_9_do_sub_return_add_generic_AC_RND_CONV_false_9_do_sub_xor_nl,
          return_add_generic_AC_RND_CONV_false_9_op2_nan_sva_mx7w0, return_add_generic_AC_RND_CONV_false_10_op2_nan_sva_1,
          return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_xnor_nl,
          return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1, {(fsm_output[6])
          , (fsm_output[14]) , (fsm_output[20]) , (fsm_output[33]) , (fsm_output[39])
          , (fsm_output[47])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_14_op2_inf_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_14_op2_inf_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_949 | or_dcpl_961 | (fsm_output[40]) | (fsm_output[15])
        | (fsm_output[42]) | (fsm_output[41]) | or_dcpl_682 | or_dcpl_906 | or_dcpl_704
        | (fsm_output[7]) | or_dcpl_953 | or_dcpl_573)) ) begin
      return_add_generic_AC_RND_CONV_false_14_op2_inf_sva <= MUX1HOT_s_1_6_2(return_extract_2_and_1_tmp,
          return_add_generic_AC_RND_CONV_false_8_do_sub_return_add_generic_AC_RND_CONV_false_8_do_sub_xor_nl,
          return_add_generic_AC_RND_CONV_false_9_op2_inf_sva_1, return_add_generic_AC_RND_CONV_false_10_op2_inf_sva_1,
          return_add_generic_AC_RND_CONV_false_21_do_sub_return_add_generic_AC_RND_CONV_false_21_do_sub_xor_nl,
          return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1, {(fsm_output[6])
          , (fsm_output[12]) , (fsm_output[20]) , (fsm_output[33]) , (fsm_output[37])
          , (fsm_output[47])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_ls_sva <= 6'b000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_ls_sva <= 6'b000000;
    end
    else if ( run_wen & (~(or_dcpl_937 | or_dcpl_560 | (fsm_output[22]) | (fsm_output[43])
        | or_dcpl_125 | or_dcpl_99 | or_dcpl_422)) ) begin
      return_add_generic_AC_RND_CONV_false_11_ls_sva <= rtn_out;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_x_im_d_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      stage_PE_1_x_im_d_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_919 | or_dcpl_556 | or_dcpl_552 | (fsm_output[37])
        | or_dcpl_840 | or_dcpl_573)) ) begin
      stage_PE_1_x_im_d_sva <= MUX_v_64_2_2(out_f_d_rsci_q_d, in_f_d_rsci_q_d, fsm_output[31]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_tmp_re_d_1_sva_1_63_57 <= 7'b0000000;
    end
    else if ( rst ) begin
      stage_PE_1_tmp_re_d_1_sva_1_63_57 <= 7'b0000000;
    end
    else if ( stage_PE_1_tmp_re_d_and_ssc ) begin
      stage_PE_1_tmp_re_d_1_sva_1_63_57 <= MUX_v_7_2_2((out_f_d_rsci_q_d[63:57]),
          (in_f_d_rsci_q_d[63:57]), fsm_output[32]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      drf_qr_lval_11_smx_lpi_3_dfm_10 <= 1'b0;
      drf_qr_lval_11_smx_lpi_3_dfm_9 <= 1'b0;
      drf_qr_lval_11_smx_lpi_3_dfm_8_5 <= 4'b0000;
      drf_qr_lval_11_smx_lpi_3_dfm_4_0 <= 5'b00000;
    end
    else if ( rst ) begin
      drf_qr_lval_11_smx_lpi_3_dfm_10 <= 1'b0;
      drf_qr_lval_11_smx_lpi_3_dfm_9 <= 1'b0;
      drf_qr_lval_11_smx_lpi_3_dfm_8_5 <= 4'b0000;
      drf_qr_lval_11_smx_lpi_3_dfm_4_0 <= 5'b00000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_8_exp_and_ssc ) begin
      drf_qr_lval_11_smx_lpi_3_dfm_10 <= MUX1HOT_s_1_6_2((drf_qr_lval_1_smx_lpi_3_dfm_mx1[10]),
          (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
          BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1, (drf_qr_lval_11_smx_lpi_3_dfm_mx2[10]),
          (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
          (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1[1]), {(fsm_output[7])
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_4_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse
          , (fsm_output[32]) , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_cse});
      drf_qr_lval_11_smx_lpi_3_dfm_9 <= MUX1HOT_s_1_6_2((drf_qr_lval_1_smx_lpi_3_dfm_mx1[9]),
          (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[9]),
          (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[4]), (drf_qr_lval_11_smx_lpi_3_dfm_mx2[9]),
          (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[9]),
          (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1[0]), {(fsm_output[7])
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_4_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse
          , (fsm_output[32]) , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_cse});
      drf_qr_lval_11_smx_lpi_3_dfm_8_5 <= MUX1HOT_v_4_6_2((drf_qr_lval_1_smx_lpi_3_dfm_mx1[8:5]),
          (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[8:5]),
          (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[3:0]), (drf_qr_lval_11_smx_lpi_3_dfm_mx2[8:5]),
          (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[8:5]),
          (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[8:5]), {(fsm_output[7])
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_4_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse
          , (fsm_output[32]) , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_cse});
      drf_qr_lval_11_smx_lpi_3_dfm_4_0 <= MUX1HOT_v_5_6_2((drf_qr_lval_1_smx_lpi_3_dfm_mx1[4:0]),
          (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[4:0]),
          reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1, (drf_qr_lval_11_smx_lpi_3_dfm_mx2[4:0]),
          (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[4:0]),
          (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[4:0]), {(fsm_output[7])
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_4_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse
          , (fsm_output[32]) , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_mux_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_mux_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_1001 | or_dcpl_999 | or_dcpl_788 | or_dcpl_750
        | or_dcpl_99 | (fsm_output[8]) | or_dcpl_953 | or_dcpl_440)) ) begin
      return_add_generic_AC_RND_CONV_false_12_mux_itm <= MUX1HOT_s_1_10_2(return_add_generic_AC_RND_CONV_false_3_if_2_return_add_generic_AC_RND_CONV_false_3_if_2_nor_1_nl,
          (stage_PE_1_x_im_d_sva[63]), (~ (out_f_d_rsci_q_d[63])), return_add_generic_AC_RND_CONV_false_12_if_2_return_add_generic_AC_RND_CONV_false_12_if_2_nor_mx4w0,
          (~ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva),
          return_add_generic_AC_RND_CONV_false_16_if_2_return_add_generic_AC_RND_CONV_false_16_if_2_nor_1_nl,
          (~ (in_f_d_rsci_q_d[63])), return_add_generic_AC_RND_CONV_false_11_if_2_return_add_generic_AC_RND_CONV_false_11_if_2_nor_mx2w0,
          (stage_PE_1_x_re_d_sva[63]), (~ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1),
          {return_add_generic_AC_RND_CONV_false_12_and_1_nl , return_add_generic_AC_RND_CONV_false_12_or_nl
          , return_add_generic_AC_RND_CONV_false_12_and_10_nl , return_extract_26_exception_and_6_cse
          , return_extract_26_exception_and_18_cse , return_add_generic_AC_RND_CONV_false_12_and_5_nl
          , return_add_generic_AC_RND_CONV_false_12_and_14_nl , return_extract_26_exception_and_11_cse
          , return_extract_26_exception_and_21_cse , return_extract_26_exception_and_22_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_16_do_sub_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_16_do_sub_sva <= 1'b0;
    end
    else if ( run_wen & (~(return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
        | or_dcpl_682 | or_dcpl_607 | return_extract_26_exception_or_3_cse)) ) begin
      return_add_generic_AC_RND_CONV_false_16_do_sub_sva <= MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_3_do_sub_return_add_generic_AC_RND_CONV_false_3_do_sub_return_add_generic_AC_RND_CONV_false_3_do_sub_xnor_nl,
          return_add_generic_AC_RND_CONV_false_7_do_sub_return_add_generic_AC_RND_CONV_false_7_do_sub_xor_nl,
          return_add_generic_AC_RND_CONV_false_16_do_sub_return_add_generic_AC_RND_CONV_false_16_do_sub_return_add_generic_AC_RND_CONV_false_16_do_sub_xnor_nl,
          return_add_generic_AC_RND_CONV_false_20_do_sub_return_add_generic_AC_RND_CONV_false_20_do_sub_xor_nl,
          {(fsm_output[7]) , (fsm_output[12]) , (fsm_output[32]) , (fsm_output[37])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_op1_inf_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_op1_inf_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_128 | or_dcpl_126 | or_dcpl_749 | or_dcpl_575
        | or_dcpl_99 | or_dcpl_1015 | or_dcpl_597 | or_dcpl_440)) ) begin
      return_add_generic_AC_RND_CONV_false_10_op1_inf_sva <= MUX1HOT_s_1_4_2(return_extract_2_and_1_tmp,
          return_extract_26_and_1_nl, return_add_generic_AC_RND_CONV_false_9_op2_inf_sva_1,
          return_add_generic_AC_RND_CONV_false_19_op1_inf_sva_1, {(fsm_output[8])
          , (fsm_output[18]) , (fsm_output[31]) , (fsm_output[35])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_op2_nan_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_op2_inf_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_op2_nan_sva <= 1'b0;
      return_add_generic_AC_RND_CONV_false_10_op2_inf_sva <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_10_op2_nan_and_cse ) begin
      return_add_generic_AC_RND_CONV_false_10_op2_nan_sva <= MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_9_op1_nan_sva_1,
          return_add_generic_AC_RND_CONV_false_6_op2_nan_sva_1, return_add_generic_AC_RND_CONV_false_10_op2_nan_sva_1,
          return_add_generic_AC_RND_CONV_false_19_op2_nan_sva_1, return_add_generic_AC_RND_CONV_false_23_op2_nan_sva_1,
          return_add_generic_AC_RND_CONV_false_22_op2_nan_sva_1, {(fsm_output[8])
          , (fsm_output[12]) , or_tmp_771 , (fsm_output[37]) , (fsm_output[41]) ,
          (fsm_output[45])});
      return_add_generic_AC_RND_CONV_false_10_op2_inf_sva <= MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_9_op1_inf_sva_1,
          return_add_generic_AC_RND_CONV_false_6_op2_inf_sva_1, return_add_generic_AC_RND_CONV_false_10_op2_inf_sva_1,
          return_add_generic_AC_RND_CONV_false_19_op2_inf_sva_1, return_add_generic_AC_RND_CONV_false_23_op2_inf_sva_1,
          return_add_generic_AC_RND_CONV_false_22_op2_inf_sva_1, {(fsm_output[8])
          , (fsm_output[12]) , or_tmp_771 , (fsm_output[37]) , (fsm_output[41]) ,
          (fsm_output[45])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0 <= 52'b0000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0 <= 52'b0000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & ((or_dcpl_48 & (~(return_add_generic_AC_RND_CONV_false_23_op1_inf_sva
        | return_add_generic_AC_RND_CONV_false_23_op1_nan_sva)) & (~(return_add_generic_AC_RND_CONV_false_14_op2_inf_sva
        | return_add_generic_AC_RND_CONV_false_14_op2_nan_sva | return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva))
        & stage_PE_1_and_1_tmp) | (or_dcpl_49 & and_dcpl_28 & (~(return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
        | operator_11_true_return_26_sva | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva))
        & stage_PE_1_and_1_tmp) | (and_dcpl_36 & (~(return_add_generic_AC_RND_CONV_false_10_op1_nan_sva
        | return_add_generic_AC_RND_CONV_false_22_op1_inf_sva)) & and_dcpl_32) |
        ((~((nand_12_cse & return_add_generic_AC_RND_CONV_false_20_acc_3_itm_11_1)
        | operator_11_true_return_15_sva)) & (~(operator_11_true_return_1_sva | all_same_out))
        & mode_lpi_1_dfm) | (or_dcpl_49 & (~ return_add_generic_AC_RND_CONV_false_10_op2_inf_sva)
        & (~(return_add_generic_AC_RND_CONV_false_10_op2_nan_sva | operator_11_true_return_17_sva))
        & and_dcpl_32) | (or_dcpl_48 & and_dcpl_28 & and_dcpl_63 & (~ return_add_generic_AC_RND_CONV_false_11_r_zero_1_sva)
        & stage_PE_1_and_1_tmp) | (or_dcpl_49 & (~(return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
        | return_add_generic_AC_RND_CONV_false_14_op2_inf_sva)) & (~(return_add_generic_AC_RND_CONV_false_14_op2_nan_sva
        | operator_11_true_return_26_sva | return_add_generic_AC_RND_CONV_false_10_r_zero_1_sva))
        & stage_PE_1_and_1_tmp) | (and_dcpl_36 & and_dcpl_63 & and_dcpl_32)) ) begin
      return_add_generic_AC_RND_CONV_false_15_res_rounded_lpi_3_dfm_51_0 <= return_add_generic_AC_RND_CONV_false_2_return_add_generic_AC_RND_CONV_false_2_and_5_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva
          <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva
          <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_449 | (fsm_output[41]) | (fsm_output[17]) | (fsm_output[16])))
        ) begin
      return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva
          <= MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_6_return_add_generic_AC_RND_CONV_false_6_if_return_add_generic_AC_RND_CONV_false_6_op1_normal_return_extract_12_nor_tmp,
          return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva_mx1,
          return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_tmp,
          return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva_mx2,
          {(fsm_output[10]) , (fsm_output[14]) , (fsm_output[35]) , (fsm_output[39])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_10_op1_nan_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_10_op1_nan_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_1001 | or_dcpl_999 | or_dcpl_789 | or_dcpl_462
        | or_dcpl_716 | or_dcpl_514 | or_dcpl_440)) ) begin
      return_add_generic_AC_RND_CONV_false_10_op1_nan_sva <= MUX1HOT_s_1_5_2(return_add_generic_AC_RND_CONV_false_6_op1_nan_sva_1,
          return_extract_26_and_2_nl, return_add_generic_AC_RND_CONV_false_9_op2_nan_sva_mx7w0,
          return_add_generic_AC_RND_CONV_false_19_op1_nan_sva_1, return_extract_56_and_2_nl,
          {(fsm_output[10]) , (fsm_output[18]) , (fsm_output[31]) , (fsm_output[35])
          , (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_22_op1_inf_sva <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_22_op1_inf_sva <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_108 | or_dcpl_465 | (fsm_output[45]) | (fsm_output[43])
        | (fsm_output[42]) | (fsm_output[13]) | (fsm_output[34]) | (fsm_output[35])
        | or_dcpl_840)) ) begin
      return_add_generic_AC_RND_CONV_false_22_op1_inf_sva <= MUX1HOT_s_1_3_2(return_add_generic_AC_RND_CONV_false_6_op1_inf_sva_1,
          return_add_generic_AC_RND_CONV_false_9_op2_inf_sva_1, return_extract_56_and_1_nl,
          {(fsm_output[10]) , (fsm_output[33]) , (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & ((~(return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_6_nl
        | or_dcpl_488 | or_dcpl_503 | (fsm_output[38]) | (fsm_output[36]) | or_dcpl_440))
        | (fsm_output[10]) | (fsm_output[12]) | (fsm_output[16]) | (fsm_output[18])
        | (fsm_output[35]) | (fsm_output[37]) | (fsm_output[41])) ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm <= MUX1HOT_v_50_15_2((stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0[50:1]),
          (stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0[49:0]), (return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1[49:0]),
          (return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1[50:1]), return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[49:0]),
          return_add_generic_AC_RND_CONV_false_10_op2_mu_1_50_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49:0]),
          (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1[50:1]), (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1[49:0]),
          (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[49:0]), (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[50:1]),
          return_add_generic_AC_RND_CONV_false_20_op2_mu_1_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0,
          {return_add_generic_AC_RND_CONV_false_11_op_smaller_and_12_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_13_cse
          , return_add_generic_AC_RND_CONV_false_12_op_bigger_and_8_cse , return_add_generic_AC_RND_CONV_false_12_op_bigger_and_9_cse
          , (fsm_output[14]) , return_add_generic_AC_RND_CONV_false_11_exp_and_2_cse
          , return_add_generic_AC_RND_CONV_false_11_exp_and_3_cse , return_add_generic_AC_RND_CONV_false_10_exp_and_2_cse
          , return_add_generic_AC_RND_CONV_false_12_op_bigger_or_4_nl , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_14_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_15_cse , return_add_generic_AC_RND_CONV_false_10_exp_and_6_cse
          , return_add_generic_AC_RND_CONV_false_10_exp_and_7_cse , (fsm_output[39])
          , return_add_generic_AC_RND_CONV_false_10_exp_and_4_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_56_50 <= 7'b0000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_56_50 <= 7'b0000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_12_res_mant_and_ssc & and_dcpl_1
        ) begin
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_56_50 <= z_out_30[56:50];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_49_0 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_49_0 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_12_res_mant_and_ssc & (~(return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse
        | and_1013_cse | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_34_cse))
        ) begin
      return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_49_0 <= MUX1HOT_v_50_12_2((return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1[50:1]),
          (return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1[49:0]), return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[49:0]),
          (return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1[50:1]), (return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1[49:0]),
          return_add_generic_AC_RND_CONV_false_20_op2_mu_1_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0,
          (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49:0]),
          return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0, (z_out_30[49:0]),
          {return_add_generic_AC_RND_CONV_false_11_op_bigger_and_24_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_23_cse
          , and_1598_cse , or_tmp_348 , return_add_generic_AC_RND_CONV_false_12_res_mant_return_add_generic_AC_RND_CONV_false_12_res_mant_return_add_generic_AC_RND_CONV_false_12_res_mant_or_nl
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_30_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_29_cse
          , and_1608_cse , or_tmp_823 , return_add_generic_AC_RND_CONV_false_10_exp_and_5_cse
          , and_1163_cse , return_add_generic_AC_RND_CONV_false_12_res_mant_or_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm <= 1'b0;
    end
    else if ( run_wen & ((~(and_dcpl_267 | return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
        | or_dcpl_788 | or_dcpl_423 | or_dcpl_940)) | (fsm_output[11]) | (fsm_output[12])
        | (fsm_output[16]) | (fsm_output[18]) | (fsm_output[35]) | (fsm_output[37])
        | (fsm_output[39]) | (fsm_output[41])) ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm <= MUX1HOT_s_1_13_2(return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm_mx0w4,
          (return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1[50]), drf_qr_lval_14_smx_0_lpi_3_dfm_mx1,
          return_add_generic_AC_RND_CONV_false_7_op2_mu_1_51_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_21_cse,
          return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1,
          return_extract_15_return_extract_15_nor_cse_sva_mx2, stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx2_50,
          return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_2_nl,
          return_add_generic_AC_RND_CONV_false_20_op2_mu_1_51_lpi_3_dfm_mx0, drf_qr_lval_13_smx_0_lpi_3_dfm,
          return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_27_cse, {(fsm_output[11])
          , return_add_generic_AC_RND_CONV_false_12_op_bigger_and_8_cse , return_add_generic_AC_RND_CONV_false_12_op_bigger_and_9_cse
          , (fsm_output[14]) , (fsm_output[16]) , return_add_generic_AC_RND_CONV_false_10_exp_and_2_cse
          , return_add_generic_AC_RND_CONV_false_10_exp_and_3_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_14_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_15_cse , (fsm_output[37])
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_cse
          , (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm <= 1'b0;
    end
    else if ( run_wen & (~ or_tmp_852) ) begin
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm <= MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_7_op1_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_31_cse,
          return_add_generic_AC_RND_CONV_false_20_op2_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_20_op1_mu_1_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_34_cse, return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
          {return_add_generic_AC_RND_CONV_false_11_op_bigger_and_33_nl , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_34_cse
          , (fsm_output[16]) , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_35_nl
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse , (fsm_output[41])
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_15_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_16_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_itm <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_itm <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_12_op_bigger_and_2_cse ) begin
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm <= MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_7_op2_mu_1_52_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_6_cse,
          return_add_generic_AC_RND_CONV_false_10_op2_mu_1_51_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[50]),
          return_add_generic_AC_RND_CONV_false_20_op2_mu_1_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm,
          return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_12_cse, {return_add_generic_AC_RND_CONV_false_11_op_smaller_and_4_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse , (fsm_output[16])
          , return_add_generic_AC_RND_CONV_false_10_exp_and_2_cse , return_add_generic_AC_RND_CONV_false_10_exp_and_3_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_cse
          , (fsm_output[41])});
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_itm <= MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_7_op2_mu_1_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_8_op1_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_31_cse,
          return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx0, drf_qr_lval_13_smx_0_lpi_3_dfm,
          return_add_generic_AC_RND_CONV_false_20_op2_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_21_op1_mu_1_0_lpi_3_dfm_1,
          return_add_generic_AC_RND_CONV_false_11_op_bigger_mux1h_34_cse, {return_add_generic_AC_RND_CONV_false_11_op_smaller_and_4_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse , (fsm_output[16])
          , return_add_generic_AC_RND_CONV_false_10_exp_and_2_cse , return_add_generic_AC_RND_CONV_false_10_exp_and_3_cse
          , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_cse
          , (fsm_output[41])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_51_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_52_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva <= 6'b000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_51_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_52_lpi_3_dfm <= 1'b0;
      return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva <= 6'b000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_12_op_smaller_and_1_cse ) begin
      return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_51_lpi_3_dfm <= MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_51_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_cse, return_add_generic_AC_RND_CONV_false_5_op_smaller_mux_1_cse,
          return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_51_lpi_3_dfm_mx3,
          return_add_generic_AC_RND_CONV_false_5_op_smaller_mux_cse, return_add_generic_AC_RND_CONV_false_9_op1_mu_mux_2_cse,
          {(fsm_output[14]) , (fsm_output[16]) , (fsm_output[18]) , (fsm_output[39])
          , (fsm_output[41]) , (fsm_output[43])});
      return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_52_lpi_3_dfm <= MUX1HOT_s_1_6_2(return_add_generic_AC_RND_CONV_false_7_op_smaller_qr_52_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_22_op1_mu_mux_cse, return_add_generic_AC_RND_CONV_false_10_exp_mux_5_cse,
          return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_52_lpi_3_dfm_mx3,
          return_add_generic_AC_RND_CONV_false_22_op1_mu_mux_1_cse, return_add_generic_AC_RND_CONV_false_13_mux_25_cse,
          {(fsm_output[14]) , (fsm_output[16]) , (fsm_output[18]) , (fsm_output[39])
          , (fsm_output[41]) , (fsm_output[43])});
      return_add_generic_AC_RND_CONV_false_12_e_dif_sat_sva <= MUX1HOT_v_6_5_2(return_add_generic_AC_RND_CONV_false_21_e_dif_sat_or_cse,
          return_add_generic_AC_RND_CONV_false_9_e_dif_sat_sva_1, return_add_generic_AC_RND_CONV_false_12_e_dif_sat_or_cse,
          return_add_generic_AC_RND_CONV_false_8_e_dif_sat_or_cse, return_add_generic_AC_RND_CONV_false_25_e_dif_sat_or_nl,
          {(fsm_output[14]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse
          , (fsm_output[18]) , (fsm_output[39]) , (fsm_output[43])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_12_ls_sva <= 6'b000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_12_ls_sva <= 6'b000000;
    end
    else if ( run_wen & (~(or_dcpl_929 | (fsm_output[46]) | (fsm_output[45]) | (fsm_output[22])
        | or_dcpl_126 | (fsm_output[21]) | or_dcpl_550)) ) begin
      return_add_generic_AC_RND_CONV_false_12_ls_sva <= rtn_out;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0 <= 5'b00000;
    end
    else if ( rst ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0 <= 5'b00000;
    end
    else if ( BUTTERFLY_1_else_1_if_and_ssc ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0 <= MUX_v_5_2_2((out_u_rsci_q_d[15:11]),
          (in_u_rsci_q_d[15:11]), or_dcpl_118);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1 <= 2'b00;
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2 <= 9'b000000000;
    end
    else if ( rst ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1 <= 2'b00;
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2 <= 9'b000000000;
    end
    else if ( BUTTERFLY_1_else_1_if_and_1_cse ) begin
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1 <= MUX1HOT_v_2_4_2((out_u_rsci_q_d[10:9]),
          (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1[10:9]),
          (return_mult_generic_AC_RND_CONV_false_4_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w2[10:9]),
          (in_u_rsci_q_d[10:9]), {or_dcpl_95 , BUTTERFLY_1_else_1_if_and_3_cse ,
          (fsm_output[37]) , or_dcpl_118});
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2 <= MUX1HOT_v_9_5_2((out_u_rsci_q_d[8:0]),
          (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1[8:0]),
          (return_mult_generic_AC_RND_CONV_false_4_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w2[8:0]),
          BUTTERFLY_n_and_nl, (in_u_rsci_q_d[8:0]), {or_dcpl_95 , BUTTERFLY_1_else_1_if_and_3_cse
          , (fsm_output[37]) , or_1355_nl , or_dcpl_118});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_0 <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_0 <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_15_op_bigger_and_ssc ) begin
      return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_0 <= MUX1HOT_s_1_7_2((return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_itm[50]),
          (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_1_itm[50]), (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_2_itm[50]),
          (return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1[50]), (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_7_itm[50]),
          (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_8_itm[50]), (return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1[50]),
          {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , (fsm_output[5])
          , (fsm_output[7]) , (fsm_output[12]) , (fsm_output[30]) , (fsm_output[32])
          , (fsm_output[35])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_15_op_bigger_and_ssc & (~ or_tmp_852)
        ) begin
      return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1 <= MUX1HOT_v_50_15_2((return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_itm[49:0]),
          (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_1_itm[49:0]),
          (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_2_itm[49:0]),
          (return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1[49:0]), return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_49_0,
          return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[49:0]),
          return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_20_op2_mu_1_50_1_lpi_3_dfm_mx0,
          (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49:0]),
          return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_23_op2_mu_1_50_1_lpi_3_dfm_mx0,
          (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_7_itm[49:0]),
          (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux1h_8_itm[49:0]),
          (return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1[49:0]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
          , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[12]) , or_1996_nl , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_34_cse
          , or_1998_nl , return_add_generic_AC_RND_CONV_false_11_exp_and_3_cse ,
          return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse , or_tmp_823
          , return_add_generic_AC_RND_CONV_false_10_exp_and_5_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_16_cse
          , (fsm_output[30]) , (fsm_output[32]) , (fsm_output[35])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_0 <= 1'b0;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_0 <= 1'b0;
    end
    else if ( return_add_generic_AC_RND_CONV_false_17_m_r_and_ssc ) begin
      return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_0 <= MUX1HOT_s_1_3_2((return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[50]),
          (return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1[50]), (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[50]),
          {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , (fsm_output[10])
          , (fsm_output[37])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1 <= 50'b00000000000000000000000000000000000000000000000000;
    end
    else if ( return_add_generic_AC_RND_CONV_false_17_m_r_and_ssc & (~ or_tmp_857)
        ) begin
      return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1 <= MUX1HOT_v_50_11_2((return_add_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[49:0]),
          (return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1[49:0]), return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm,
          return_add_generic_AC_RND_CONV_false_7_op2_mu_1_50_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[49:0]),
          return_add_generic_AC_RND_CONV_false_9_op2_mu_1_50_1_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[49:0]),
          return_add_generic_AC_RND_CONV_false_10_op2_mu_1_50_1_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_20_op2_mu_1_50_1_lpi_3_dfm_mx0,
          return_add_generic_AC_RND_CONV_false_22_op2_mu_1_50_1_lpi_3_dfm_mx0, (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1[49:0]),
          {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , (fsm_output[10])
          , or_2005_nl , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_5_cse
          , or_tmp_348 , return_add_generic_AC_RND_CONV_false_11_exp_and_3_cse ,
          or_2010_nl , return_add_generic_AC_RND_CONV_false_10_exp_and_3_cse , return_add_generic_AC_RND_CONV_false_11_op_smaller_and_7_cse
          , return_add_generic_AC_RND_CONV_false_10_exp_and_5_cse , (fsm_output[37])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_1 <= 1'b0;
    end
    else if ( rst ) begin
      BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_1 <= 1'b0;
    end
    else if ( run_wen & ((~ or_1670_ssc) | BUTTERFLY_1_else_2_or_cse | BUTTERFLY_1_else_2_and_27_cse)
        ) begin
      BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_1 <= MUX1HOT_s_1_14_2((z_out_40[10]),
          (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[5]), (out_f_d_rsci_q_d[62]), (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w3_10_1[9]),
          (stage_PE_1_tmp_re_d_1_sva_1_63_57[5]), (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5[5]),
          (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
          (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1[1]), (in_f_d_rsci_q_d[62]),
          (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w9_10_1[9]), (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5[5]),
          (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
          BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1, (z_out_45[10]), {BUTTERFLY_1_else_2_or_cse
          , or_tmp_561 , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
          , or_tmp_564 , return_add_generic_AC_RND_CONV_false_17_e_r_and_cse , or_1673_ssc
          , and_1598_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_34_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse , or_tmp_570
          , or_1678_ssc , and_1608_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse
          , BUTTERFLY_1_else_2_and_27_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd <= 1'b0;
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1 <= 4'b0000;
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2 <= 4'b0000;
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3 <= 1'b0;
    end
    else if ( rst ) begin
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd <= 1'b0;
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1 <= 4'b0000;
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2 <= 4'b0000;
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3 <= 1'b0;
    end
    else if ( BUTTERFLY_1_else_2_and_46_cse ) begin
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd <= MUX1HOT_s_1_20_2((O_1_out_1[61]),
          (O_1_out[61]), (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1[9]),
          (stage_PE_1_x_re_d_sva[62]), (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[9]),
          (stage_PE_1_x_im_d_sva[62]), (z_out_40[9]), (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[4]),
          (out_f_d_rsci_q_d[61]), (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w3_10_1[8]),
          (stage_PE_1_tmp_re_d_1_sva_1_63_57[4]), (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5[4]),
          (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[9]),
          (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1[0]), (in_f_d_rsci_q_d[61]),
          (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w9_10_1[8]), (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5[4]),
          (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[9]),
          (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[4]), (z_out_45[9]), {and_1153_rgt
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_6_cse , or_tmp_348
          , return_add_generic_AC_RND_CONV_false_11_exp_and_3_cse , and_1163_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_16_cse , BUTTERFLY_1_else_2_or_cse
          , or_tmp_561 , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
          , or_tmp_564 , return_add_generic_AC_RND_CONV_false_17_e_r_and_cse , or_1673_ssc
          , and_1598_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_34_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse , or_tmp_570
          , or_1678_ssc , and_1608_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse
          , BUTTERFLY_1_else_2_and_27_cse});
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1 <= MUX1HOT_v_4_20_2((O_1_out_1[60:57]),
          (O_1_out[60:57]), (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1[8:5]),
          (stage_PE_1_x_re_d_sva[61:58]), (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[8:5]),
          (stage_PE_1_x_im_d_sva[61:58]), (z_out_40[8:5]), (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[3:0]),
          (out_f_d_rsci_q_d[60:57]), (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w3_10_1[7:4]),
          (stage_PE_1_tmp_re_d_1_sva_1_63_57[3:0]), (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5[3:0]),
          (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[8:5]),
          (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[8:5]), (in_f_d_rsci_q_d[60:57]),
          (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w9_10_1[7:4]), (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5[3:0]),
          (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[8:5]),
          (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[3:0]), (z_out_45[8:5]), {and_1153_rgt
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_6_cse , or_tmp_348
          , return_add_generic_AC_RND_CONV_false_11_exp_and_3_cse , and_1163_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_16_cse , BUTTERFLY_1_else_2_or_cse
          , or_tmp_561 , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
          , or_tmp_564 , return_add_generic_AC_RND_CONV_false_17_e_r_and_cse , or_1673_ssc
          , and_1598_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_34_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse , or_tmp_570
          , or_1678_ssc , and_1608_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse
          , BUTTERFLY_1_else_2_and_27_cse});
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2 <= MUX1HOT_v_4_20_2((O_1_out_1[56:53]),
          (O_1_out[56:53]), (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1[4:1]),
          (stage_PE_1_x_re_d_sva[57:54]), (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[4:1]),
          (stage_PE_1_x_im_d_sva[57:54]), (z_out_40[4:1]), (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[56:53]),
          (out_f_d_rsci_q_d[56:53]), (stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w3_10_1[3:0]),
          (stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_0[5:2]), stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1,
          (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[4:1]),
          (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[4:1]), (in_f_d_rsci_q_d[56:53]),
          (stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w9_10_1[3:0]), stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1,
          (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[4:1]),
          (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[4:1]), (z_out_45[4:1]), {and_1153_rgt
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_6_cse , or_tmp_348
          , return_add_generic_AC_RND_CONV_false_11_exp_and_3_cse , and_1163_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_16_cse , BUTTERFLY_1_else_2_or_cse
          , or_tmp_561 , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
          , or_tmp_564 , return_add_generic_AC_RND_CONV_false_17_e_r_and_cse , or_1673_ssc
          , and_1598_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_34_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse , or_tmp_570
          , or_1678_ssc , and_1608_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse
          , BUTTERFLY_1_else_2_and_27_cse});
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3 <= MUX1HOT_s_1_20_2((O_1_out_1[52]),
          (O_1_out[52]), (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1[0]),
          (stage_PE_1_x_re_d_sva[53]), (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[0]),
          (stage_PE_1_x_im_d_sva[53]), (z_out_40[0]), (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[52]),
          (out_f_d_rsci_q_d[52]), stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0w3_0, (stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_0[1]),
          stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0, (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[0]),
          (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[0]), (in_f_d_rsci_q_d[52]),
          stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0w9_0, stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0,
          (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[0]),
          (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[0]), (z_out_45[0]), {and_1153_rgt
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_6_cse , or_tmp_348
          , return_add_generic_AC_RND_CONV_false_11_exp_and_3_cse , and_1163_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_16_cse , BUTTERFLY_1_else_2_or_cse
          , or_tmp_561 , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
          , or_tmp_564 , return_add_generic_AC_RND_CONV_false_17_e_r_and_cse , or_1673_ssc
          , and_1598_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_34_cse
          , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse , or_tmp_570
          , or_1678_ssc , and_1608_cse , return_add_generic_AC_RND_CONV_false_11_op_bigger_and_36_cse
          , BUTTERFLY_1_else_2_and_27_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_0 <= 3'b000;
    end
    else if ( rst ) begin
      BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_0 <= 3'b000;
    end
    else if ( BUTTERFLY_1_else_3_else_and_1_ssc ) begin
      BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_0 <= MUX1HOT_v_3_3_2((BUTTERFLY_1_else_3_else_mux1h_itm[13:11]),
          (z_out_4_31_16[13:11]), (z_out_38[13:11]), {or_1540_itm , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
          , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1 <= 1'b0;
    end
    else if ( rst ) begin
      BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1 <= 1'b0;
    end
    else if ( BUTTERFLY_1_else_3_else_and_1_ssc & (~ or_tmp_403) ) begin
      BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1 <= MUX1HOT_s_1_9_2((BUTTERFLY_1_else_3_else_mux1h_itm[10]),
          (z_out_4_31_16[10]), (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[5]), (out_f_d_rsci_q_d[62]),
          (stage_PE_1_x_im_d_sva[62]), (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w3[10]),
          (in_f_d_rsci_q_d[62]), (return_mult_generic_AC_RND_CONV_false_3_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w6[10]),
          (z_out_38[10]), {or_1540_itm , BUTTERFLY_1_else_3_else_and_11_cse , BUTTERFLY_1_else_3_else_and_26_cse
          , BUTTERFLY_1_else_3_else_and_27_cse , BUTTERFLY_1_else_3_else_and_28_cse
          , (fsm_output[12]) , BUTTERFLY_1_else_3_else_and_30_cse , (fsm_output[35])
          , BUTTERFLY_1_else_2_and_27_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd <= 5'b00000;
      reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1 <= 5'b00000;
    end
    else if ( rst ) begin
      reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd <= 5'b00000;
      reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1 <= 5'b00000;
    end
    else if ( BUTTERFLY_1_else_3_else_and_24_cse ) begin
      reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd <= MUX1HOT_v_5_13_2((BUTTERFLY_1_else_3_else_mux1h_itm[9:5]),
          (z_out_4_31_16[9:5]), (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[4:0]), (out_f_d_rsci_q_d[61:57]),
          (stage_PE_1_x_im_d_sva[61:57]), (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w3[9:5]),
          (in_f_d_rsci_q_d[61:57]), (return_mult_generic_AC_RND_CONV_false_3_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w6[9:5]),
          (z_out_38[9:5]), (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1[9:5]),
          (stage_PE_1_x_im_d_sva[62:58]), (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1[9:5]),
          (stage_PE_1_x_re_d_sva[62:58]), {or_1540_itm , BUTTERFLY_1_else_3_else_and_11_cse
          , BUTTERFLY_1_else_3_else_and_26_cse , BUTTERFLY_1_else_3_else_and_27_cse
          , BUTTERFLY_1_else_3_else_and_28_cse , (fsm_output[12]) , BUTTERFLY_1_else_3_else_and_30_cse
          , (fsm_output[35]) , BUTTERFLY_1_else_2_and_27_cse , and_2281_cse , return_add_generic_AC_RND_CONV_false_10_exp_and_3_cse
          , or_tmp_823 , return_add_generic_AC_RND_CONV_false_10_exp_and_5_cse});
      reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1 <= MUX1HOT_v_5_13_2((BUTTERFLY_1_else_3_else_mux1h_itm[4:0]),
          (z_out_4_31_16[4:0]), (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[56:52]), (out_f_d_rsci_q_d[56:52]),
          (stage_PE_1_x_im_d_sva[56:52]), (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w3[4:0]),
          (in_f_d_rsci_q_d[56:52]), (return_mult_generic_AC_RND_CONV_false_3_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w6[4:0]),
          (z_out_38[4:0]), (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1[4:0]),
          (stage_PE_1_x_im_d_sva[57:53]), (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1[4:0]),
          (stage_PE_1_x_re_d_sva[57:53]), {or_1540_itm , BUTTERFLY_1_else_3_else_and_11_cse
          , BUTTERFLY_1_else_3_else_and_26_cse , BUTTERFLY_1_else_3_else_and_27_cse
          , BUTTERFLY_1_else_3_else_and_28_cse , (fsm_output[12]) , BUTTERFLY_1_else_3_else_and_30_cse
          , (fsm_output[35]) , BUTTERFLY_1_else_2_and_27_cse , and_2281_cse , return_add_generic_AC_RND_CONV_false_10_exp_and_3_cse
          , or_tmp_823 , return_add_generic_AC_RND_CONV_false_10_exp_and_5_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_tmp_im_d_1_sva_1_rsp_0 <= 7'b0000000;
    end
    else if ( rst ) begin
      stage_PE_1_tmp_im_d_1_sva_1_rsp_0 <= 7'b0000000;
    end
    else if ( stage_PE_1_tmp_im_d_and_ssc ) begin
      stage_PE_1_tmp_im_d_1_sva_1_rsp_0 <= MUX_v_7_2_2((out_f_d_rsci_q_d[63:57]),
          (in_f_d_rsci_q_d[63:57]), fsm_output[29]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_tmp_im_d_1_sva_1_rsp_1 <= 57'b000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      stage_PE_1_tmp_im_d_1_sva_1_rsp_1 <= 57'b000000000000000000000000000000000000000000000000000000000;
    end
    else if ( stage_PE_1_tmp_im_d_and_ssc & (~(or_dcpl_660 | (fsm_output[45]) | or_dcpl_985
        | (fsm_output[10]) | (fsm_output[34]) | (fsm_output[9]) | (fsm_output[35])
        | (fsm_output[19]))) ) begin
      stage_PE_1_tmp_im_d_1_sva_1_rsp_1 <= MUX1HOT_v_57_3_2((out_f_d_rsci_q_d[56:0]),
          z_out_30, (in_f_d_rsci_q_d[56:0]), {(fsm_output[4]) , stage_PE_1_tmp_im_d_or_1_nl
          , (fsm_output[29])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_0 <= 6'b000000;
    end
    else if ( rst ) begin
      stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_0 <= 6'b000000;
    end
    else if ( stage_PE_1_tmp_re_d_and_ssc & stage_PE_1_tmp_re_d_or_6_cse ) begin
      stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_0 <= MUX1HOT_v_6_3_2((z_out_30[56:51]),
          (out_f_d_rsci_q_d[56:51]), (in_f_d_rsci_q_d[56:51]), {stage_PE_1_tmp_re_d_or_4_rgt
          , stage_PE_1_tmp_re_d_and_5_rgt , stage_PE_1_tmp_re_d_and_7_rgt});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_1 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( rst ) begin
      stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_1 <= 51'b000000000000000000000000000000000000000000000000000;
    end
    else if ( stage_PE_1_tmp_re_d_and_ssc & (~(return_add_generic_AC_RND_CONV_false_17_e_r_and_cse
        | or_dcpl_418)) & stage_PE_1_tmp_re_d_or_6_cse ) begin
      stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_1 <= MUX1HOT_v_51_5_2((z_out_30[50:0]),
          (out_f_d_rsci_q_d[50:0]), stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0w0, stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx0w3,
          (in_f_d_rsci_q_d[50:0]), {stage_PE_1_tmp_re_d_or_4_rgt , stage_PE_1_tmp_re_d_and_5_rgt
          , stage_PE_1_tmp_re_d_and_3_nl , or_tmp_570 , stage_PE_1_tmp_re_d_and_7_rgt});
    end
  end
  assign nl_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_acc_nl = return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3
      + 11'b00000000001;
  assign return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_acc_nl = nl_return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_acc_nl[10:0];
  assign return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl = (~ return_mult_generic_AC_RND_CONV_false_6_e_incr_lpi_2_dfm_2)
      & return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1;
  assign return_mult_generic_AC_RND_CONV_false_6_else_2_else_mux_nl = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_6_exp_plus_1_acc_nl,
      return_mult_generic_AC_RND_CONV_false_6_exp_1_10_0_lpi_2_dfm_3, return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl);
  assign return_mult_generic_AC_RND_CONV_false_6_else_2_else_return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl
      = MUX_v_11_2_2(11'b00000000000, return_mult_generic_AC_RND_CONV_false_6_else_2_else_mux_nl,
      return_mult_generic_AC_RND_CONV_false_6_zero_m_return_mult_generic_AC_RND_CONV_false_6_zero_m_oelse_return_mult_generic_AC_RND_CONV_false_6_r_zero_return_extract_64_nand_mdf_sva_1);
  assign return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_or_nl
      = MUX_v_11_2_2(return_mult_generic_AC_RND_CONV_false_6_else_2_else_return_mult_generic_AC_RND_CONV_false_6_else_2_else_and_nl,
      11'b11111111111, return_mult_generic_AC_RND_CONV_false_6_lor_lpi_2_dfm_1);
  assign BUTTERFLY_if_1_and_nl = (~ return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1)
      & out1_rsci_idat_63_0_mx0c1;
  assign BUTTERFLY_if_1_and_1_nl = return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1
      & out1_rsci_idat_63_0_mx0c1;
  assign return_mult_generic_AC_RND_CONV_false_6_oelse_3_not_1_nl = ~ return_mult_generic_AC_RND_CONV_false_6_lor_3_lpi_2_dfm_1;
  assign return_mult_generic_AC_RND_CONV_false_6_return_mult_generic_AC_RND_CONV_false_6_and_1_nl
      = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000, (z_out_6[50:0]),
      return_mult_generic_AC_RND_CONV_false_6_oelse_3_not_1_nl);
  assign or_1606_nl = (fsm_output[42]) | (fsm_output[36]) | or_dcpl_712;
  assign stage_PE_qif_qelse_or_nl = (stage_PE_1_and_cse & (fsm_output[2])) | or_tmp_208;
  assign stage_PE_qif_qelse_mux_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_10, t_in_10_0_lpi_1_dfm_1_9,
      mode_lpi_1_dfm);
  assign stage_PE_qif_qelse_mux_1_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_13, m_in_15_1_lpi_1_dfm_1_14,
      mode_lpi_1_dfm);
  assign stage_PE_qif_qelse_mux_14_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_12, m_in_15_1_lpi_1_dfm_1_13,
      mode_lpi_1_dfm);
  assign stage_PE_qif_qelse_mux_13_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_11, m_in_15_1_lpi_1_dfm_1_12,
      mode_lpi_1_dfm);
  assign stage_PE_qif_qelse_mux_12_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_10, m_in_15_1_lpi_1_dfm_1_11,
      mode_lpi_1_dfm);
  assign stage_PE_qif_qelse_mux_11_nl = MUX_s_1_2_2(m_in_15_1_lpi_1_dfm_1_9, m_in_15_1_lpi_1_dfm_1_10,
      mode_lpi_1_dfm);
  assign BUTTERFLY_fry_BUTTERFLY_fry_mux_nl = MUX_v_10_2_2(z_out_2, (z_out_19[9:0]),
      fsm_output[55]);
  assign not_709_nl = ~ or_dcpl_395;
  assign return_extract_15_return_extract_15_nor_nl = ~((return_add_generic_AC_RND_CONV_false_4_e_r_qelse_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1);
  assign return_extract_47_return_extract_47_nor_nl = ~((return_add_generic_AC_RND_CONV_false_17_e_r_qelse_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm_1);
  assign return_add_generic_AC_RND_CONV_false_17_e_r_and_1_nl = inverse_lpi_1_dfm_1
      & or_dcpl_548;
  assign return_extract_20_m_zero_return_extract_20_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_11_mux_2_itm_mx3
      | (return_mult_generic_AC_RND_CONV_false_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_25_m_zero_return_extract_25_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_54_m_zero_return_extract_54_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_11_mux_2_itm_mx9
      | (return_mult_generic_AC_RND_CONV_false_4_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign operator_11_true_15_operator_11_true_15_and_nl = (return_add_generic_AC_RND_CONV_false_4_e_r_qelse_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1;
  assign operator_11_true_21_operator_11_true_21_and_nl = (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1==11'b11111111111);
  assign operator_11_true_27_operator_11_true_27_and_nl = (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1;
  assign operator_11_true_53_operator_11_true_53_and_nl = (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1==11'b11111111111);
  assign operator_11_true_59_operator_11_true_59_and_nl = (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_3_nl
      = return_add_generic_AC_RND_CONV_false_11_mux_2_itm_mx3 | return_add_generic_AC_RND_CONV_false_7_return_add_generic_AC_RND_CONV_false_7_or_tmp;
  assign return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_3_nl
      = drf_qr_lval_14_smx_0_lpi_3_dfm_mx3 | return_add_generic_AC_RND_CONV_false_20_return_add_generic_AC_RND_CONV_false_20_or_tmp;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_5_nl = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_7_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_11_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_8_nl = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_7_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_11_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_or_10_nl = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_16_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_or_nl = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_7_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_10_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_or_5_nl = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_8_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_9_cse | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_12_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_13_cse | return_add_generic_AC_RND_CONV_false_11_op_smaller_and_6_cse;
  assign return_add_generic_AC_RND_CONV_false_11_op_smaller_or_6_nl = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_11_cse
      | return_add_generic_AC_RND_CONV_false_11_op_bigger_and_14_cse;
  assign return_add_generic_AC_RND_CONV_false_11_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_11_e_dif_qr_lpi_3_dfm_mx0_10_0[10:6]!=5'b00000)
      | return_add_generic_AC_RND_CONV_false_9_e_dif_qelse_return_add_generic_AC_RND_CONV_false_9_e_dif_qelse_and_cse;
  assign return_add_generic_AC_RND_CONV_false_11_e_dif_sat_or_nl = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_11_e_dif_qr_lpi_3_dfm_mx0_10_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_11_e_dif_sat_or_1_nl);
  assign return_extract_15_return_extract_15_or_1_nl = (return_add_generic_AC_RND_CONV_false_4_e_r_qelse_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_4_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_2_nl
      = drf_qr_lval_14_smx_0_lpi_3_dfm_mx1 | return_add_generic_AC_RND_CONV_false_8_return_add_generic_AC_RND_CONV_false_8_or_tmp;
  assign return_extract_47_return_extract_47_or_1_nl = (return_add_generic_AC_RND_CONV_false_17_e_r_qelse_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_17_if_2_return_add_generic_AC_RND_CONV_false_17_if_2_nor_1_nl
      = ~(inverse_lpi_1_dfm_1 | (~ (O_1_out[63])));
  assign return_add_generic_AC_RND_CONV_false_17_and_1_nl = (~ or_dcpl_549) & return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  assign return_add_generic_AC_RND_CONV_false_17_and_7_nl = (~ or_590_cse) & return_add_generic_AC_RND_CONV_false_17_and_2_m1c;
  assign return_add_generic_AC_RND_CONV_false_17_and_8_nl = or_590_cse & return_add_generic_AC_RND_CONV_false_17_and_2_m1c;
  assign return_add_generic_AC_RND_CONV_false_18_if_2_return_add_generic_AC_RND_CONV_false_18_if_2_and_2_nl
      = inverse_lpi_1_dfm_1 & (O_1_out[63]);
  assign return_add_generic_AC_RND_CONV_false_18_r_sign_mux_1_nl = MUX_s_1_2_2((O_1_out[63]),
      inverse_lpi_1_dfm_1, or_590_cse);
  assign return_add_generic_AC_RND_CONV_false_5_do_sub_return_add_generic_AC_RND_CONV_false_5_do_sub_xor_nl
      = (O_1_out[63]) ^ inverse_lpi_1_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_10_do_sub_return_add_generic_AC_RND_CONV_false_10_do_sub_xor_nl
      = (stage_PE_1_x_im_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva_mx1;
  assign return_add_generic_AC_RND_CONV_false_23_do_sub_return_add_generic_AC_RND_CONV_false_23_do_sub_xor_nl
      = (stage_PE_1_x_im_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva_mx2;
  assign return_extract_18_and_nl = return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_if_1_return_add_generic_AC_RND_CONV_false_4_op2_normal_return_extract_9_nor_tmp
      & (O_1_out_1[51:0]==52'b0000000000000000000000000000000000000000000000000000);
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_or_10_nl = return_add_generic_AC_RND_CONV_false_13_op2_mu_or_3_rgt
      | (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_1_op_bigger_return_add_generic_AC_RND_CONV_false_13_op2_mu_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_1_op1_smaller_oelse_and_1_cse
      | (z_out_25[11]) | (~ inverse_lpi_1_dfm_1));
  assign return_add_generic_AC_RND_CONV_false_13_op2_mu_or_nl = (return_add_generic_AC_RND_CONV_false_13_return_add_generic_AC_RND_CONV_false_13_or_1_tmp
      & (~ inverse_lpi_1_dfm_1)) | return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx6c1
      | return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_mx6c2;
  assign return_add_generic_AC_RND_CONV_false_14_op_bigger_return_add_generic_AC_RND_CONV_false_13_op2_mu_nor_nl
      = ~(return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_return_add_generic_AC_RND_CONV_false_14_op1_smaller_oelse_and_1_cse
      | (z_out_25[11]) | (~ inverse_lpi_1_dfm_1));
  assign reg_return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm_rgt_nl
      = MUX1HOT_s_1_4_2(return_add_generic_AC_RND_CONV_false_1_op_bigger_return_add_generic_AC_RND_CONV_false_13_op2_mu_nor_nl,
      return_add_generic_AC_RND_CONV_false_13_op2_mu_or_nl, inverse_lpi_1_dfm_1,
      return_add_generic_AC_RND_CONV_false_14_op_bigger_return_add_generic_AC_RND_CONV_false_13_op2_mu_nor_nl,
      {(fsm_output[7]) , (fsm_output[30]) , (fsm_output[31]) , (fsm_output[32])});
  assign return_extract_22_m_zero_return_extract_22_m_zero_nor_nl = ~(drf_qr_lval_14_smx_0_lpi_3_dfm_mx1
      | (return_mult_generic_AC_RND_CONV_false_1_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_53_m_zero_return_extract_53_m_zero_nor_nl = ~(return_mult_generic_AC_RND_CONV_false_5_m_r_51_lpi_3_dfm_mx1
      | (return_mult_generic_AC_RND_CONV_false_5_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_59_m_zero_return_extract_59_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_21_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign operator_11_true_20_operator_11_true_20_and_nl = (return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_3_10_0_1==11'b11111111111);
  assign operator_11_true_25_operator_11_true_25_and_nl = (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_12_r_nan_and_nl = return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva & return_add_generic_AC_RND_CONV_false_12_do_sub_sva;
  assign operator_11_true_52_operator_11_true_52_and_nl = (return_mult_generic_AC_RND_CONV_false_3_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w6==11'b11111111111);
  assign operator_11_true_57_operator_11_true_57_and_nl = (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1;
  assign return_add_generic_AC_RND_CONV_false_25_r_nan_and_nl = return_add_generic_AC_RND_CONV_false_23_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_14_op2_inf_sva & return_add_generic_AC_RND_CONV_false_12_do_sub_sva;
  assign return_extract_21_m_zero_return_extract_21_m_zero_nor_nl = ~(return_mult_generic_AC_RND_CONV_false_2_m_r_51_lpi_3_dfm_mx1
      | (return_mult_generic_AC_RND_CONV_false_2_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_27_m_zero_return_extract_27_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_8_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_17_m_zero_or_2_nl = (fsm_output[29]) | or_200_cse;
  assign return_extract_17_m_zero_mux_nl = MUX_s_1_2_2((~ inverse_lpi_1_dfm_1), inverse_lpi_1_dfm_1,
      fsm_output[32]);
  assign operator_11_true_22_operator_11_true_22_and_nl = (return_mult_generic_AC_RND_CONV_false_1_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w3==11'b11111111111);
  assign operator_11_true_47_operator_11_true_47_and_nl = (return_add_generic_AC_RND_CONV_false_17_e_r_qelse_qr_10_1_lpi_3_dfm_1==10'b1111111111)
      & return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm_1;
  assign operator_11_true_54_operator_11_true_54_and_nl = (return_mult_generic_AC_RND_CONV_false_4_exp_1_11_0_lpi_3_dfm_3_10_0_mx0w2==11'b11111111111);
  assign return_extract_17_return_extract_17_or_1_nl = (return_add_generic_AC_RND_CONV_false_5_e_r_qelse_qr_10_1_lpi_3_dfm_1!=10'b0000000000)
      | return_add_generic_AC_RND_CONV_false_5_e_r_qr_0_lpi_3_dfm_1;
  assign or_1586_nl = (fsm_output[31]) | (fsm_output[29]);
  assign return_extract_52_m_zero_return_extract_52_m_zero_nor_nl = ~(drf_qr_lval_14_smx_0_lpi_3_dfm_mx3
      | (return_mult_generic_AC_RND_CONV_false_3_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_extract_57_m_zero_return_extract_57_m_zero_nor_nl = ~(return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0
      | (return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1!=51'b000000000000000000000000000000000000000000000000000));
  assign return_add_generic_AC_RND_CONV_false_11_and_7_nl = (~ return_add_generic_AC_RND_CONV_false_16_do_sub_sva)
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_11_and_8_nl = return_add_generic_AC_RND_CONV_false_16_do_sub_sva
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_11_and_9_nl = (~ return_add_generic_AC_RND_CONV_false_14_op2_nan_sva)
      & (fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_11_and_10_nl = return_add_generic_AC_RND_CONV_false_14_op2_nan_sva
      & (fsm_output[16]);
  assign return_add_generic_AC_RND_CONV_false_11_and_11_nl = (~ return_add_generic_AC_RND_CONV_false_11_do_sub_sva)
      & (fsm_output[17]);
  assign return_add_generic_AC_RND_CONV_false_11_and_12_nl = return_add_generic_AC_RND_CONV_false_11_do_sub_sva
      & (fsm_output[17]);
  assign return_add_generic_AC_RND_CONV_false_11_and_17_nl = (~ return_add_generic_AC_RND_CONV_false_16_do_sub_sva)
      & (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_11_and_18_nl = return_add_generic_AC_RND_CONV_false_16_do_sub_sva
      & (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_11_and_19_nl = (~ return_add_generic_AC_RND_CONV_false_11_do_sub_sva)
      & (fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_11_and_20_nl = return_add_generic_AC_RND_CONV_false_11_do_sub_sva
      & (fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_11_and_21_nl = (~ return_add_generic_AC_RND_CONV_false_14_op2_nan_sva)
      & (fsm_output[42]);
  assign return_add_generic_AC_RND_CONV_false_11_and_22_nl = return_add_generic_AC_RND_CONV_false_14_op2_nan_sva
      & (fsm_output[42]);
  assign return_add_generic_AC_RND_CONV_false_13_or_nl = (fsm_output[5]) | (fsm_output[19])
      | (fsm_output[21]) | (fsm_output[23]) | (fsm_output[25]) | (fsm_output[30])
      | (fsm_output[44]) | (fsm_output[46]) | (fsm_output[48]) | (fsm_output[50]);
  assign return_add_generic_AC_RND_CONV_false_2_if_2_return_add_generic_AC_RND_CONV_false_2_if_2_nor_1_nl
      = ~((stage_PE_1_tmp_im_d_1_sva_1_rsp_0[6]) | (~ (out_f_d_rsci_q_d[63])));
  assign return_add_generic_AC_RND_CONV_false_15_if_2_return_add_generic_AC_RND_CONV_false_15_if_2_nor_1_nl
      = ~((stage_PE_1_tmp_im_d_1_sva_1_rsp_0[6]) | (~ (in_f_d_rsci_q_d[63])));
  assign return_add_generic_AC_RND_CONV_false_11_or_nl = return_add_generic_AC_RND_CONV_false_11_and_32_cse
      | (return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse
      & return_add_generic_AC_RND_CONV_false_11_and_28_m1c);
  assign return_add_generic_AC_RND_CONV_false_11_and_27_nl = (~ or_dcpl_876) & (fsm_output[30]);
  assign return_add_generic_AC_RND_CONV_false_11_and_35_nl = (~ return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse)
      & return_add_generic_AC_RND_CONV_false_11_and_28_m1c;
  assign return_add_generic_AC_RND_CONV_false_2_do_sub_return_add_generic_AC_RND_CONV_false_2_do_sub_return_add_generic_AC_RND_CONV_false_2_do_sub_xnor_nl
      = ~((out_f_d_rsci_q_d[63]) ^ (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[6]));
  assign return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_return_add_generic_AC_RND_CONV_false_11_do_sub_xnor_nl
      = ~((stage_PE_1_x_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1);
  assign return_add_generic_AC_RND_CONV_false_15_do_sub_return_add_generic_AC_RND_CONV_false_15_do_sub_return_add_generic_AC_RND_CONV_false_15_do_sub_xnor_nl
      = ~((in_f_d_rsci_q_d[63]) ^ (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[6]));
  assign return_add_generic_AC_RND_CONV_false_22_do_sub_return_add_generic_AC_RND_CONV_false_22_do_sub_xor_nl
      = (stage_PE_1_x_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2;
  assign return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_return_add_generic_AC_RND_CONV_false_12_do_sub_xnor_nl
      = ~((stage_PE_1_x_im_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva_mx1);
  assign return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_return_add_generic_AC_RND_CONV_false_25_do_sub_xnor_nl
      = ~((stage_PE_1_x_im_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_19_return_add_generic_AC_RND_CONV_false_19_if_return_add_generic_AC_RND_CONV_false_19_op1_normal_return_extract_44_nor_cse_sva_mx2);
  assign return_add_generic_AC_RND_CONV_false_10_or_3_nl = or_dcpl_401 | return_add_generic_AC_RND_CONV_false_10_or_cse;
  assign return_add_generic_AC_RND_CONV_false_if_2_return_add_generic_AC_RND_CONV_false_if_2_and_2_nl
      = (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[6]) & (out_f_d_rsci_q_d[63]);
  assign return_add_generic_AC_RND_CONV_false_1_if_2_return_add_generic_AC_RND_CONV_false_1_if_2_and_2_nl
      = (out_f_d_rsci_q_d[63]) & (stage_PE_1_x_im_d_sva[63]);
  assign return_add_generic_AC_RND_CONV_false_13_if_2_return_add_generic_AC_RND_CONV_false_13_if_2_and_2_nl
      = (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[6]) & (in_f_d_rsci_q_d[63]);
  assign return_add_generic_AC_RND_CONV_false_14_if_2_return_add_generic_AC_RND_CONV_false_14_if_2_and_2_nl
      = (in_f_d_rsci_q_d[63]) & (stage_PE_1_x_im_d_sva[63]);
  assign return_extract_26_exception_or_nl = return_add_generic_AC_RND_CONV_false_11_and_31_cse
      | (return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse
      & return_extract_26_exception_and_5_m1c);
  assign return_extract_26_exception_or_4_nl = return_add_generic_AC_RND_CONV_false_11_and_32_cse
      | (return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse
      & and_494_m1c & (fsm_output[30]));
  assign return_extract_26_exception_and_4_nl = (~ and_491_tmp) & (fsm_output[7]);
  assign return_extract_26_exception_or_5_nl = ((~ return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse)
      & return_extract_26_exception_and_5_m1c) | return_extract_26_exception_and_17_cse
      | ((~ return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse)
      & return_extract_26_exception_and_10_m1c);
  assign return_extract_26_exception_and_8_nl = (~ inverse_lpi_1_dfm_1) & (fsm_output[30]);
  assign and_493_nl = return_add_generic_AC_RND_CONV_false_15_aif_equal_tmp & return_add_generic_AC_RND_CONV_false_13_e1_eq_e2_equal_tmp
      & inverse_lpi_1_dfm_1 & (fsm_output[30]);
  assign return_extract_26_exception_or_6_nl = ((~ return_add_generic_AC_RND_CONV_false_15_op1_smaller_return_add_generic_AC_RND_CONV_false_15_op1_smaller_or_cse)
      & and_494_m1c & (fsm_output[30])) | (return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse
      & return_extract_26_exception_and_10_m1c);
  assign return_extract_26_exception_and_9_nl = (~ and_497_tmp) & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_10_or_4_nl = (inverse_lpi_1_dfm_1 &
      (fsm_output[5])) | (fsm_output[19]) | (fsm_output[21]) | (fsm_output[23]) |
      (fsm_output[25]) | (fsm_output[30]) | (fsm_output[44]) | (fsm_output[46]) |
      (fsm_output[48]) | (fsm_output[50]);
  assign and_498_nl = (~ inverse_lpi_1_dfm_1) & return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp
      & (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_10_and_4_nl = (~(inverse_lpi_1_dfm_1
      | return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp))
      & (fsm_output[5]);
  assign return_add_generic_AC_RND_CONV_false_3_r_nan_and_nl = return_add_generic_AC_RND_CONV_false_10_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva & return_add_generic_AC_RND_CONV_false_16_do_sub_sva;
  assign return_add_generic_AC_RND_CONV_false_16_r_nan_and_nl = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_14_op2_inf_sva & return_add_generic_AC_RND_CONV_false_16_do_sub_sva;
  assign return_add_generic_AC_RND_CONV_false_24_r_nan_and_nl = return_add_generic_AC_RND_CONV_false_22_op1_inf_sva
      & return_add_generic_AC_RND_CONV_false_10_op2_inf_sva & return_add_generic_AC_RND_CONV_false_14_op2_nan_sva;
  assign return_extract_58_and_2_nl = return_add_generic_AC_RND_CONV_false_11_mux_itm
      & (~ return_extract_26_m_zero_sva);
  assign return_extract_58_and_1_nl = return_add_generic_AC_RND_CONV_false_11_mux_itm
      & return_extract_26_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_9_do_sub_return_add_generic_AC_RND_CONV_false_9_do_sub_xor_nl
      = (stage_PE_1_x_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx1;
  assign return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_return_add_generic_AC_RND_CONV_false_24_do_sub_xnor_nl
      = ~((stage_PE_1_x_re_d_sva[63]) ^ return_add_generic_AC_RND_CONV_false_20_r_sign_lpi_3_dfm_1_mx2);
  assign return_add_generic_AC_RND_CONV_false_8_do_sub_return_add_generic_AC_RND_CONV_false_8_do_sub_xor_nl
      = stage_d_mul_return_d_4_63_sva_1 ^ stage_d_mul_return_d_2_63_sva_1;
  assign return_add_generic_AC_RND_CONV_false_21_do_sub_return_add_generic_AC_RND_CONV_false_21_do_sub_xor_nl
      = stage_d_mul_return_d_4_63_sva_1 ^ stage_d_mul_return_d_5_63_sva_1;
  assign return_add_generic_AC_RND_CONV_false_3_if_2_return_add_generic_AC_RND_CONV_false_3_if_2_nor_1_nl
      = ~((out_f_d_rsci_q_d[63]) | (~ (stage_PE_1_x_im_d_sva[63])));
  assign return_add_generic_AC_RND_CONV_false_16_if_2_return_add_generic_AC_RND_CONV_false_16_if_2_nor_1_nl
      = ~((in_f_d_rsci_q_d[63]) | (~ (stage_PE_1_x_im_d_sva[63])));
  assign return_add_generic_AC_RND_CONV_false_12_and_1_nl = (~ or_dcpl_911) & (fsm_output[7]);
  assign return_add_generic_AC_RND_CONV_false_12_or_nl = ((~ return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse)
      & return_add_generic_AC_RND_CONV_false_12_and_2_m1c) | return_extract_26_exception_and_17_cse
      | ((~ return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse)
      & return_add_generic_AC_RND_CONV_false_12_and_6_m1c);
  assign return_add_generic_AC_RND_CONV_false_12_and_10_nl = return_add_generic_AC_RND_CONV_false_3_op1_smaller_return_add_generic_AC_RND_CONV_false_3_op1_smaller_or_cse
      & return_add_generic_AC_RND_CONV_false_12_and_2_m1c;
  assign return_add_generic_AC_RND_CONV_false_12_and_5_nl = (~ or_dcpl_913) & (fsm_output[32]);
  assign return_add_generic_AC_RND_CONV_false_12_and_14_nl = return_add_generic_AC_RND_CONV_false_16_op1_smaller_return_add_generic_AC_RND_CONV_false_16_op1_smaller_or_cse
      & return_add_generic_AC_RND_CONV_false_12_and_6_m1c;
  assign return_add_generic_AC_RND_CONV_false_3_do_sub_return_add_generic_AC_RND_CONV_false_3_do_sub_return_add_generic_AC_RND_CONV_false_3_do_sub_xnor_nl
      = ~((stage_PE_1_x_im_d_sva[63]) ^ (out_f_d_rsci_q_d[63]));
  assign return_add_generic_AC_RND_CONV_false_7_do_sub_return_add_generic_AC_RND_CONV_false_7_do_sub_xor_nl
      = stage_d_mul_return_d_63_sva_1 ^ stage_d_mul_return_d_2_63_sva_1;
  assign return_add_generic_AC_RND_CONV_false_16_do_sub_return_add_generic_AC_RND_CONV_false_16_do_sub_return_add_generic_AC_RND_CONV_false_16_do_sub_xnor_nl
      = ~((stage_PE_1_x_im_d_sva[63]) ^ (in_f_d_rsci_q_d[63]));
  assign return_add_generic_AC_RND_CONV_false_20_do_sub_return_add_generic_AC_RND_CONV_false_20_do_sub_xor_nl
      = stage_d_mul_return_d_63_sva_1 ^ stage_d_mul_return_d_5_63_sva_1;
  assign return_extract_26_and_1_nl = operator_11_true_return_26_sva & return_extract_26_m_zero_sva;
  assign return_extract_26_and_2_nl = operator_11_true_return_26_sva & (~ return_extract_26_m_zero_sva);
  assign return_extract_56_and_2_nl = operator_11_true_return_26_sva & (~ return_extract_17_m_zero_sva);
  assign return_extract_56_and_1_nl = operator_11_true_return_26_sva & return_extract_17_m_zero_sva;
  assign return_add_generic_AC_RND_CONV_false_12_op_bigger_or_4_nl = return_add_generic_AC_RND_CONV_false_10_exp_and_3_cse
      | return_add_generic_AC_RND_CONV_false_10_exp_and_5_cse;
  assign return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_6_nl = MUX_s_1_2_2(and_dcpl_267,
      and_dcpl_268, fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_12_res_mant_return_add_generic_AC_RND_CONV_false_12_res_mant_return_add_generic_AC_RND_CONV_false_12_res_mant_or_nl
      = return_add_generic_AC_RND_CONV_false_11_op_bigger_and_16_cse | return_add_generic_AC_RND_CONV_false_11_exp_and_3_cse;
  assign return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_2_nl
      = return_add_generic_AC_RND_CONV_false_11_mux_2_itm_mx9 | return_add_generic_AC_RND_CONV_false_21_return_add_generic_AC_RND_CONV_false_21_or_tmp;
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_33_nl = (~ and_dcpl_260)
      & (fsm_output[14]);
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_and_35_nl = (~ and_dcpl_264)
      & (fsm_output[39]);
  assign return_add_generic_AC_RND_CONV_false_25_e_dif_sat_or_1_nl = (return_add_generic_AC_RND_CONV_false_25_e_dif_qr_lpi_3_dfm_mx0_10_0[10:6]!=5'b00000)
      | return_add_generic_AC_RND_CONV_false_9_e_dif_qelse_return_add_generic_AC_RND_CONV_false_9_e_dif_qelse_and_cse;
  assign return_add_generic_AC_RND_CONV_false_25_e_dif_sat_or_nl = MUX_v_6_2_2((return_add_generic_AC_RND_CONV_false_25_e_dif_qr_lpi_3_dfm_mx0_10_0[5:0]),
      6'b111111, return_add_generic_AC_RND_CONV_false_25_e_dif_sat_or_1_nl);
  assign BUTTERFLY_n_mux1h_1_nl = MUX1HOT_v_9_3_2((BUTTERFLY_1_fry_9_0_sva[8:0]),
      (BUTTERFLY_1_i_9_0_sva[8:0]), (BUTTERFLY_1_n_9_0_sva_1[8:0]), {BUTTERFLY_1_fiy_or_1_cse
      , or_tmp_234 , or_dcpl_395});
  assign BUTTERFLY_1_fiy_nand_nl = ~(nor_24_cse & (~((fsm_output[50]) | (fsm_output[46])))
      & (~((fsm_output[25]) | (fsm_output[42]))) & (~((fsm_output[21]) | (fsm_output[17]))));
  assign BUTTERFLY_n_and_nl = MUX_v_9_2_2(9'b000000000, BUTTERFLY_n_mux1h_1_nl, BUTTERFLY_1_fiy_nand_nl);
  assign or_1355_nl = or_dcpl_395 | (fsm_output[2]) | or_dcpl_106 | (fsm_output[25])
      | (fsm_output[42]) | (fsm_output[21]) | (fsm_output[17]);
  assign or_1996_nl = and_1608_cse | and_1598_cse;
  assign or_1998_nl = and_1163_cse | or_tmp_348;
  assign or_2005_nl = (or_1144_cse & (fsm_output[39])) | (return_add_generic_AC_RND_CONV_false_8_op1_smaller_return_add_generic_AC_RND_CONV_false_8_op1_smaller_or_cse
      & (fsm_output[14]));
  assign or_2010_nl = or_tmp_823 | and_2281_cse;
  assign stage_PE_1_tmp_im_d_or_1_nl = or_dcpl_571 | stage_PE_1_tmp_im_d_1_sva_1_mx0c3;
  assign stage_PE_1_tmp_re_d_and_3_nl = (~ or_tmp_570) & stage_PE_1_tmp_re_d_1_sva_1_mx0c4;
  assign operator_6_false_1_mux1h_9_nl = MUX1HOT_s_1_7_2(BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1,
      BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_1, drf_qr_lval_11_smx_lpi_3_dfm_10,
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd, (drf_qr_lval_13_smx_10_1_lpi_3_dfm[9]),
      (drf_qr_lval_14_smx_10_1_lpi_3_dfm[9]), (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[4]),
      {or_tmp_927 , operator_6_false_1_or_1_ssc , or_tmp_929 , operator_6_false_1_or_8_cse
      , or_dcpl_751 , operator_6_false_1_or_4_cse , operator_6_false_1_or_6_cse});
  assign operator_6_false_1_mux1h_10_nl = MUX1HOT_s_1_7_2((reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[4]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd, drf_qr_lval_11_smx_lpi_3_dfm_9,
      (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1[3]), (drf_qr_lval_13_smx_10_1_lpi_3_dfm[8]),
      (drf_qr_lval_14_smx_10_1_lpi_3_dfm[8]), (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[3]),
      {or_tmp_927 , operator_6_false_1_or_1_ssc , or_tmp_929 , operator_6_false_1_or_8_cse
      , or_dcpl_751 , operator_6_false_1_or_4_cse , operator_6_false_1_or_6_cse});
  assign operator_6_false_1_mux1h_11_nl = MUX1HOT_v_3_7_2((reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[3:1]),
      (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1[3:1]), (drf_qr_lval_11_smx_lpi_3_dfm_8_5[3:1]),
      (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1[2:0]), (drf_qr_lval_13_smx_10_1_lpi_3_dfm[7:5]),
      (drf_qr_lval_14_smx_10_1_lpi_3_dfm[7:5]), (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[2:0]),
      {or_tmp_927 , operator_6_false_1_or_1_ssc , or_tmp_929 , operator_6_false_1_or_8_cse
      , or_dcpl_751 , operator_6_false_1_or_4_cse , operator_6_false_1_or_6_cse});
  assign operator_6_false_1_mux1h_12_nl = MUX1HOT_s_1_7_2((reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[0]),
      (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1[0]), (drf_qr_lval_11_smx_lpi_3_dfm_8_5[0]),
      (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2[3]), (drf_qr_lval_13_smx_10_1_lpi_3_dfm[4]),
      (drf_qr_lval_14_smx_10_1_lpi_3_dfm[4]), (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[4]),
      {or_tmp_927 , operator_6_false_1_or_1_ssc , or_tmp_929 , operator_6_false_1_or_8_cse
      , or_dcpl_751 , operator_6_false_1_or_4_cse , operator_6_false_1_or_6_cse});
  assign operator_6_false_1_mux1h_13_nl = MUX1HOT_v_3_7_2((reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[4:2]),
      (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2[3:1]), (drf_qr_lval_11_smx_lpi_3_dfm_4_0[4:2]),
      (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2[2:0]), (drf_qr_lval_13_smx_10_1_lpi_3_dfm[3:1]),
      (drf_qr_lval_14_smx_10_1_lpi_3_dfm[3:1]), (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[3:1]),
      {or_tmp_927 , operator_6_false_1_or_1_ssc , or_tmp_929 , operator_6_false_1_or_8_cse
      , or_dcpl_751 , operator_6_false_1_or_4_cse , operator_6_false_1_or_6_cse});
  assign operator_6_false_1_mux1h_14_nl = MUX1HOT_s_1_7_2((reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[1]),
      (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2[0]), (drf_qr_lval_11_smx_lpi_3_dfm_4_0[1]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3, (drf_qr_lval_13_smx_10_1_lpi_3_dfm[0]),
      (drf_qr_lval_14_smx_10_1_lpi_3_dfm[0]), (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[0]),
      {or_tmp_927 , operator_6_false_1_or_1_ssc , or_tmp_929 , operator_6_false_1_or_8_cse
      , or_dcpl_751 , operator_6_false_1_or_4_cse , operator_6_false_1_or_6_cse});
  assign operator_6_false_1_or_16_nl = (fsm_output[22]) | (fsm_output[47]);
  assign operator_6_false_1_or_17_nl = (fsm_output[24]) | (fsm_output[49]);
  assign operator_6_false_1_or_18_nl = (fsm_output[26]) | (fsm_output[51]);
  assign operator_6_false_1_mux1h_15_nl = MUX1HOT_s_1_7_2((reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[0]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3, (drf_qr_lval_11_smx_lpi_3_dfm_4_0[0]),
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm, drf_qr_lval_13_smx_0_lpi_3_dfm,
      drf_qr_lval_14_smx_0_lpi_3_dfm, drf_qr_lval_15_smx_0_lpi_3_dfm, {or_tmp_927
      , operator_6_false_1_or_1_ssc , or_tmp_929 , return_add_generic_AC_RND_CONV_false_12_res_mant_or_cse
      , operator_6_false_1_or_16_nl , operator_6_false_1_or_17_nl , operator_6_false_1_or_18_nl});
  assign operator_6_false_1_or_19_nl = or_tmp_927 | or_tmp_929 | or_tmp_930 | (fsm_output[22])
      | (fsm_output[47]);
  assign operator_6_false_1_or_20_nl = or_dcpl_548 | (fsm_output[24]) | (fsm_output[45])
      | (fsm_output[51]);
  assign operator_6_false_1_or_21_nl = (fsm_output[20]) | (fsm_output[26]) | (fsm_output[49]);
  assign operator_6_false_1_mux1h_16_nl = MUX1HOT_v_6_3_2((~ return_add_generic_AC_RND_CONV_false_10_ls_sva),
      (~ return_add_generic_AC_RND_CONV_false_11_ls_sva), (~ return_add_generic_AC_RND_CONV_false_12_ls_sva),
      {operator_6_false_1_or_19_nl , operator_6_false_1_or_20_nl , operator_6_false_1_or_21_nl});
  assign nl_acc_1_nl = conv_u2u_12_13({operator_6_false_1_mux1h_9_nl , operator_6_false_1_mux1h_10_nl
      , operator_6_false_1_mux1h_11_nl , operator_6_false_1_mux1h_12_nl , operator_6_false_1_mux1h_13_nl
      , operator_6_false_1_mux1h_14_nl , operator_6_false_1_mux1h_15_nl , 1'b1})
      + conv_s2u_8_13({1'b1 , operator_6_false_1_mux1h_16_nl , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[12:0];
  assign z_out_1 = readslicef_13_12_1(acc_1_nl);
  assign BUTTERFLY_fry_mux_10_nl = MUX_s_1_2_2(stage_PE_1_qr_0_lpi_2_dfm, stage_PE_1_qr_10_1_lpi_2_dfm_8,
      or_tmp_940);
  assign BUTTERFLY_fry_mux_11_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_8, reg_stage_PE_1_qr_10_1_lpi_2_dfm_7_0_ftd,
      or_tmp_940);
  assign BUTTERFLY_fry_mux_12_nl = MUX_s_1_2_2(reg_stage_PE_1_qr_10_1_lpi_2_dfm_7_0_ftd,
      reg_stage_PE_1_qr_10_1_lpi_2_dfm_7_0_ftd_1, or_tmp_940);
  assign BUTTERFLY_fry_mux_13_nl = MUX_s_1_2_2(reg_stage_PE_1_qr_10_1_lpi_2_dfm_7_0_ftd_1,
      stage_PE_1_qr_10_1_lpi_2_dfm_5, or_tmp_940);
  assign BUTTERFLY_fry_mux_14_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_5, stage_PE_1_qr_10_1_lpi_2_dfm_4,
      or_tmp_940);
  assign BUTTERFLY_fry_mux_15_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_4, stage_PE_1_qr_10_1_lpi_2_dfm_3,
      or_tmp_940);
  assign BUTTERFLY_fry_mux_16_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_3, stage_PE_1_qr_10_1_lpi_2_dfm_2,
      or_tmp_940);
  assign BUTTERFLY_fry_mux_17_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_2, stage_PE_1_qr_10_1_lpi_2_dfm_1,
      or_tmp_940);
  assign BUTTERFLY_fry_mux_18_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_1, stage_PE_1_qr_10_1_lpi_2_dfm_0,
      or_tmp_940);
  assign BUTTERFLY_fry_mux_19_nl = MUX_s_1_2_2(stage_PE_1_qr_10_1_lpi_2_dfm_0, stage_PE_1_qr_0_lpi_2_dfm,
      or_tmp_940);
  assign nl_z_out_2 = BUTTERFLY_i_9_0_sva_1 + ({BUTTERFLY_fry_mux_10_nl , BUTTERFLY_fry_mux_11_nl
      , BUTTERFLY_fry_mux_12_nl , BUTTERFLY_fry_mux_13_nl , BUTTERFLY_fry_mux_14_nl
      , BUTTERFLY_fry_mux_15_nl , BUTTERFLY_fry_mux_16_nl , BUTTERFLY_fry_mux_17_nl
      , BUTTERFLY_fry_mux_18_nl , BUTTERFLY_fry_mux_19_nl});
  assign z_out_2 = nl_z_out_2[9:0];
  assign nl_z_out_3 = conv_s2u_17_18(z_out_40) + conv_u2u_14_18(signext_14_13({(z_out_40[16])
      , 11'b00000000000 , (z_out_40[16])}));
  assign z_out_3 = nl_z_out_3[17:0];
  assign nl_operator_32_false_acc_nl = conv_u2u_16_32(z_out_5) + conv_u2u_28_32({(~
      z_out_5) , 12'b000000000000}) + conv_u2u_30_32({z_out_5 , 14'b01000000000000})
      + (z_out_21[31:0]) + 32'b11110000000000000000000000000000;
  assign operator_32_false_acc_nl = nl_operator_32_false_acc_nl[31:0];
  assign z_out_4_31_16 = readslicef_32_16_16(operator_32_false_acc_nl);
  assign nl_z_out_5 = ({(z_out_19[3:0]) , 12'b000000000001}) + (~ (z_out_21[15:0]));
  assign z_out_5 = nl_z_out_5[15:0];
  assign return_add_generic_AC_RND_CONV_false_4_res_rounded_return_add_generic_AC_RND_CONV_false_4_res_rounded_and_1_nl
      = (z_out_15[56]) & (~((fsm_output[10]) | (fsm_output[12]) | (fsm_output[14])
      | (fsm_output[35]) | (fsm_output[37]) | (fsm_output[39]) | (fsm_output[54])));
  assign return_add_generic_AC_RND_CONV_false_4_res_rounded_mux1h_2_nl = MUX1HOT_v_52_8_2((z_out_15[55:4]),
      (return_mult_generic_AC_RND_CONV_false_res_bef_rnd_3_53_1_lpi_3_dfm_1[52:1]),
      (return_mult_generic_AC_RND_CONV_false_1_res_bef_rnd_3_53_1_lpi_3_dfm_1[52:1]),
      (return_mult_generic_AC_RND_CONV_false_2_res_bef_rnd_3_53_1_lpi_3_dfm_1[52:1]),
      (return_mult_generic_AC_RND_CONV_false_3_res_bef_rnd_3_53_1_lpi_3_dfm_1[52:1]),
      (return_mult_generic_AC_RND_CONV_false_4_res_bef_rnd_3_53_1_lpi_3_dfm_1[52:1]),
      (return_mult_generic_AC_RND_CONV_false_5_res_bef_rnd_3_53_1_lpi_3_dfm_1[52:1]),
      (return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1[52:1]),
      {return_add_generic_AC_RND_CONV_false_4_res_rounded_or_1_cse , (fsm_output[10])
      , (fsm_output[12]) , (fsm_output[14]) , (fsm_output[35]) , (fsm_output[37])
      , (fsm_output[39]) , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_4_res_rounded_and_1_nl = (z_out_15[3])
      & ((z_out_15[0]) | (z_out_15[1]) | (z_out_15[2]) | (z_out_15[4]));
  assign return_mult_generic_AC_RND_CONV_false_if_1_or_4_nl = (z_out_18[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_if_1_aelse_return_mult_generic_AC_RND_CONV_false_if_1_aelse_or_2
      & (z_out_18[51]));
  assign return_mult_generic_AC_RND_CONV_false_mux_14_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_if_1_or_4_nl,
      return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_or_cse,
      z_out_27[12]);
  assign return_mult_generic_AC_RND_CONV_false_and_3_nl = (return_mult_generic_AC_RND_CONV_false_res_bef_rnd_3_53_1_lpi_3_dfm_1[0])
      & (return_mult_generic_AC_RND_CONV_false_mux_14_nl | (return_mult_generic_AC_RND_CONV_false_res_bef_rnd_3_53_1_lpi_3_dfm_1[1]));
  assign return_mult_generic_AC_RND_CONV_false_1_if_1_or_1_nl = (z_out_18[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_return_mult_generic_AC_RND_CONV_false_1_if_1_aelse_or_2
      & (z_out_18[51]));
  assign return_mult_generic_AC_RND_CONV_false_1_mux_14_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_1_if_1_or_1_nl,
      return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_or_cse,
      z_out_27[12]);
  assign return_mult_generic_AC_RND_CONV_false_1_and_3_nl = (return_mult_generic_AC_RND_CONV_false_1_res_bef_rnd_3_53_1_lpi_3_dfm_1[0])
      & (return_mult_generic_AC_RND_CONV_false_1_mux_14_nl | (return_mult_generic_AC_RND_CONV_false_1_res_bef_rnd_3_53_1_lpi_3_dfm_1[1]));
  assign return_mult_generic_AC_RND_CONV_false_2_if_1_or_1_nl = (z_out_18[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_return_mult_generic_AC_RND_CONV_false_2_if_1_aelse_or_2
      & (z_out_18[51]));
  assign return_mult_generic_AC_RND_CONV_false_2_mux_14_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_2_if_1_or_1_nl,
      return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_or_cse,
      z_out_27[12]);
  assign return_mult_generic_AC_RND_CONV_false_2_and_3_nl = (return_mult_generic_AC_RND_CONV_false_2_res_bef_rnd_3_53_1_lpi_3_dfm_1[0])
      & (return_mult_generic_AC_RND_CONV_false_2_mux_14_nl | (return_mult_generic_AC_RND_CONV_false_2_res_bef_rnd_3_53_1_lpi_3_dfm_1[1]));
  assign return_mult_generic_AC_RND_CONV_false_3_if_1_or_1_nl = (z_out_18[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_3_if_1_aelse_return_mult_generic_AC_RND_CONV_false_3_if_1_aelse_or_2
      & (z_out_18[51]));
  assign return_mult_generic_AC_RND_CONV_false_3_mux_14_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_3_if_1_or_1_nl,
      return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_or_cse,
      z_out_27[12]);
  assign return_mult_generic_AC_RND_CONV_false_3_and_3_nl = (return_mult_generic_AC_RND_CONV_false_3_res_bef_rnd_3_53_1_lpi_3_dfm_1[0])
      & (return_mult_generic_AC_RND_CONV_false_3_mux_14_nl | (return_mult_generic_AC_RND_CONV_false_3_res_bef_rnd_3_53_1_lpi_3_dfm_1[1]));
  assign return_mult_generic_AC_RND_CONV_false_4_if_1_or_1_nl = (z_out_18[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_return_mult_generic_AC_RND_CONV_false_4_if_1_aelse_or_2
      & (z_out_18[51]));
  assign return_mult_generic_AC_RND_CONV_false_4_mux_14_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_4_if_1_or_1_nl,
      return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_or_cse,
      z_out_27[12]);
  assign return_mult_generic_AC_RND_CONV_false_4_and_3_nl = (return_mult_generic_AC_RND_CONV_false_4_res_bef_rnd_3_53_1_lpi_3_dfm_1[0])
      & (return_mult_generic_AC_RND_CONV_false_4_mux_14_nl | (return_mult_generic_AC_RND_CONV_false_4_res_bef_rnd_3_53_1_lpi_3_dfm_1[1]));
  assign return_mult_generic_AC_RND_CONV_false_5_if_1_or_1_nl = (z_out_18[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_return_mult_generic_AC_RND_CONV_false_5_if_1_aelse_or_2
      & (z_out_18[51]));
  assign return_mult_generic_AC_RND_CONV_false_5_mux_14_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_5_if_1_or_1_nl,
      return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_else_1_sticky_bit_or_cse,
      z_out_27[12]);
  assign return_mult_generic_AC_RND_CONV_false_5_and_3_nl = (return_mult_generic_AC_RND_CONV_false_5_res_bef_rnd_3_53_1_lpi_3_dfm_1[0])
      & (return_mult_generic_AC_RND_CONV_false_5_mux_14_nl | (return_mult_generic_AC_RND_CONV_false_5_res_bef_rnd_3_53_1_lpi_3_dfm_1[1]));
  assign return_mult_generic_AC_RND_CONV_false_6_if_1_or_1_nl = (z_out_18[50:0]!=51'b000000000000000000000000000000000000000000000000000)
      | (return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_return_mult_generic_AC_RND_CONV_false_6_if_1_aelse_or_2
      & (z_out_18[51]));
  assign return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_or_1_nl
      = (return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp
      & (~ (z_out_17[51]))) | ((out_f_d_rsci_q_d[51]) & (~ (z_out_17[50]))) | ((out_f_d_rsci_q_d[50])
      & (~ (z_out_17[49]))) | ((out_f_d_rsci_q_d[49]) & (~ (z_out_17[48]))) | ((out_f_d_rsci_q_d[48])
      & (~ (z_out_17[47]))) | ((out_f_d_rsci_q_d[47]) & (~ (z_out_17[46]))) | ((out_f_d_rsci_q_d[46])
      & (~ (z_out_17[45]))) | ((out_f_d_rsci_q_d[45]) & (~ (z_out_17[44]))) | ((out_f_d_rsci_q_d[44])
      & (~ (z_out_17[43]))) | ((out_f_d_rsci_q_d[43]) & (~ (z_out_17[42]))) | ((out_f_d_rsci_q_d[42])
      & (~ (z_out_17[41]))) | ((out_f_d_rsci_q_d[41]) & (~ (z_out_17[40]))) | ((out_f_d_rsci_q_d[40])
      & (~ (z_out_17[39]))) | ((out_f_d_rsci_q_d[39]) & (~ (z_out_17[38]))) | ((out_f_d_rsci_q_d[38])
      & (~ (z_out_17[37]))) | ((out_f_d_rsci_q_d[37]) & (~ (z_out_17[36]))) | ((out_f_d_rsci_q_d[36])
      & (~ (z_out_17[35]))) | ((out_f_d_rsci_q_d[35]) & (~ (z_out_17[34]))) | ((out_f_d_rsci_q_d[34])
      & (~ (z_out_17[33]))) | ((out_f_d_rsci_q_d[33]) & (~ (z_out_17[32]))) | ((out_f_d_rsci_q_d[32])
      & (~ (z_out_17[31]))) | ((out_f_d_rsci_q_d[31]) & (~ (z_out_17[30]))) | ((out_f_d_rsci_q_d[30])
      & (~ (z_out_17[29]))) | ((out_f_d_rsci_q_d[29]) & (~ (z_out_17[28]))) | ((out_f_d_rsci_q_d[28])
      & (~ (z_out_17[27]))) | ((out_f_d_rsci_q_d[27]) & (~ (z_out_17[26]))) | ((out_f_d_rsci_q_d[26])
      & (~ (z_out_17[25]))) | ((out_f_d_rsci_q_d[25]) & (~ (z_out_17[24]))) | ((out_f_d_rsci_q_d[24])
      & (~ (z_out_17[23]))) | ((out_f_d_rsci_q_d[23]) & (~ (z_out_17[22]))) | ((out_f_d_rsci_q_d[22])
      & (~ (z_out_17[21]))) | ((out_f_d_rsci_q_d[21]) & (~ (z_out_17[20]))) | ((out_f_d_rsci_q_d[20])
      & (~ (z_out_17[19]))) | ((out_f_d_rsci_q_d[19]) & (~ (z_out_17[18]))) | ((out_f_d_rsci_q_d[18])
      & (~ (z_out_17[17]))) | ((out_f_d_rsci_q_d[17]) & (~ (z_out_17[16]))) | ((out_f_d_rsci_q_d[16])
      & (~ (z_out_17[15]))) | ((out_f_d_rsci_q_d[15]) & (~ (z_out_17[14]))) | ((out_f_d_rsci_q_d[14])
      & (~ (z_out_17[13]))) | ((out_f_d_rsci_q_d[13]) & (~ (z_out_17[12]))) | ((out_f_d_rsci_q_d[12])
      & (~ (z_out_17[11]))) | ((out_f_d_rsci_q_d[11]) & (~ (z_out_17[10]))) | ((out_f_d_rsci_q_d[10])
      & (~ (z_out_17[9]))) | ((out_f_d_rsci_q_d[9]) & (~ (z_out_17[8]))) | ((out_f_d_rsci_q_d[8])
      & (~ (z_out_17[7]))) | ((out_f_d_rsci_q_d[7]) & (~ (z_out_17[6]))) | ((out_f_d_rsci_q_d[6])
      & (~ (z_out_17[5]))) | ((out_f_d_rsci_q_d[5]) & (~ (z_out_17[4]))) | ((out_f_d_rsci_q_d[4])
      & (~ (z_out_17[3]))) | ((out_f_d_rsci_q_d[3]) & (~ (z_out_17[2]))) | ((out_f_d_rsci_q_d[2])
      & (~ (z_out_17[1]))) | ((out_f_d_rsci_q_d[1]) & (~ (z_out_17[0]))) | (out_f_d_rsci_q_d[0]);
  assign return_mult_generic_AC_RND_CONV_false_6_mux_12_nl = MUX_s_1_2_2(return_mult_generic_AC_RND_CONV_false_6_if_1_or_1_nl,
      return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_return_mult_generic_AC_RND_CONV_false_6_else_1_sticky_bit_or_1_nl,
      z_out_27[11]);
  assign return_mult_generic_AC_RND_CONV_false_6_and_3_nl = (return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1[0])
      & (return_mult_generic_AC_RND_CONV_false_6_mux_12_nl | (return_mult_generic_AC_RND_CONV_false_6_res_bef_rnd_3_53_1_lpi_2_dfm_1[1]));
  assign return_add_generic_AC_RND_CONV_false_4_res_rounded_mux1h_3_nl = MUX1HOT_s_1_8_2(return_add_generic_AC_RND_CONV_false_4_res_rounded_and_1_nl,
      return_mult_generic_AC_RND_CONV_false_and_3_nl, return_mult_generic_AC_RND_CONV_false_1_and_3_nl,
      return_mult_generic_AC_RND_CONV_false_2_and_3_nl, return_mult_generic_AC_RND_CONV_false_3_and_3_nl,
      return_mult_generic_AC_RND_CONV_false_4_and_3_nl, return_mult_generic_AC_RND_CONV_false_5_and_3_nl,
      return_mult_generic_AC_RND_CONV_false_6_and_3_nl, {return_add_generic_AC_RND_CONV_false_4_res_rounded_or_1_cse
      , (fsm_output[10]) , (fsm_output[12]) , (fsm_output[14]) , (fsm_output[35])
      , (fsm_output[37]) , (fsm_output[39]) , (fsm_output[54])});
  assign nl_z_out_6 = conv_u2u_53_54({return_add_generic_AC_RND_CONV_false_4_res_rounded_return_add_generic_AC_RND_CONV_false_4_res_rounded_and_1_nl
      , return_add_generic_AC_RND_CONV_false_4_res_rounded_mux1h_2_nl}) + conv_u2u_1_54(return_add_generic_AC_RND_CONV_false_4_res_rounded_mux1h_3_nl);
  assign z_out_6 = nl_z_out_6[53:0];
  assign stage_PE_stage_PE_stage_PE_mux_3_nl = MUX_s_1_2_2(t_in_10_0_lpi_1_dfm_1_10,
      t_in_10_0_lpi_1_dfm_1_9, return_extract_26_m_zero_sva);
  assign BUTTERFLY_if_mux_14_nl = MUX_s_1_2_2(stage_PE_stage_PE_stage_PE_mux_3_nl,
      stage_PE_1_qr_1_10_1_lpi_2_dfm_8, or_tmp_979);
  assign BUTTERFLY_if_mux_15_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_8, stage_PE_1_qr_1_10_1_lpi_2_dfm_7,
      or_tmp_979);
  assign BUTTERFLY_if_mux_16_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_7, stage_PE_1_qr_1_10_1_lpi_2_dfm_6,
      or_tmp_979);
  assign BUTTERFLY_if_mux_17_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_6, stage_PE_1_qr_1_10_1_lpi_2_dfm_5,
      or_tmp_979);
  assign BUTTERFLY_if_mux_18_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_5, stage_PE_1_qr_1_10_1_lpi_2_dfm_4,
      or_tmp_979);
  assign BUTTERFLY_if_mux_19_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_4, stage_PE_1_qr_1_10_1_lpi_2_dfm_3,
      or_tmp_979);
  assign BUTTERFLY_if_mux_20_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_3, stage_PE_1_qr_1_10_1_lpi_2_dfm_2,
      or_tmp_979);
  assign BUTTERFLY_if_mux_21_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_2, stage_PE_1_qr_1_10_1_lpi_2_dfm_1,
      or_tmp_979);
  assign BUTTERFLY_if_mux_22_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_1, stage_PE_1_qr_1_10_1_lpi_2_dfm_0,
      or_tmp_979);
  assign BUTTERFLY_if_mux_23_nl = MUX_s_1_2_2(stage_PE_1_qr_1_10_1_lpi_2_dfm_0, stage_PE_1_qr_1_0_lpi_2_dfm,
      or_tmp_979);
  assign nl_z_out_7 = ({BUTTERFLY_if_mux_14_nl , BUTTERFLY_if_mux_15_nl , BUTTERFLY_if_mux_16_nl
      , BUTTERFLY_if_mux_17_nl , BUTTERFLY_if_mux_18_nl , BUTTERFLY_if_mux_19_nl
      , BUTTERFLY_if_mux_20_nl , BUTTERFLY_if_mux_21_nl , BUTTERFLY_if_mux_22_nl
      , BUTTERFLY_if_mux_23_nl}) + conv_u2u_9_10(BUTTERFLY_i_div_psp_sva_1);
  assign z_out_7 = nl_z_out_7[9:0];
  assign operator_6_false_mux1h_9_nl = MUX1HOT_s_1_10_2((drf_qr_lval_smx_lpi_3_dfm_mx0_10_5[5]),
      (drf_qr_lval_1_smx_lpi_3_dfm_mx1[10]), BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_1,
      drf_qr_lval_11_smx_lpi_3_dfm_10, reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd,
      (drf_qr_lval_13_smx_10_1_lpi_3_dfm[9]), (drf_qr_lval_14_smx_10_1_lpi_3_dfm[9]),
      (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[4]), (drf_qr_lval_16_smx_lpi_3_dfm_mx0_10_5[5]),
      (drf_qr_lval_11_smx_lpi_3_dfm_mx2[10]), {(fsm_output[5]) , (fsm_output[7])
      , operator_6_false_or_3_ssc , or_tmp_983 , operator_6_false_or_15_cse , operator_6_false_or_6_cse
      , or_dcpl_769 , operator_6_false_or_12_cse , (fsm_output[30]) , (fsm_output[32])});
  assign operator_6_false_mux1h_10_nl = MUX1HOT_s_1_10_2((drf_qr_lval_smx_lpi_3_dfm_mx0_10_5[4]),
      (drf_qr_lval_1_smx_lpi_3_dfm_mx1[9]), reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd,
      drf_qr_lval_11_smx_lpi_3_dfm_9, (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1[3]),
      (drf_qr_lval_13_smx_10_1_lpi_3_dfm[8]), (drf_qr_lval_14_smx_10_1_lpi_3_dfm[8]),
      (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[3]), (drf_qr_lval_16_smx_lpi_3_dfm_mx0_10_5[4]),
      (drf_qr_lval_11_smx_lpi_3_dfm_mx2[9]), {(fsm_output[5]) , (fsm_output[7]) ,
      operator_6_false_or_3_ssc , or_tmp_983 , operator_6_false_or_15_cse , operator_6_false_or_6_cse
      , or_dcpl_769 , operator_6_false_or_12_cse , (fsm_output[30]) , (fsm_output[32])});
  assign operator_6_false_mux1h_11_nl = MUX1HOT_v_3_10_2((drf_qr_lval_smx_lpi_3_dfm_mx0_10_5[3:1]),
      (drf_qr_lval_1_smx_lpi_3_dfm_mx1[8:6]), (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1[3:1]),
      (drf_qr_lval_11_smx_lpi_3_dfm_8_5[3:1]), (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1[2:0]),
      (drf_qr_lval_13_smx_10_1_lpi_3_dfm[7:5]), (drf_qr_lval_14_smx_10_1_lpi_3_dfm[7:5]),
      (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[2:0]), (drf_qr_lval_16_smx_lpi_3_dfm_mx0_10_5[3:1]),
      (drf_qr_lval_11_smx_lpi_3_dfm_mx2[8:6]), {(fsm_output[5]) , (fsm_output[7])
      , operator_6_false_or_3_ssc , or_tmp_983 , operator_6_false_or_15_cse , operator_6_false_or_6_cse
      , or_dcpl_769 , operator_6_false_or_12_cse , (fsm_output[30]) , (fsm_output[32])});
  assign operator_6_false_mux1h_12_nl = MUX1HOT_s_1_10_2((drf_qr_lval_smx_lpi_3_dfm_mx0_10_5[0]),
      (drf_qr_lval_1_smx_lpi_3_dfm_mx1[5]), (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1[0]),
      (drf_qr_lval_11_smx_lpi_3_dfm_8_5[0]), (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2[3]),
      (drf_qr_lval_13_smx_10_1_lpi_3_dfm[4]), (drf_qr_lval_14_smx_10_1_lpi_3_dfm[4]),
      (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[4]), (drf_qr_lval_16_smx_lpi_3_dfm_mx0_10_5[0]),
      (drf_qr_lval_11_smx_lpi_3_dfm_mx2[5]), {(fsm_output[5]) , (fsm_output[7]) ,
      operator_6_false_or_3_ssc , or_tmp_983 , operator_6_false_or_15_cse , operator_6_false_or_6_cse
      , or_dcpl_769 , operator_6_false_or_12_cse , (fsm_output[30]) , (fsm_output[32])});
  assign operator_6_false_mux1h_13_nl = MUX1HOT_v_3_10_2((drf_qr_lval_smx_lpi_3_dfm_mx0_4_0[4:2]),
      (drf_qr_lval_1_smx_lpi_3_dfm_mx1[4:2]), (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2[3:1]),
      (drf_qr_lval_11_smx_lpi_3_dfm_4_0[4:2]), (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2[2:0]),
      (drf_qr_lval_13_smx_10_1_lpi_3_dfm[3:1]), (drf_qr_lval_14_smx_10_1_lpi_3_dfm[3:1]),
      (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[3:1]), (drf_qr_lval_16_smx_lpi_3_dfm_mx0_4_0[4:2]),
      (drf_qr_lval_11_smx_lpi_3_dfm_mx2[4:2]), {(fsm_output[5]) , (fsm_output[7])
      , operator_6_false_or_3_ssc , or_tmp_983 , operator_6_false_or_15_cse , operator_6_false_or_6_cse
      , or_dcpl_769 , operator_6_false_or_12_cse , (fsm_output[30]) , (fsm_output[32])});
  assign operator_6_false_mux1h_14_nl = MUX1HOT_s_1_10_2((drf_qr_lval_smx_lpi_3_dfm_mx0_4_0[1]),
      (drf_qr_lval_1_smx_lpi_3_dfm_mx1[1]), (reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2[0]),
      (drf_qr_lval_11_smx_lpi_3_dfm_4_0[1]), reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3,
      (drf_qr_lval_13_smx_10_1_lpi_3_dfm[0]), (drf_qr_lval_14_smx_10_1_lpi_3_dfm[0]),
      (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[0]), (drf_qr_lval_16_smx_lpi_3_dfm_mx0_4_0[1]),
      (drf_qr_lval_11_smx_lpi_3_dfm_mx2[1]), {(fsm_output[5]) , (fsm_output[7]) ,
      operator_6_false_or_3_ssc , or_tmp_983 , operator_6_false_or_15_cse , operator_6_false_or_6_cse
      , or_dcpl_769 , operator_6_false_or_12_cse , (fsm_output[30]) , (fsm_output[32])});
  assign operator_6_false_or_23_nl = (fsm_output[19]) | (fsm_output[44]);
  assign operator_6_false_mux1h_15_nl = MUX1HOT_s_1_10_2((drf_qr_lval_smx_lpi_3_dfm_mx0_4_0[0]),
      (drf_qr_lval_1_smx_lpi_3_dfm_mx1[0]), reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3,
      (drf_qr_lval_11_smx_lpi_3_dfm_4_0[0]), BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm,
      drf_qr_lval_13_smx_0_lpi_3_dfm, drf_qr_lval_14_smx_0_lpi_3_dfm, drf_qr_lval_15_smx_0_lpi_3_dfm,
      (drf_qr_lval_16_smx_lpi_3_dfm_mx0_4_0[0]), (drf_qr_lval_11_smx_lpi_3_dfm_mx2[0]),
      {(fsm_output[5]) , (fsm_output[7]) , operator_6_false_or_3_ssc , or_tmp_983
      , operator_6_false_or_23_nl , or_tmp_234 , or_dcpl_661 , or_dcpl_397 , (fsm_output[30])
      , (fsm_output[32])});
  assign nl_operator_6_false_acc_1_nl = ({1'b1 , (~ (rtn_out[5:1]))}) + 6'b000001;
  assign operator_6_false_acc_1_nl = nl_operator_6_false_acc_1_nl[5:0];
  assign nl_operator_6_false_2_acc_1_nl = ({1'b1 , (~ (rtn_out[5:1]))}) + 6'b000001;
  assign operator_6_false_2_acc_1_nl = nl_operator_6_false_2_acc_1_nl[5:0];
  assign nl_operator_6_false_4_acc_3_nl = ({1'b1 , (~ (return_add_generic_AC_RND_CONV_false_11_ls_sva[5:1]))})
      + 6'b000001;
  assign operator_6_false_4_acc_3_nl = nl_operator_6_false_4_acc_3_nl[5:0];
  assign nl_operator_6_false_23_acc_3_nl = ({1'b1 , (~ (return_add_generic_AC_RND_CONV_false_10_ls_sva[5:1]))})
      + 6'b000001;
  assign operator_6_false_23_acc_3_nl = nl_operator_6_false_23_acc_3_nl[5:0];
  assign nl_operator_6_false_17_acc_3_nl = ({1'b1 , (~ (rtn_out[5:1]))}) + 6'b000001;
  assign operator_6_false_17_acc_3_nl = nl_operator_6_false_17_acc_3_nl[5:0];
  assign nl_operator_6_false_21_acc_3_nl = ({1'b1 , (~ (return_add_generic_AC_RND_CONV_false_12_ls_sva[5:1]))})
      + 6'b000001;
  assign operator_6_false_21_acc_3_nl = nl_operator_6_false_21_acc_3_nl[5:0];
  assign nl_operator_6_false_29_acc_1_nl = ({1'b1 , (~ (rtn_out[5:1]))}) + 6'b000001;
  assign operator_6_false_29_acc_1_nl = nl_operator_6_false_29_acc_1_nl[5:0];
  assign nl_operator_6_false_31_acc_1_nl = ({1'b1 , (~ (rtn_out[5:1]))}) + 6'b000001;
  assign operator_6_false_31_acc_1_nl = nl_operator_6_false_31_acc_1_nl[5:0];
  assign operator_6_false_mux1h_16_nl = MUX1HOT_v_6_8_2(operator_6_false_acc_1_nl,
      operator_6_false_2_acc_1_nl, operator_6_false_4_acc_3_nl, operator_6_false_23_acc_3_nl,
      operator_6_false_17_acc_3_nl, operator_6_false_21_acc_3_nl, operator_6_false_29_acc_1_nl,
      operator_6_false_31_acc_1_nl, {(fsm_output[5]) , (fsm_output[7]) , operator_6_false_or_ssc
      , operator_6_false_or_1_ssc , return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
      , operator_6_false_or_20_cse , (fsm_output[30]) , (fsm_output[32])});
  assign operator_6_false_or_24_nl = (fsm_output[5]) | (fsm_output[7]) | return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
      | (fsm_output[30]) | (fsm_output[32]);
  assign operator_6_false_mux1h_17_nl = MUX1HOT_s_1_4_2((~ (rtn_out[0])), (~ (return_add_generic_AC_RND_CONV_false_11_ls_sva[0])),
      (~ (return_add_generic_AC_RND_CONV_false_10_ls_sva[0])), (~ (return_add_generic_AC_RND_CONV_false_12_ls_sva[0])),
      {operator_6_false_or_24_nl , operator_6_false_or_ssc , operator_6_false_or_1_ssc
      , operator_6_false_or_20_cse});
  assign nl_z_out_8 = conv_u2u_11_13({operator_6_false_mux1h_9_nl , operator_6_false_mux1h_10_nl
      , operator_6_false_mux1h_11_nl , operator_6_false_mux1h_12_nl , operator_6_false_mux1h_13_nl
      , operator_6_false_mux1h_14_nl , operator_6_false_mux1h_15_nl}) + conv_s2u_7_13({operator_6_false_mux1h_16_nl
      , operator_6_false_mux1h_17_nl});
  assign z_out_8 = nl_z_out_8[12:0];
  assign BUTTERFLY_1_mux_1_nl = MUX_s_1_2_2((~ (in_u_rsci_q_d[9])), (BUTTERFLY_1_fry_9_0_sva[9]),
      fsm_output[55]);
  assign BUTTERFLY_1_and_2_nl = BUTTERFLY_1_mux_1_nl & (~ return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse)
      & BUTTERFLY_1_nor_1_seb;
  assign BUTTERFLY_1_mux1h_5_nl = MUX1HOT_v_5_3_2((BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[8:4]),
      (~ (in_u_rsci_q_d[8:4])), (BUTTERFLY_1_fry_9_0_sva[8:4]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , (fsm_output[54]) , (fsm_output[55])});
  assign BUTTERFLY_1_and_3_nl = MUX_v_5_2_2(5'b00000, BUTTERFLY_1_mux1h_5_nl, BUTTERFLY_1_nor_1_seb);
  assign BUTTERFLY_1_mux1h_6_nl = MUX1HOT_v_4_4_2((BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[3:0]),
      (~ (z_out_21[3:0])), (~ (in_u_rsci_q_d[3:0])), (BUTTERFLY_1_fry_9_0_sva[3:0]),
      {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , (fsm_output[54]) , (fsm_output[55])});
  assign BUTTERFLY_1_nor_2_nl = ~(return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      | (fsm_output[55:54]!=2'b00));
  assign BUTTERFLY_1_BUTTERFLY_1_and_2_nl = MUX_v_2_2_2(2'b00, (z_out_21[1:0]), BUTTERFLY_1_nor_2_nl);
  assign nl_z_out_19 = conv_u2u_10_11({BUTTERFLY_1_and_2_nl , BUTTERFLY_1_and_3_nl
      , BUTTERFLY_1_mux1h_6_nl}) + conv_u2u_4_11({BUTTERFLY_1_BUTTERFLY_1_and_2_nl
      , 2'b01});
  assign z_out_19 = nl_z_out_19[10:0];
  assign nl_z_out_20 = (z_out_28[10:1]) + 10'b0000000001;
  assign z_out_20 = nl_z_out_20[9:0];
  assign BUTTERFLY_i_mux1h_24_nl = MUX1HOT_s_1_5_2(return_extract_12_return_extract_12_or_1_cse_sva_1,
      return_extract_13_return_extract_13_or_1_cse_sva_1, BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm,
      return_extract_44_return_extract_44_or_1_cse_sva_1, return_extract_45_return_extract_45_or_1_cse_sva_1,
      {(fsm_output[10]) , (fsm_output[12]) , BUTTERFLY_i_or_4_cse , (fsm_output[35])
      , (fsm_output[37])});
  assign BUTTERFLY_i_and_14_nl = BUTTERFLY_i_mux1h_24_nl & BUTTERFLY_i_nor_2_cse_1;
  assign BUTTERFLY_i_mux1h_25_nl = MUX1HOT_s_1_5_2(return_extract_15_return_extract_15_nor_cse_sva_mx1,
      return_add_generic_AC_RND_CONV_false_3_r_nan_mux1h_cse, (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[51]),
      return_extract_15_return_extract_15_nor_cse_sva_mx2, return_add_generic_AC_RND_CONV_false_16_r_nan_mux1h_cse,
      {(fsm_output[10]) , (fsm_output[12]) , BUTTERFLY_i_or_4_cse , (fsm_output[35])
      , (fsm_output[37])});
  assign BUTTERFLY_i_and_15_nl = BUTTERFLY_i_mux1h_25_nl & BUTTERFLY_i_nor_2_cse_1;
  assign BUTTERFLY_i_mux1h_26_nl = MUX1HOT_v_37_5_2((stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0[50:14]),
      (stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0[50:14]), (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[50:14]),
      (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1[50:14]), (stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0[50:14]),
      {(fsm_output[10]) , (fsm_output[12]) , BUTTERFLY_i_or_4_cse , (fsm_output[35])
      , (fsm_output[37])});
  assign BUTTERFLY_i_and_16_nl = MUX_v_37_2_2(37'b0000000000000000000000000000000000000,
      BUTTERFLY_i_mux1h_26_nl, BUTTERFLY_i_nor_2_cse_1);
  assign BUTTERFLY_i_mux1h_27_nl = MUX1HOT_v_3_6_2(BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_0,
      (stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0[13:11]), (stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0[13:11]),
      (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[13:11]), (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1[13:11]),
      (stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0[13:11]), {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , (fsm_output[10]) , (fsm_output[12]) , BUTTERFLY_i_or_4_cse , (fsm_output[35])
      , (fsm_output[37])});
  assign not_815_nl = ~ return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  assign BUTTERFLY_i_and_17_nl = MUX_v_3_2_2(3'b000, BUTTERFLY_i_mux1h_27_nl, not_815_nl);
  assign BUTTERFLY_i_mux1h_28_nl = MUX1HOT_s_1_6_2(BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1,
      (stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0[10]), (stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0[10]),
      (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[10]), (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1[10]),
      (stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0[10]), {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , (fsm_output[10]) , (fsm_output[12]) , BUTTERFLY_i_or_4_cse , (fsm_output[35])
      , (fsm_output[37])});
  assign BUTTERFLY_i_and_18_nl = BUTTERFLY_i_mux1h_28_nl & (~ return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse);
  assign BUTTERFLY_i_mux1h_29_nl = MUX1HOT_v_5_7_2(({1'b0, BUTTERFLY_i_div_psp_sva_1[8:5]}),
      reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd, (stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0[9:5]),
      (stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0[9:5]), (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[9:5]),
      (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1[9:5]), (stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0[9:5]),
      {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , (fsm_output[10]) , (fsm_output[12]) , BUTTERFLY_i_or_4_cse , (fsm_output[35])
      , (fsm_output[37])});
  assign BUTTERFLY_i_mux1h_30_nl = MUX1HOT_v_5_7_2((BUTTERFLY_i_div_psp_sva_1[4:0]),
      reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1, (stage_PE_tmp_re_d_1_lpi_3_dfm_50_0_mx0[4:0]),
      (stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0[4:0]), (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[4:0]),
      (stage_PE_1_tmp_re_d_1_lpi_3_dfm_50_0_mx1[4:0]), (stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0[4:0]),
      {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , (fsm_output[10]) , (fsm_output[12]) , BUTTERFLY_i_or_4_cse , (fsm_output[35])
      , (fsm_output[37])});
  assign BUTTERFLY_i_BUTTERFLY_i_and_1_nl = (BUTTERFLY_else_1_BUTTERFLY_else_1_and_cse[1])
      & (~(return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse | (fsm_output[10])
      | (fsm_output[12]) | (fsm_output[14]) | (fsm_output[35]) | (fsm_output[37])
      | (fsm_output[39])));
  assign BUTTERFLY_i_mux1h_31_nl = MUX1HOT_s_1_5_2((BUTTERFLY_else_1_BUTTERFLY_else_1_and_cse[1]),
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_12_op_smaller_qr_0_lpi_3_dfm,
      return_extract_19_return_extract_19_or_sva_1, return_extract_51_return_extract_51_or_sva_1,
      {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , or_dcpl_548 , or_dcpl_404
      , (fsm_output[14]) , (fsm_output[39])});
  assign BUTTERFLY_i_and_19_nl = BUTTERFLY_i_mux1h_31_nl & (~ return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse);
  assign BUTTERFLY_i_mux1h_32_nl = MUX1HOT_s_1_5_2((BUTTERFLY_else_1_BUTTERFLY_else_1_and_cse[1]),
      drf_qr_lval_14_smx_0_lpi_3_dfm, drf_qr_lval_15_smx_0_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_6_m_r_51_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_19_m_r_51_lpi_3_dfm_mx0, {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , or_dcpl_548 , or_dcpl_404 , (fsm_output[14]) , (fsm_output[39])});
  assign BUTTERFLY_i_and_20_nl = BUTTERFLY_i_mux1h_32_nl & (~ return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse);
  assign BUTTERFLY_i_mux1h_33_nl = MUX1HOT_s_1_5_2((BUTTERFLY_else_1_BUTTERFLY_else_1_and_cse[1]),
      return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_0, (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[50]),
      (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[50]), (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[50]),
      {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , or_dcpl_548 , or_dcpl_404
      , (fsm_output[14]) , (fsm_output[39])});
  assign BUTTERFLY_i_and_21_nl = BUTTERFLY_i_mux1h_33_nl & (~ return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse);
  assign BUTTERFLY_i_mux1h_34_nl = MUX1HOT_v_33_5_2((signext_33_1(BUTTERFLY_else_1_BUTTERFLY_else_1_and_cse[1])),
      (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[49:17]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[49:17]), (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[49:17]),
      (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[49:17]), {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , or_dcpl_548 , or_dcpl_404 , (fsm_output[14]) , (fsm_output[39])});
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_not_10_nl = ~ return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  assign BUTTERFLY_i_and_22_nl = MUX_v_33_2_2(33'b000000000000000000000000000000000,
      BUTTERFLY_i_mux1h_34_nl, return_add_generic_AC_RND_CONV_false_11_op_bigger_not_10_nl);
  assign BUTTERFLY_i_mux1h_35_nl = MUX1HOT_s_1_5_2((BUTTERFLY_else_1_BUTTERFLY_else_1_and_cse[0]),
      (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[16]), (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[16]),
      (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[16]), (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[16]),
      {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , or_dcpl_548 , or_dcpl_404
      , (fsm_output[14]) , (fsm_output[39])});
  assign BUTTERFLY_i_and_23_nl = BUTTERFLY_i_mux1h_35_nl & (~ return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse);
  assign BUTTERFLY_i_and_25_nl = (~ inverse_lpi_1_dfm_1) & return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse;
  assign BUTTERFLY_i_and_26_nl = inverse_lpi_1_dfm_1 & return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse;
  assign BUTTERFLY_i_mux1h_36_nl = MUX1HOT_v_5_6_2(BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0,
      (z_out_3[15:11]), (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[15:11]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[15:11]), (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[15:11]),
      (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[15:11]), {BUTTERFLY_i_and_25_nl
      , BUTTERFLY_i_and_26_nl , or_dcpl_548 , or_dcpl_404 , (fsm_output[14]) , (fsm_output[39])});
  assign return_add_generic_AC_RND_CONV_false_11_op_bigger_not_12_nl = ~ return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse;
  assign BUTTERFLY_i_and_24_nl = MUX_v_5_2_2(5'b00000, BUTTERFLY_i_mux1h_36_nl, return_add_generic_AC_RND_CONV_false_11_op_bigger_not_12_nl);
  assign BUTTERFLY_i_mux1h_37_nl = MUX1HOT_s_1_5_2((BUTTERFLY_i_conc_3_itm_10_9[1]),
      (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[10]), (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[10]),
      (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[10]), (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[10]),
      {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , or_dcpl_548 , or_dcpl_404
      , (fsm_output[14]) , (fsm_output[39])});
  assign BUTTERFLY_i_and_27_nl = BUTTERFLY_i_mux1h_37_nl & (~ return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse);
  assign BUTTERFLY_i_mux1h_38_nl = MUX1HOT_s_1_6_2(stage_PE_1_index_const_9_1_lpi_2_dfm_8,
      (BUTTERFLY_i_conc_3_itm_10_9[0]), (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[9]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[9]), (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[9]),
      (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[9]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , or_dcpl_548 ,
      or_dcpl_404 , (fsm_output[14]) , (fsm_output[39])});
  assign BUTTERFLY_i_mux1h_39_nl = MUX1HOT_s_1_6_2(stage_PE_1_index_const_9_1_lpi_2_dfm_7,
      (BUTTERFLY_i_conc_3_itm_8_0[8]), (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[8]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[8]), (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[8]),
      (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[8]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , or_dcpl_548 ,
      or_dcpl_404 , (fsm_output[14]) , (fsm_output[39])});
  assign BUTTERFLY_i_mux1h_40_nl = MUX1HOT_s_1_6_2(stage_PE_1_index_const_9_1_lpi_2_dfm_6,
      (BUTTERFLY_i_conc_3_itm_8_0[7]), (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[7]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[7]), (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[7]),
      (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[7]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , or_dcpl_548 ,
      or_dcpl_404 , (fsm_output[14]) , (fsm_output[39])});
  assign BUTTERFLY_i_mux1h_41_nl = MUX1HOT_s_1_6_2(stage_PE_1_index_const_9_1_lpi_2_dfm_5,
      (BUTTERFLY_i_conc_3_itm_8_0[6]), (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[6]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[6]), (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[6]),
      (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[6]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , or_dcpl_548 ,
      or_dcpl_404 , (fsm_output[14]) , (fsm_output[39])});
  assign BUTTERFLY_i_mux1h_42_nl = MUX1HOT_s_1_6_2(stage_PE_1_index_const_9_1_lpi_2_dfm_4,
      (BUTTERFLY_i_conc_3_itm_8_0[5]), (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[5]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[5]), (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[5]),
      (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[5]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , or_dcpl_548 ,
      or_dcpl_404 , (fsm_output[14]) , (fsm_output[39])});
  assign BUTTERFLY_i_mux1h_43_nl = MUX1HOT_s_1_6_2(stage_PE_1_index_const_9_1_lpi_2_dfm_3,
      (BUTTERFLY_i_conc_3_itm_8_0[4]), (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[4]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[4]), (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[4]),
      (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[4]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , or_dcpl_548 ,
      or_dcpl_404 , (fsm_output[14]) , (fsm_output[39])});
  assign BUTTERFLY_i_mux1h_44_nl = MUX1HOT_s_1_6_2(stage_PE_1_index_const_9_1_lpi_2_dfm_2,
      (BUTTERFLY_i_conc_3_itm_8_0[3]), (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[3]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[3]), (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[3]),
      (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[3]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , or_dcpl_548 ,
      or_dcpl_404 , (fsm_output[14]) , (fsm_output[39])});
  assign BUTTERFLY_i_mux1h_45_nl = MUX1HOT_s_1_6_2(stage_PE_1_index_const_9_1_lpi_2_dfm_1,
      (BUTTERFLY_i_conc_3_itm_8_0[2]), (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[2]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[2]), (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[2]),
      (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[2]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , or_dcpl_548 ,
      or_dcpl_404 , (fsm_output[14]) , (fsm_output[39])});
  assign BUTTERFLY_i_mux1h_46_nl = MUX1HOT_s_1_6_2(stage_PE_1_index_const_9_1_lpi_2_dfm_0,
      (BUTTERFLY_i_conc_3_itm_8_0[1]), (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[1]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[1]), (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[1]),
      (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[1]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , or_dcpl_548 ,
      or_dcpl_404 , (fsm_output[14]) , (fsm_output[39])});
  assign BUTTERFLY_i_mux1h_47_nl = MUX1HOT_s_1_6_2(stage_PE_1_index_const_0_lpi_2_dfm,
      (BUTTERFLY_i_conc_3_itm_8_0[0]), (return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1[0]),
      (return_add_generic_AC_RND_CONV_false_18_m_r_50_0_lpi_3_dfm[0]), (return_add_generic_AC_RND_CONV_false_6_m_r_50_0_lpi_3_dfm_1[0]),
      (return_add_generic_AC_RND_CONV_false_19_m_r_50_0_lpi_3_dfm_1[0]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , or_dcpl_548 ,
      or_dcpl_404 , (fsm_output[14]) , (fsm_output[39])});
  assign nl_z_out_21 = $signed(conv_u2s_53_54({BUTTERFLY_i_and_14_nl , BUTTERFLY_i_and_15_nl
      , BUTTERFLY_i_and_16_nl , BUTTERFLY_i_and_17_nl , BUTTERFLY_i_and_18_nl , BUTTERFLY_i_mux1h_29_nl
      , BUTTERFLY_i_mux1h_30_nl})) * $signed(({BUTTERFLY_i_BUTTERFLY_i_and_1_nl ,
      BUTTERFLY_i_and_19_nl , BUTTERFLY_i_and_20_nl , BUTTERFLY_i_and_21_nl , BUTTERFLY_i_and_22_nl
      , BUTTERFLY_i_and_23_nl , BUTTERFLY_i_and_24_nl , BUTTERFLY_i_and_27_nl , BUTTERFLY_i_mux1h_38_nl
      , BUTTERFLY_i_mux1h_39_nl , BUTTERFLY_i_mux1h_40_nl , BUTTERFLY_i_mux1h_41_nl
      , BUTTERFLY_i_mux1h_42_nl , BUTTERFLY_i_mux1h_43_nl , BUTTERFLY_i_mux1h_44_nl
      , BUTTERFLY_i_mux1h_45_nl , BUTTERFLY_i_mux1h_46_nl , BUTTERFLY_i_mux1h_47_nl}));
  assign z_out_21 = nl_z_out_21[105:0];
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_10_nl = MUX1HOT_s_1_6_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_0[5]),
      (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
      (stage_PE_1_x_re_d_sva[62]), (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1[9]),
      (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
      (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[9]), {return_add_generic_AC_RND_CONV_false_e_dif_qif_or_cse
      , (fsm_output[14]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse
      , return_add_generic_AC_RND_CONV_false_e_dif_qif_and_1_cse , (fsm_output[39])
      , (fsm_output[43])});
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_and_7_nl = return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_10_nl
      & (~ (fsm_output[54]));
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_11_nl = MUX1HOT_v_5_7_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_0[4:0]),
      (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[9:5]),
      (stage_PE_1_x_re_d_sva[61:57]), (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1[8:4]),
      (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[9:5]),
      (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[8:4]), (~
      (z_out_19[9:5])), {return_add_generic_AC_RND_CONV_false_e_dif_qif_or_cse ,
      (fsm_output[14]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse
      , return_add_generic_AC_RND_CONV_false_e_dif_qif_and_1_cse , (fsm_output[39])
      , (fsm_output[43]) , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_12_nl = MUX1HOT_v_4_7_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_1[56:53]),
      (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[4:1]),
      (stage_PE_1_x_re_d_sva[56:53]), (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0w0_10_1[3:0]),
      (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[4:1]),
      (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[3:0]), (~
      (z_out_19[4:1])), {return_add_generic_AC_RND_CONV_false_e_dif_qif_or_cse ,
      (fsm_output[14]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse
      , return_add_generic_AC_RND_CONV_false_e_dif_qif_and_1_cse , (fsm_output[39])
      , (fsm_output[43]) , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_13_nl = MUX1HOT_s_1_7_2((stage_PE_1_tmp_im_d_1_sva_1_rsp_1[52]),
      (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[0]),
      (stage_PE_1_x_re_d_sva[52]), stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0, (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[0]),
      return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1, (~ (z_out_19[0])),
      {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , (fsm_output[14])
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse , (fsm_output[37])
      , (fsm_output[39]) , (fsm_output[43]) , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_14_nl = MUX1HOT_s_1_7_2((out_f_d_rsci_q_d[62]),
      BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1, (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1[9]),
      (in_f_d_rsci_q_d[62]), BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_1, (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1[9]),
      (stage_PE_1_x_im_d_sva[62]), {(fsm_output[5]) , BUTTERFLY_i_or_4_cse , (fsm_output[16])
      , (fsm_output[30]) , (fsm_output[37]) , (fsm_output[41]) , (fsm_output[43])});
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_nor_1_nl = ~(return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_14_nl
      | (fsm_output[54]));
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_15_nl = MUX1HOT_s_1_7_2((out_f_d_rsci_q_d[61]),
      (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[4]), (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1[8]),
      (in_f_d_rsci_q_d[61]), reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd, (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1[8]),
      (stage_PE_1_x_im_d_sva[61]), {(fsm_output[5]) , BUTTERFLY_i_or_4_cse , (fsm_output[16])
      , (fsm_output[30]) , (fsm_output[37]) , (fsm_output[41]) , (fsm_output[43])});
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_return_add_generic_AC_RND_CONV_false_e_dif_qif_nor_2_nl
      = ~(return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_15_nl | (fsm_output[54]));
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_16_nl = MUX1HOT_v_4_7_2((out_f_d_rsci_q_d[60:57]),
      (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[3:0]), (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1[7:4]),
      (in_f_d_rsci_q_d[60:57]), reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1, (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1[7:4]),
      (stage_PE_1_x_im_d_sva[60:57]), {(fsm_output[5]) , BUTTERFLY_i_or_4_cse , (fsm_output[16])
      , (fsm_output[30]) , (fsm_output[37]) , (fsm_output[41]) , (fsm_output[43])});
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_return_add_generic_AC_RND_CONV_false_e_dif_qif_nor_3_nl
      = ~(MUX_v_4_2_2(return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_16_nl,
      4'b1111, (fsm_output[54])));
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_17_nl = MUX1HOT_v_4_8_2((~
      (out_f_d_rsci_q_d[56:53])), (~ (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[4:1])),
      (~ (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1[3:0])),
      (~ (in_f_d_rsci_q_d[56:53])), (~ reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2),
      (~ (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1[3:0])),
      (~ (stage_PE_1_x_im_d_sva[56:53])), ({1'b0, in_u_rsci_q_d[15:13]}), {(fsm_output[5])
      , BUTTERFLY_i_or_4_cse , (fsm_output[16]) , (fsm_output[30]) , (fsm_output[37])
      , (fsm_output[41]) , (fsm_output[43]) , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_18_nl = MUX1HOT_s_1_8_2((~
      (out_f_d_rsci_q_d[52])), (~ (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1[0])),
      (~ return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1), (~ (in_f_d_rsci_q_d[52])),
      (~ reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3), (~ return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1),
      (~ (stage_PE_1_x_im_d_sva[52])), (in_u_rsci_q_d[12]), {(fsm_output[5]) , BUTTERFLY_i_or_4_cse
      , (fsm_output[16]) , (fsm_output[30]) , (fsm_output[37]) , (fsm_output[41])
      , (fsm_output[43]) , (fsm_output[54])});
  assign nl_acc_12_nl = ({(~ (fsm_output[54])) , return_add_generic_AC_RND_CONV_false_e_dif_qif_and_7_nl
      , return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_11_nl , return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_12_nl
      , return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_13_nl , (~ (fsm_output[54]))})
      + conv_u2u_12_13({return_add_generic_AC_RND_CONV_false_e_dif_qif_nor_1_nl ,
      return_add_generic_AC_RND_CONV_false_e_dif_qif_return_add_generic_AC_RND_CONV_false_e_dif_qif_nor_2_nl
      , return_add_generic_AC_RND_CONV_false_e_dif_qif_return_add_generic_AC_RND_CONV_false_e_dif_qif_nor_3_nl
      , return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_17_nl , return_add_generic_AC_RND_CONV_false_e_dif_qif_mux1h_18_nl
      , 1'b1});
  assign acc_12_nl = nl_acc_12_nl[12:0];
  assign z_out_23 = readslicef_13_12_1(acc_12_nl);
  assign return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_10_nl = MUX1HOT_s_1_6_2((out_f_d_rsci_q_d[62]),
      BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_1, (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
      (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1[9]), (in_f_d_rsci_q_d[62]),
      (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
      {or_219_cse , or_dcpl_404 , (fsm_output[14]) , (fsm_output[18]) , or_200_cse
      , (fsm_output[39])});
  assign return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_11_nl = MUX1HOT_s_1_6_2((out_f_d_rsci_q_d[61]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd, (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[9]),
      (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1[8]), (in_f_d_rsci_q_d[61]),
      (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[9]),
      {or_219_cse , or_dcpl_404 , (fsm_output[14]) , (fsm_output[18]) , or_200_cse
      , (fsm_output[39])});
  assign return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_12_nl = MUX1HOT_v_4_6_2((out_f_d_rsci_q_d[60:57]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1, (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[8:5]),
      (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1[7:4]), (in_f_d_rsci_q_d[60:57]),
      (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[8:5]),
      {or_219_cse , or_dcpl_404 , (fsm_output[14]) , (fsm_output[18]) , or_200_cse
      , (fsm_output[39])});
  assign return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_13_nl = MUX1HOT_v_4_6_2((out_f_d_rsci_q_d[56:53]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2, (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[4:1]),
      (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1[3:0]), (in_f_d_rsci_q_d[56:53]),
      (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[4:1]),
      {or_219_cse , or_dcpl_404 , (fsm_output[14]) , (fsm_output[18]) , or_200_cse
      , (fsm_output[39])});
  assign return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_14_nl = MUX1HOT_s_1_6_2((out_f_d_rsci_q_d[52]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3, (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[0]),
      return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1, (in_f_d_rsci_q_d[52]),
      (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[0]),
      {or_219_cse , or_dcpl_404 , (fsm_output[14]) , (fsm_output[18]) , or_200_cse
      , (fsm_output[39])});
  assign return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_15_nl = MUX1HOT_v_2_5_2((~
      (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[5:4])), (~ (stage_PE_1_x_im_d_sva[62:61])),
      (~ (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5[5:4])), (~ BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1),
      (~ (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5[5:4])), {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_add_generic_AC_RND_CONV_false_e_dif1_or_1_ssc , (fsm_output[12]) ,
      BUTTERFLY_i_or_4_cse , (fsm_output[37])});
  assign return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_16_nl = MUX1HOT_v_4_5_2((~
      (stage_PE_1_tmp_im_d_1_sva_1_rsp_0[3:0])), (~ (stage_PE_1_x_im_d_sva[60:57])),
      (~ (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5[3:0])), (~ (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[8:5])),
      (~ (stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5[3:0])), {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_add_generic_AC_RND_CONV_false_e_dif1_or_1_ssc , (fsm_output[12]) ,
      BUTTERFLY_i_or_4_cse , (fsm_output[37])});
  assign return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_17_nl = MUX1HOT_v_4_5_2((~
      (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[56:53])), (~ (stage_PE_1_x_im_d_sva[56:53])),
      (~ stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1), (~ (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[4:1])),
      (~ stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1), {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_add_generic_AC_RND_CONV_false_e_dif1_or_1_ssc , (fsm_output[12]) ,
      BUTTERFLY_i_or_4_cse , (fsm_output[37])});
  assign return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_18_nl = MUX1HOT_s_1_5_2((~
      (stage_PE_1_tmp_im_d_1_sva_1_rsp_1[52])), (~ (stage_PE_1_x_im_d_sva[52])),
      (~ stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0), (~ (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[0])),
      (~ stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0), {return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_add_generic_AC_RND_CONV_false_e_dif1_or_1_ssc , (fsm_output[12]) ,
      BUTTERFLY_i_or_4_cse , (fsm_output[37])});
  assign nl_acc_13_nl = ({1'b1 , return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_10_nl
      , return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_11_nl , return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_12_nl
      , return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_13_nl , return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_14_nl
      , 1'b1}) + conv_u2u_12_13({return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_15_nl
      , return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_16_nl , return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_17_nl
      , return_add_generic_AC_RND_CONV_false_e_dif1_mux1h_18_nl , 1'b1});
  assign acc_13_nl = nl_acc_13_nl[12:0];
  assign z_out_24 = readslicef_13_12_1(acc_13_nl);
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_10_nl = MUX1HOT_v_2_6_2((stage_PE_1_x_im_d_sva[62:61]),
      (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5[5:4]), BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1,
      (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1[9:8]), (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1[9:8]),
      (z_out_23[10:9]), {return_add_generic_AC_RND_CONV_false_1_e_dif1_or_6_cse ,
      (fsm_output[12]) , BUTTERFLY_i_or_4_cse , (fsm_output[16]) , (fsm_output[41])
      , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_11_nl = MUX1HOT_v_4_6_2((stage_PE_1_x_im_d_sva[60:57]),
      (stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5[3:0]), (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[8:5]),
      (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1[7:4]), (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1[7:4]),
      (z_out_23[8:5]), {return_add_generic_AC_RND_CONV_false_1_e_dif1_or_6_cse ,
      (fsm_output[12]) , BUTTERFLY_i_or_4_cse , (fsm_output[16]) , (fsm_output[41])
      , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_12_nl = MUX1HOT_v_4_6_2((stage_PE_1_x_im_d_sva[56:53]),
      stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1, (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[4:1]),
      (return_add_generic_AC_RND_CONV_false_7_e_r_qr_10_1_lpi_3_dfm_1[3:0]), (return_add_generic_AC_RND_CONV_false_20_e_r_qr_10_1_lpi_3_dfm_1[3:0]),
      (z_out_23[4:1]), {return_add_generic_AC_RND_CONV_false_1_e_dif1_or_6_cse ,
      (fsm_output[12]) , BUTTERFLY_i_or_4_cse , (fsm_output[16]) , (fsm_output[41])
      , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_13_nl = MUX1HOT_s_1_6_2((stage_PE_1_x_im_d_sva[52]),
      stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0, (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[0]),
      return_add_generic_AC_RND_CONV_false_7_e_r_qr_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_20_e_r_qr_0_lpi_3_dfm_1,
      (z_out_23[0]), {return_add_generic_AC_RND_CONV_false_1_e_dif1_or_6_cse , (fsm_output[12])
      , BUTTERFLY_i_or_4_cse , (fsm_output[16]) , (fsm_output[41]) , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_14_nl = MUX1HOT_s_1_8_2((out_f_d_rsci_q_d[62]),
      BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_1, (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
      (stage_PE_1_x_re_d_sva[62]), (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1[9]),
      (in_f_d_rsci_q_d[62]), (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[10]),
      (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[9]), {(fsm_output[7])
      , (fsm_output[12]) , (fsm_output[14]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse
      , (fsm_output[18]) , (fsm_output[32]) , (fsm_output[39]) , (fsm_output[43])});
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_return_add_generic_AC_RND_CONV_false_1_e_dif1_nand_2_nl
      = ~(return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_14_nl & (~ (fsm_output[54])));
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_15_nl = MUX1HOT_s_1_8_2((out_f_d_rsci_q_d[61]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd, (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[9]),
      (stage_PE_1_x_re_d_sva[61]), (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1[8]),
      (in_f_d_rsci_q_d[61]), (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[9]),
      (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[8]), {(fsm_output[7])
      , (fsm_output[12]) , (fsm_output[14]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse
      , (fsm_output[18]) , (fsm_output[32]) , (fsm_output[39]) , (fsm_output[43])});
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_nor_3_nl = ~(return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_15_nl
      | (fsm_output[54]));
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_16_nl = MUX1HOT_v_4_8_2((out_f_d_rsci_q_d[60:57]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1, (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[8:5]),
      (stage_PE_1_x_re_d_sva[60:57]), (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1[7:4]),
      (in_f_d_rsci_q_d[60:57]), (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[8:5]),
      (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[7:4]), {(fsm_output[7])
      , (fsm_output[12]) , (fsm_output[14]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse
      , (fsm_output[18]) , (fsm_output[32]) , (fsm_output[39]) , (fsm_output[43])});
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_nor_4_nl = ~(MUX_v_4_2_2(return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_16_nl,
      4'b1111, (fsm_output[54])));
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_17_nl = MUX1HOT_v_4_8_2((out_f_d_rsci_q_d[56:53]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2, (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[4:1]),
      (stage_PE_1_x_re_d_sva[56:53]), (return_add_generic_AC_RND_CONV_false_8_e_r_qr_10_1_lpi_3_dfm_1[3:0]),
      (in_f_d_rsci_q_d[56:53]), (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[4:1]),
      (return_add_generic_AC_RND_CONV_false_21_e_r_qr_10_1_lpi_3_dfm_1[3:0]), {(fsm_output[7])
      , (fsm_output[12]) , (fsm_output[14]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse
      , (fsm_output[18]) , (fsm_output[32]) , (fsm_output[39]) , (fsm_output[43])});
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_nor_5_nl = ~(MUX_v_4_2_2(return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_17_nl,
      4'b1111, (fsm_output[54])));
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_18_nl = MUX1HOT_s_1_8_2((out_f_d_rsci_q_d[52]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3, (return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1[0]),
      (stage_PE_1_x_re_d_sva[52]), return_add_generic_AC_RND_CONV_false_8_e_r_qr_0_lpi_3_dfm_1,
      (in_f_d_rsci_q_d[52]), (return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1[0]),
      return_add_generic_AC_RND_CONV_false_21_e_r_qr_0_lpi_3_dfm_1, {(fsm_output[7])
      , (fsm_output[12]) , (fsm_output[14]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse
      , (fsm_output[18]) , (fsm_output[32]) , (fsm_output[39]) , (fsm_output[43])});
  assign return_add_generic_AC_RND_CONV_false_1_e_dif1_return_add_generic_AC_RND_CONV_false_1_e_dif1_nand_3_nl
      = ~(return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_18_nl & (~ (fsm_output[54])));
  assign nl_acc_14_nl = ({(~ (fsm_output[54])) , return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_10_nl
      , return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_11_nl , return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_12_nl
      , return_add_generic_AC_RND_CONV_false_1_e_dif1_mux1h_13_nl , (~ (fsm_output[54]))})
      + conv_u2u_12_13({return_add_generic_AC_RND_CONV_false_1_e_dif1_return_add_generic_AC_RND_CONV_false_1_e_dif1_nand_2_nl
      , return_add_generic_AC_RND_CONV_false_1_e_dif1_nor_3_nl , return_add_generic_AC_RND_CONV_false_1_e_dif1_nor_4_nl
      , return_add_generic_AC_RND_CONV_false_1_e_dif1_nor_5_nl , return_add_generic_AC_RND_CONV_false_1_e_dif1_return_add_generic_AC_RND_CONV_false_1_e_dif1_nand_3_nl
      , 1'b1});
  assign acc_14_nl = nl_acc_14_nl[12:0];
  assign z_out_25 = readslicef_13_12_1(acc_14_nl);
  assign return_add_generic_AC_RND_CONV_false_8_e_dif1_mux_4_nl = MUX_v_11_2_2((~
      return_mult_generic_AC_RND_CONV_false_2_exp_1_11_0_lpi_3_dfm_3_10_0_1), (~
      return_mult_generic_AC_RND_CONV_false_5_exp_1_11_0_lpi_3_dfm_3_10_0_1), fsm_output[39]);
  assign nl_acc_15_nl = ({1'b1 , BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1 , reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd
      , reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1 , 1'b1}) + conv_u2u_12_13({return_add_generic_AC_RND_CONV_false_8_e_dif1_mux_4_nl
      , 1'b1});
  assign acc_15_nl = nl_acc_15_nl[12:0];
  assign z_out_26 = readslicef_13_12_1(acc_15_nl);
  assign return_mult_generic_AC_RND_CONV_false_exp_return_mult_generic_AC_RND_CONV_false_exp_and_1_nl
      = (z_out_44[11]) & (~((fsm_output[10]) | (fsm_output[12]) | (fsm_output[35])
      | (fsm_output[37]) | (fsm_output[54])));
  assign return_mult_generic_AC_RND_CONV_false_exp_mux1h_12_nl = MUX1HOT_v_6_6_2(stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_5,
      stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5, (z_out_44[10:5]), stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_10_5,
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_10_5, (out_f_d_rsci_q_d[62:57]),
      {(fsm_output[10]) , (fsm_output[12]) , BUTTERFLY_i_or_4_cse , (fsm_output[35])
      , (fsm_output[37]) , (fsm_output[54])});
  assign return_mult_generic_AC_RND_CONV_false_exp_mux1h_13_nl = MUX1HOT_v_4_6_2(stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_4_1,
      stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1, (z_out_44[4:1]), stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_4_1,
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_4_1, (out_f_d_rsci_q_d[56:53]), {(fsm_output[10])
      , (fsm_output[12]) , BUTTERFLY_i_or_4_cse , (fsm_output[35]) , (fsm_output[37])
      , (fsm_output[54])});
  assign return_mult_generic_AC_RND_CONV_false_exp_mux1h_14_nl = MUX1HOT_s_1_6_2(stage_PE_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0,
      stage_PE_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0, (z_out_44[0]), stage_PE_1_tmp_re_d_1_lpi_3_dfm_62_52_mx0_0,
      stage_PE_1_tmp_im_d_1_lpi_3_dfm_62_52_mx0_0, (out_f_d_rsci_q_d[52]), {(fsm_output[10])
      , (fsm_output[12]) , BUTTERFLY_i_or_4_cse , (fsm_output[35]) , (fsm_output[37])
      , (fsm_output[54])});
  assign return_mult_generic_AC_RND_CONV_false_exp_mux1h_15_nl = MUX1HOT_s_1_4_2(return_extract_15_return_extract_15_nor_cse_sva,
      return_extract_17_return_extract_17_nor_cse_sva, return_extract_19_return_extract_19_nor_tmp,
      return_extract_51_return_extract_51_nor_tmp, {or_dcpl_548 , or_dcpl_404 , (fsm_output[14])
      , (fsm_output[39])});
  assign return_mult_generic_AC_RND_CONV_false_exp_or_12_nl = return_mult_generic_AC_RND_CONV_false_exp_mux1h_15_nl
      | (fsm_output[54]);
  assign return_mult_generic_AC_RND_CONV_false_exp_or_13_nl = (fsm_output[14]) |
      (fsm_output[39]) | (fsm_output[54]);
  assign return_mult_generic_AC_RND_CONV_false_exp_return_mult_generic_AC_RND_CONV_false_exp_or_1_nl
      = MUX_v_2_2_2((z_out_39[11:10]), 2'b11, return_mult_generic_AC_RND_CONV_false_exp_or_13_nl);
  assign return_mult_generic_AC_RND_CONV_false_exp_mux1h_16_nl = MUX1HOT_v_9_3_2((z_out_39[9:1]),
      (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[61:53]), 9'b111111011, {return_mult_generic_AC_RND_CONV_false_exp_or_4_itm
      , BUTTERFLY_i_or_4_cse , (fsm_output[54])});
  assign return_mult_generic_AC_RND_CONV_false_exp_mux1h_17_nl = MUX1HOT_s_1_3_2((z_out_39[0]),
      (stage_PE_1_gm_im_d_61_0_lpi_3_dfm[52]), (~ return_add_generic_AC_RND_CONV_false_10_return_add_generic_AC_RND_CONV_false_10_or_tmp),
      {return_mult_generic_AC_RND_CONV_false_exp_or_4_itm , BUTTERFLY_i_or_4_cse
      , (fsm_output[54])});
  assign nl_acc_16_nl = conv_u2u_13_14({return_mult_generic_AC_RND_CONV_false_exp_return_mult_generic_AC_RND_CONV_false_exp_and_1_nl
      , return_mult_generic_AC_RND_CONV_false_exp_mux1h_12_nl , return_mult_generic_AC_RND_CONV_false_exp_mux1h_13_nl
      , return_mult_generic_AC_RND_CONV_false_exp_mux1h_14_nl , return_mult_generic_AC_RND_CONV_false_exp_or_12_nl})
      + conv_s2u_13_14({return_mult_generic_AC_RND_CONV_false_exp_return_mult_generic_AC_RND_CONV_false_exp_or_1_nl
      , return_mult_generic_AC_RND_CONV_false_exp_mux1h_16_nl , return_mult_generic_AC_RND_CONV_false_exp_mux1h_17_nl
      , 1'b1});
  assign acc_16_nl = nl_acc_16_nl[13:0];
  assign z_out_27 = readslicef_14_13_1(acc_16_nl);
  assign operator_6_false_9_mux_4_nl = MUX_s_1_2_2((drf_qr_lval_4_smx_9_0_lpi_3_dfm_mx0[9]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd, or_38_cse);
  assign operator_6_false_9_mux_5_nl = MUX_v_4_2_2((drf_qr_lval_4_smx_9_0_lpi_3_dfm_mx0[8:5]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1, or_38_cse);
  assign operator_6_false_9_mux_6_nl = MUX_v_4_2_2((drf_qr_lval_4_smx_9_0_lpi_3_dfm_mx0[4:1]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2, or_38_cse);
  assign operator_6_false_9_mux_7_nl = MUX_s_1_2_2((drf_qr_lval_4_smx_9_0_lpi_3_dfm_mx0[0]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3, or_38_cse);
  assign nl_acc_17_nl = conv_u2u_11_12({operator_6_false_9_mux_4_nl , operator_6_false_9_mux_5_nl
      , operator_6_false_9_mux_6_nl , operator_6_false_9_mux_7_nl , 1'b1}) + conv_s2u_8_12({1'b1
      , (~ rtn_out) , 1'b1});
  assign acc_17_nl = nl_acc_17_nl[11:0];
  assign z_out_28 = readslicef_12_11_1(acc_17_nl);
  assign operator_6_false_14_operator_6_false_14_mux_2_nl = MUX_s_1_2_2((z_out_27[12]),
      (z_out_27[11]), fsm_output[54]);
  assign nl_acc_18_nl = ({operator_6_false_14_operator_6_false_14_mux_2_nl , (z_out_27[11:0])
      , 1'b1}) + conv_s2u_8_14({1'b1 , (~ rtn_out_1) , 1'b1});
  assign acc_18_nl = nl_acc_18_nl[13:0];
  assign z_out_29 = readslicef_14_13_1(acc_18_nl);
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_25_nl = MUX1HOT_v_45_13_2((return_add_generic_AC_RND_CONV_false_4_mux_24_cse[55:11]),
      (return_add_generic_AC_RND_CONV_false_5_mux_18_cse[55:11]), (return_add_generic_AC_RND_CONV_false_res_mant_conc_2_itm_56_1[55:11]),
      (return_add_generic_AC_RND_CONV_false_5_mux_19_cse[55:11]), (return_add_generic_AC_RND_CONV_false_12_mux_19_cse[55:11]),
      (return_add_generic_AC_RND_CONV_false_1_res_mant_conc_2_itm_56_1[55:11]), (return_add_generic_AC_RND_CONV_false_5_mux_20_cse[55:11]),
      (return_add_generic_AC_RND_CONV_false_6_mux_33_cse[55:11]), (return_add_generic_AC_RND_CONV_false_8_res_mant_conc_7_itm_56_1[55:11]),
      (return_add_generic_AC_RND_CONV_false_14_res_mant_conc_2_itm_56_1[55:11]),
      (return_add_generic_AC_RND_CONV_false_12_mux_21_cse[55:11]), (return_add_generic_AC_RND_CONV_false_13_res_mant_conc_2_itm_56_1[55:11]),
      (signext_45_11(z_out_25[10:0])), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_4_or_35_cse , (fsm_output[5]) , return_add_generic_AC_RND_CONV_false_4_or_33_cse
      , return_add_generic_AC_RND_CONV_false_4_or_43_cse , (fsm_output[7]) , return_add_generic_AC_RND_CONV_false_4_or_47_cse
      , or_dcpl_404 , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse
      , (fsm_output[32]) , return_add_generic_AC_RND_CONV_false_12_res_mant_or_cse
      , (fsm_output[30]) , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_26_nl = MUX1HOT_v_11_13_2((return_add_generic_AC_RND_CONV_false_4_mux_24_cse[10:0]),
      (return_add_generic_AC_RND_CONV_false_5_mux_18_cse[10:0]), (return_add_generic_AC_RND_CONV_false_res_mant_conc_2_itm_56_1[10:0]),
      (return_add_generic_AC_RND_CONV_false_5_mux_19_cse[10:0]), (return_add_generic_AC_RND_CONV_false_12_mux_19_cse[10:0]),
      (return_add_generic_AC_RND_CONV_false_1_res_mant_conc_2_itm_56_1[10:0]), (return_add_generic_AC_RND_CONV_false_5_mux_20_cse[10:0]),
      (return_add_generic_AC_RND_CONV_false_6_mux_33_cse[10:0]), (return_add_generic_AC_RND_CONV_false_8_res_mant_conc_7_itm_56_1[10:0]),
      (return_add_generic_AC_RND_CONV_false_14_res_mant_conc_2_itm_56_1[10:0]), (return_add_generic_AC_RND_CONV_false_12_mux_21_cse[10:0]),
      (return_add_generic_AC_RND_CONV_false_13_res_mant_conc_2_itm_56_1[10:0]), (in_u_rsci_q_d[11:1]),
      {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , return_add_generic_AC_RND_CONV_false_4_or_35_cse
      , (fsm_output[5]) , return_add_generic_AC_RND_CONV_false_4_or_33_cse , return_add_generic_AC_RND_CONV_false_4_or_43_cse
      , (fsm_output[7]) , return_add_generic_AC_RND_CONV_false_4_or_47_cse , or_dcpl_404
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse , (fsm_output[32])
      , return_add_generic_AC_RND_CONV_false_12_res_mant_or_cse , (fsm_output[30])
      , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_4_and_137_nl = (~ return_add_generic_AC_RND_CONV_false_17_do_sub_sva_1)
      & (fsm_output[3]);
  assign return_add_generic_AC_RND_CONV_false_4_and_138_nl = return_add_generic_AC_RND_CONV_false_17_do_sub_sva_1
      & (fsm_output[3]);
  assign return_add_generic_AC_RND_CONV_false_4_and_139_nl = (~ return_add_generic_AC_RND_CONV_false_10_do_sub_sva)
      & or_38_cse;
  assign return_add_generic_AC_RND_CONV_false_4_and_140_nl = return_add_generic_AC_RND_CONV_false_10_do_sub_sva
      & or_38_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_117_nl = or_dcpl_401 | (fsm_output[17])
      | (fsm_output[19]) | return_extract_26_exception_or_3_cse | (fsm_output[42])
      | (fsm_output[44]) | return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse;
  assign return_add_generic_AC_RND_CONV_false_4_and_141_nl = (~ return_add_generic_AC_RND_CONV_false_10_do_sub_sva)
      & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_4_and_142_nl = return_add_generic_AC_RND_CONV_false_10_do_sub_sva
      & (fsm_output[43]);
  assign return_add_generic_AC_RND_CONV_false_4_and_143_nl = (~ not_tmp_302) & (fsm_output[12]);
  assign return_add_generic_AC_RND_CONV_false_4_and_144_nl = not_tmp_302 & (fsm_output[12]);
  assign return_add_generic_AC_RND_CONV_false_4_and_145_nl = (~ return_add_generic_AC_RND_CONV_false_14_op2_inf_sva)
      & return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse;
  assign return_add_generic_AC_RND_CONV_false_4_and_146_nl = return_add_generic_AC_RND_CONV_false_14_op2_inf_sva
      & return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse;
  assign return_add_generic_AC_RND_CONV_false_4_and_147_nl = (~ return_add_generic_AC_RND_CONV_false_10_do_sub_sva)
      & (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_4_and_148_nl = return_add_generic_AC_RND_CONV_false_10_do_sub_sva
      & (fsm_output[18]);
  assign return_add_generic_AC_RND_CONV_false_4_and_149_nl = (~ not_tmp_302) & (fsm_output[37]);
  assign return_add_generic_AC_RND_CONV_false_4_and_150_nl = not_tmp_302 & (fsm_output[37]);
  assign return_add_generic_AC_RND_CONV_false_4_and_151_nl = (~ return_add_generic_AC_RND_CONV_false_12_do_sub_sva)
      & (fsm_output[20]);
  assign return_add_generic_AC_RND_CONV_false_4_and_152_nl = return_add_generic_AC_RND_CONV_false_12_do_sub_sva
      & (fsm_output[20]);
  assign return_add_generic_AC_RND_CONV_false_4_and_153_nl = (~ return_add_generic_AC_RND_CONV_false_12_do_sub_sva)
      & (fsm_output[45]);
  assign return_add_generic_AC_RND_CONV_false_4_and_154_nl = return_add_generic_AC_RND_CONV_false_12_do_sub_sva
      & (fsm_output[45]);
  assign return_add_generic_AC_RND_CONV_false_4_and_155_nl = (~ return_add_generic_AC_RND_CONV_false_17_do_sub_sva_1)
      & (fsm_output[28]);
  assign return_add_generic_AC_RND_CONV_false_4_and_156_nl = return_add_generic_AC_RND_CONV_false_17_do_sub_sva_1
      & (fsm_output[28]);
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_27_nl = MUX1HOT_s_1_30_2(return_add_generic_AC_RND_CONV_false_4_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_4_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_5_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_5_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_res_mant_3_0_sva_1,
      (~ return_add_generic_AC_RND_CONV_false_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_11_mux_2_itm,
      return_add_generic_AC_RND_CONV_false_23_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_23_res_mant_3_0_sva_1),
      return_add_generic_AC_RND_CONV_false_1_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_1_res_mant_3_0_sva_1),
      (~ return_add_generic_AC_RND_CONV_false_6_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_6_res_mant_3_0_sva_1,
      return_add_generic_AC_RND_CONV_false_8_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_8_res_mant_3_0_sva_1),
      return_add_generic_AC_RND_CONV_false_10_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_10_res_mant_3_0_sva_1),
      return_add_generic_AC_RND_CONV_false_14_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_14_res_mant_3_0_sva_1),
      (~ return_add_generic_AC_RND_CONV_false_19_res_mant_3_0_sva_1), return_add_generic_AC_RND_CONV_false_19_res_mant_3_0_sva_1,
      return_add_generic_AC_RND_CONV_false_12_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_12_res_mant_3_0_sva_1),
      return_add_generic_AC_RND_CONV_false_25_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_25_res_mant_3_0_sva_1),
      return_add_generic_AC_RND_CONV_false_17_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_17_res_mant_3_0_sva_1),
      return_add_generic_AC_RND_CONV_false_13_res_mant_3_0_sva_1, (~ return_add_generic_AC_RND_CONV_false_13_res_mant_3_0_sva_1),
      (in_u_rsci_q_d[0]), {return_add_generic_AC_RND_CONV_false_4_and_137_nl , return_add_generic_AC_RND_CONV_false_4_and_138_nl
      , return_add_generic_AC_RND_CONV_false_4_and_139_nl , return_add_generic_AC_RND_CONV_false_4_and_140_nl
      , return_add_generic_AC_RND_CONV_false_11_and_3_cse , return_add_generic_AC_RND_CONV_false_11_and_4_cse
      , return_add_generic_AC_RND_CONV_false_4_or_117_nl , return_add_generic_AC_RND_CONV_false_4_and_141_nl
      , return_add_generic_AC_RND_CONV_false_4_and_142_nl , return_add_generic_AC_RND_CONV_false_11_and_5_cse
      , return_add_generic_AC_RND_CONV_false_11_and_6_cse , return_add_generic_AC_RND_CONV_false_4_and_143_nl
      , return_add_generic_AC_RND_CONV_false_4_and_144_nl , return_add_generic_AC_RND_CONV_false_4_and_145_nl
      , return_add_generic_AC_RND_CONV_false_4_and_146_nl , return_add_generic_AC_RND_CONV_false_4_and_147_nl
      , return_add_generic_AC_RND_CONV_false_4_and_148_nl , return_add_generic_AC_RND_CONV_false_11_and_15_cse
      , return_add_generic_AC_RND_CONV_false_11_and_16_cse , return_add_generic_AC_RND_CONV_false_4_and_149_nl
      , return_add_generic_AC_RND_CONV_false_4_and_150_nl , return_add_generic_AC_RND_CONV_false_4_and_151_nl
      , return_add_generic_AC_RND_CONV_false_4_and_152_nl , return_add_generic_AC_RND_CONV_false_4_and_153_nl
      , return_add_generic_AC_RND_CONV_false_4_and_154_nl , return_add_generic_AC_RND_CONV_false_4_and_155_nl
      , return_add_generic_AC_RND_CONV_false_4_and_156_nl , return_add_generic_AC_RND_CONV_false_11_and_13_cse
      , return_add_generic_AC_RND_CONV_false_11_and_14_cse , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_28_nl = MUX1HOT_s_1_12_2(return_add_generic_AC_RND_CONV_false_17_do_sub_sva_1,
      return_add_generic_AC_RND_CONV_false_10_do_sub_sva, xor_cse, return_add_generic_AC_RND_CONV_false_11_do_sub_sva,
      return_add_generic_AC_RND_CONV_false_14_op2_nan_sva, xor_2_cse, return_add_generic_AC_RND_CONV_false_16_do_sub_sva,
      return_add_generic_AC_RND_CONV_false_6_do_sub_sva_1, return_add_generic_AC_RND_CONV_false_14_op2_inf_sva,
      xor_4_cse, return_add_generic_AC_RND_CONV_false_12_do_sub_sva, xor_3_cse, {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_4_or_35_cse , (fsm_output[5]) , return_add_generic_AC_RND_CONV_false_4_or_33_cse
      , return_add_generic_AC_RND_CONV_false_4_or_43_cse , (fsm_output[7]) , return_add_generic_AC_RND_CONV_false_4_or_47_cse
      , or_dcpl_404 , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse
      , (fsm_output[32]) , return_add_generic_AC_RND_CONV_false_12_res_mant_or_cse
      , (fsm_output[30])});
  assign return_add_generic_AC_RND_CONV_false_4_and_157_nl = return_add_generic_AC_RND_CONV_false_4_mux1h_28_nl
      & (~ (fsm_output[54]));
  assign return_add_generic_AC_RND_CONV_false_4_or_121_nl = and_1583_cse | return_add_generic_AC_RND_CONV_false_4_and_69_cse
      | return_add_generic_AC_RND_CONV_false_4_and_73_cse | return_add_generic_AC_RND_CONV_false_4_and_75_cse
      | and_1584_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_122_nl = or_dcpl_401 | return_extract_26_exception_or_3_cse
      | return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_123_nl = return_add_generic_AC_RND_CONV_false_4_and_67_cse
      | return_add_generic_AC_RND_CONV_false_4_and_71_cse;
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_29_nl = MUX1HOT_s_1_16_2(return_add_generic_AC_RND_CONV_false_17_op1_mu_52_lpi_3_dfm_1,
      stage_PE_1_gm_im_d_mux_cse, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm,
      return_add_generic_AC_RND_CONV_false_op2_mu_52_lpi_3_dfm_1, drf_qr_lval_13_smx_0_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm, return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_itm,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm, return_add_generic_AC_RND_CONV_false_13_slc_return_add_generic_AC_RND_CONV_false_13_res_rounded_51_0_itm,
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_52_lpi_3_dfm_mx0, return_add_generic_AC_RND_CONV_false_6_op2_mu_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm, return_add_generic_AC_RND_CONV_false_10_op2_mu_1_52_lpi_3_dfm_mx0,
      return_add_generic_AC_RND_CONV_false_13_op1_mu_52_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm,
      return_add_generic_AC_RND_CONV_false_19_op2_mu_52_lpi_3_dfm_mx0, {return_add_generic_AC_RND_CONV_false_4_and_105_cse
      , and_1153_rgt , or_38_cse , return_add_generic_AC_RND_CONV_false_4_or_70_cse
      , return_add_generic_AC_RND_CONV_false_4_or_121_nl , return_add_generic_AC_RND_CONV_false_4_or_122_nl
      , return_extract_1_exception_or_cse , return_add_generic_AC_RND_CONV_false_10_or_cse
      , return_add_generic_AC_RND_CONV_false_4_or_123_nl , and_1163_cse , or_1673_ssc
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse , and_2281_cse
      , return_add_generic_AC_RND_CONV_false_4_or_73_cse , return_add_generic_AC_RND_CONV_false_4_and_77_cse
      , or_1678_ssc});
  assign return_add_generic_AC_RND_CONV_false_4_and_158_nl = return_add_generic_AC_RND_CONV_false_4_mux1h_29_nl
      & (~ (fsm_output[54]));
  assign return_add_generic_AC_RND_CONV_false_4_or_124_nl = return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse
      | return_add_generic_AC_RND_CONV_false_4_and_77_cse;
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_30_nl = MUX1HOT_s_1_17_2((z_out_11[50]),
      return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_0, (return_add_generic_AC_RND_CONV_false_conc_6_itm_54_4[50]),
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_1_itm, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm,
      (return_add_generic_AC_RND_CONV_false_10_slc_return_add_generic_AC_RND_CONV_false_10_res_rounded_51_0_1_itm[50]),
      return_add_generic_AC_RND_CONV_false_23_op2_mu_1_51_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_1_conc_6_itm_54_4[50]),
      return_add_generic_AC_RND_CONV_false_11_op_smaller_qr_52_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_6_op2_mu_51_1_lpi_3_dfm_50_mx0,
      return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm, (return_add_generic_AC_RND_CONV_false_13_op2_mu_51_1_lpi_3_dfm[50]),
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_51_lpi_3_dfm_mx0, (return_add_generic_AC_RND_CONV_false_14_conc_6_itm_54_4[50]),
      return_add_generic_AC_RND_CONV_false_19_op2_mu_51_1_lpi_3_dfm_50_mx0, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm,
      (return_add_generic_AC_RND_CONV_false_13_conc_6_itm_54_4[50]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_4_or_99_cse , (fsm_output[5]) , return_extract_1_exception_or_cse
      , return_add_generic_AC_RND_CONV_false_10_or_cse , return_add_generic_AC_RND_CONV_false_4_and_67_cse
      , and_1163_cse , (fsm_output[7]) , return_add_generic_AC_RND_CONV_false_4_and_71_cse
      , or_1673_ssc , return_add_generic_AC_RND_CONV_false_4_or_124_nl , return_add_generic_AC_RND_CONV_false_4_and_73_cse
      , and_2281_cse , (fsm_output[32]) , or_1678_ssc , return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
      , (fsm_output[30])});
  assign return_add_generic_AC_RND_CONV_false_4_and_159_nl = return_add_generic_AC_RND_CONV_false_4_mux1h_30_nl
      & (~ (fsm_output[54]));
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_31_nl = MUX1HOT_v_30_12_2((z_out_11[49:20]),
      (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[49:20]),
      (return_add_generic_AC_RND_CONV_false_conc_6_itm_54_4[49:20]), (return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm[49:20]),
      (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_49_0[49:20]), (return_add_generic_AC_RND_CONV_false_23_conc_6_itm_53_4[49:20]),
      (return_add_generic_AC_RND_CONV_false_1_conc_6_itm_54_4[49:20]), (return_add_generic_AC_RND_CONV_false_6_conc_6_itm_53_4[49:20]),
      (return_add_generic_AC_RND_CONV_false_10_conc_6_itm_53_4[49:20]), (return_add_generic_AC_RND_CONV_false_14_conc_6_itm_54_4[49:20]),
      (return_add_generic_AC_RND_CONV_false_19_conc_6_itm_53_4[49:20]), (return_add_generic_AC_RND_CONV_false_13_conc_6_itm_54_4[49:20]),
      {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , return_add_generic_AC_RND_CONV_false_4_or_99_cse
      , (fsm_output[5]) , return_add_generic_AC_RND_CONV_false_4_or_27_cse , return_add_generic_AC_RND_CONV_false_4_or_31_cse
      , (fsm_output[43]) , (fsm_output[7]) , (fsm_output[12]) , (fsm_output[18])
      , (fsm_output[32]) , (fsm_output[37]) , (fsm_output[30])});
  assign return_add_generic_AC_RND_CONV_false_4_not_59_nl = ~ (fsm_output[54]);
  assign return_add_generic_AC_RND_CONV_false_4_and_160_nl = MUX_v_30_2_2(30'b000000000000000000000000000000,
      return_add_generic_AC_RND_CONV_false_4_mux1h_31_nl, return_add_generic_AC_RND_CONV_false_4_not_59_nl);
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_32_nl = MUX1HOT_v_10_13_2((z_out_11[19:10]),
      (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[19:10]),
      (return_add_generic_AC_RND_CONV_false_conc_6_itm_54_4[19:10]), (return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm[19:10]),
      (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_49_0[19:10]), (return_add_generic_AC_RND_CONV_false_23_conc_6_itm_53_4[19:10]),
      (return_add_generic_AC_RND_CONV_false_1_conc_6_itm_54_4[19:10]), (return_add_generic_AC_RND_CONV_false_6_conc_6_itm_53_4[19:10]),
      (return_add_generic_AC_RND_CONV_false_10_conc_6_itm_53_4[19:10]), (return_add_generic_AC_RND_CONV_false_14_conc_6_itm_54_4[19:10]),
      (return_add_generic_AC_RND_CONV_false_19_conc_6_itm_53_4[19:10]), (return_add_generic_AC_RND_CONV_false_13_conc_6_itm_54_4[19:10]),
      (z_out_19[9:0]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_4_or_99_cse , (fsm_output[5]) , return_add_generic_AC_RND_CONV_false_4_or_27_cse
      , return_add_generic_AC_RND_CONV_false_4_or_31_cse , (fsm_output[43]) , (fsm_output[7])
      , (fsm_output[12]) , (fsm_output[18]) , (fsm_output[32]) , (fsm_output[37])
      , (fsm_output[30]) , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_33_nl = MUX1HOT_v_4_12_2((z_out_11[9:6]),
      (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[9:6]), (return_add_generic_AC_RND_CONV_false_conc_6_itm_54_4[9:6]),
      (return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm[9:6]), (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_49_0[9:6]),
      (return_add_generic_AC_RND_CONV_false_23_conc_6_itm_53_4[9:6]), (return_add_generic_AC_RND_CONV_false_1_conc_6_itm_54_4[9:6]),
      (return_add_generic_AC_RND_CONV_false_6_conc_6_itm_53_4[9:6]), (return_add_generic_AC_RND_CONV_false_10_conc_6_itm_53_4[9:6]),
      (return_add_generic_AC_RND_CONV_false_14_conc_6_itm_54_4[9:6]), (return_add_generic_AC_RND_CONV_false_19_conc_6_itm_53_4[9:6]),
      (return_add_generic_AC_RND_CONV_false_13_conc_6_itm_54_4[9:6]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , return_add_generic_AC_RND_CONV_false_4_or_99_cse , (fsm_output[5]) , return_add_generic_AC_RND_CONV_false_4_or_27_cse
      , return_add_generic_AC_RND_CONV_false_4_or_31_cse , (fsm_output[43]) , (fsm_output[7])
      , (fsm_output[12]) , (fsm_output[18]) , (fsm_output[32]) , (fsm_output[37])
      , (fsm_output[30])});
  assign return_add_generic_AC_RND_CONV_false_4_not_60_nl = ~ (fsm_output[54]);
  assign return_add_generic_AC_RND_CONV_false_4_and_161_nl = MUX_v_4_2_2(4'b0000,
      return_add_generic_AC_RND_CONV_false_4_mux1h_33_nl, return_add_generic_AC_RND_CONV_false_4_not_60_nl);
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_34_nl = MUX1HOT_v_6_13_2((z_out_11[5:0]),
      (return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1[5:0]), (return_add_generic_AC_RND_CONV_false_conc_6_itm_54_4[5:0]),
      (return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_2_itm[5:0]), (return_add_generic_AC_RND_CONV_false_12_res_mant_4_sva_49_0[5:0]),
      (return_add_generic_AC_RND_CONV_false_23_conc_6_itm_53_4[5:0]), (return_add_generic_AC_RND_CONV_false_1_conc_6_itm_54_4[5:0]),
      (return_add_generic_AC_RND_CONV_false_6_conc_6_itm_53_4[5:0]), (return_add_generic_AC_RND_CONV_false_10_conc_6_itm_53_4[5:0]),
      (return_add_generic_AC_RND_CONV_false_14_conc_6_itm_54_4[5:0]), (return_add_generic_AC_RND_CONV_false_19_conc_6_itm_53_4[5:0]),
      (return_add_generic_AC_RND_CONV_false_13_conc_6_itm_54_4[5:0]), (z_out_19[9:4]),
      {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse , return_add_generic_AC_RND_CONV_false_4_or_99_cse
      , (fsm_output[5]) , return_add_generic_AC_RND_CONV_false_4_or_27_cse , return_add_generic_AC_RND_CONV_false_4_or_31_cse
      , (fsm_output[43]) , (fsm_output[7]) , (fsm_output[12]) , (fsm_output[18])
      , (fsm_output[32]) , (fsm_output[37]) , (fsm_output[30]) , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_4_or_125_nl = or_dcpl_401 | (fsm_output[19])
      | return_extract_26_exception_or_3_cse | (fsm_output[42]) | (fsm_output[45]);
  assign return_add_generic_AC_RND_CONV_false_4_or_126_nl = (fsm_output[17]) | (fsm_output[44])
      | (fsm_output[20]) | return_add_generic_AC_RND_CONV_false_4_and_71_cse;
  assign return_add_generic_AC_RND_CONV_false_4_or_127_nl = return_add_generic_AC_RND_CONV_false_4_and_67_cse
      | return_add_generic_AC_RND_CONV_false_4_and_69_cse | return_add_generic_AC_RND_CONV_false_4_and_73_cse
      | return_add_generic_AC_RND_CONV_false_4_and_75_cse;
  assign return_add_generic_AC_RND_CONV_false_4_mux1h_35_nl = MUX1HOT_s_1_17_2(return_add_generic_AC_RND_CONV_false_17_op1_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_17_op2_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_1_itm,
      return_add_generic_AC_RND_CONV_false_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_op2_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_3_itm, return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_3_itm,
      return_add_generic_AC_RND_CONV_false_1_op1_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_23_op2_mu_1_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_6_op2_mu_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_12_op_bigger_mux_itm,
      return_add_generic_AC_RND_CONV_false_10_op2_mu_1_0_lpi_3_dfm_1, return_add_generic_AC_RND_CONV_false_13_op1_mu_0_lpi_3_dfm_1,
      drf_qr_lval_13_smx_0_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_19_op2_mu_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_11_op_bigger_mux_itm, (z_out_19[3]), {return_add_generic_AC_RND_CONV_false_4_and_105_cse
      , and_1153_rgt , or_38_cse , return_add_generic_AC_RND_CONV_false_4_or_70_cse
      , or_tmp_561 , return_add_generic_AC_RND_CONV_false_4_or_125_nl , return_add_generic_AC_RND_CONV_false_4_or_126_nl
      , return_add_generic_AC_RND_CONV_false_4_or_127_nl , and_1163_cse , or_1673_ssc
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse , and_2281_cse
      , return_add_generic_AC_RND_CONV_false_4_or_73_cse , return_add_generic_AC_RND_CONV_false_4_and_77_cse
      , or_1678_ssc , return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
      , (fsm_output[54])});
  assign return_add_generic_AC_RND_CONV_false_4_nor_1_nl = ~((fsm_output[3]) | or_38_cse
      | (fsm_output[5]) | or_dcpl_401 | (fsm_output[17]) | (fsm_output[19]) | (fsm_output[43])
      | (fsm_output[7]) | return_extract_26_exception_or_3_cse | (fsm_output[12])
      | return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_4_cse | (fsm_output[18])
      | (fsm_output[32]) | (fsm_output[37]) | (fsm_output[42]) | (fsm_output[44])
      | (fsm_output[20]) | (fsm_output[45]) | return_add_generic_AC_RND_CONV_false_15_res_rounded_or_1_cse
      | (fsm_output[28]) | (fsm_output[30]));
  assign return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_8_nl
      = MUX_v_3_2_2(3'b000, (z_out_19[2:0]), return_add_generic_AC_RND_CONV_false_4_nor_1_nl);
  assign nl_acc_19_nl = ({return_add_generic_AC_RND_CONV_false_4_mux1h_25_nl , return_add_generic_AC_RND_CONV_false_4_mux1h_26_nl
      , return_add_generic_AC_RND_CONV_false_4_mux1h_27_nl , return_add_generic_AC_RND_CONV_false_4_and_157_nl})
      + conv_u2u_57_58({return_add_generic_AC_RND_CONV_false_4_and_158_nl , return_add_generic_AC_RND_CONV_false_4_and_159_nl
      , return_add_generic_AC_RND_CONV_false_4_and_160_nl , return_add_generic_AC_RND_CONV_false_4_mux1h_32_nl
      , return_add_generic_AC_RND_CONV_false_4_and_161_nl , return_add_generic_AC_RND_CONV_false_4_mux1h_34_nl
      , return_add_generic_AC_RND_CONV_false_4_mux1h_35_nl , return_add_generic_AC_RND_CONV_false_4_return_add_generic_AC_RND_CONV_false_4_and_8_nl
      , 1'b1});
  assign acc_19_nl = nl_acc_19_nl[57:0];
  assign z_out_30 = readslicef_58_57_1(acc_19_nl);
  assign nl_acc_20_nl = ({1'b1 , drf_qr_lval_14_smx_0_lpi_3_dfm , return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_0
      , return_add_generic_AC_RND_CONV_false_15_op_bigger_mux_2_itm_rsp_1 , 1'b1})
      + conv_u2u_53_54({return_add_generic_AC_RND_CONV_false_20_ma1_lt_ma2_mux_1_cse
      , return_add_generic_AC_RND_CONV_false_20_ma1_lt_ma2_mux_4_cse , 1'b1});
  assign acc_20_nl = nl_acc_20_nl[53:0];
  assign z_out_31_52 = readslicef_54_1_53(acc_20_nl);
  assign return_add_generic_AC_RND_CONV_false_6_ma1_lt_ma2_mux_5_nl = MUX_s_1_2_2((~
      return_add_generic_AC_RND_CONV_false_3_r_nan_mux1h_cse), (~ return_add_generic_AC_RND_CONV_false_16_r_nan_mux1h_cse),
      fsm_output[37]);
  assign return_add_generic_AC_RND_CONV_false_6_ma1_lt_ma2_mux_6_nl = MUX_v_51_2_2((~
      stage_PE_tmp_im_d_1_lpi_3_dfm_50_0_mx0), (~ stage_PE_1_tmp_im_d_1_lpi_3_dfm_50_0_mx0),
      fsm_output[37]);
  assign nl_acc_21_nl = ({1'b1 , return_extract_15_return_extract_15_nor_cse_sva
      , stage_PE_1_tmp_re_d_1_sva_1_56_0_rsp_1 , 1'b1}) + conv_u2u_53_54({return_add_generic_AC_RND_CONV_false_6_ma1_lt_ma2_mux_5_nl
      , return_add_generic_AC_RND_CONV_false_6_ma1_lt_ma2_mux_6_nl , 1'b1});
  assign acc_21_nl = nl_acc_21_nl[53:0];
  assign z_out_32_52 = readslicef_54_1_53(acc_21_nl);
  assign return_add_generic_AC_RND_CONV_false_9_ma1_lt_ma2_mux_4_nl = MUX_s_1_2_2((~
      return_add_generic_AC_RND_CONV_false_7_m_r_51_lpi_3_dfm_mx0), (~ return_add_generic_AC_RND_CONV_false_20_m_r_51_lpi_3_dfm_mx0),
      fsm_output[41]);
  assign return_add_generic_AC_RND_CONV_false_9_ma1_lt_ma2_mux_5_nl = MUX_v_51_2_2((~
      return_add_generic_AC_RND_CONV_false_7_m_r_50_0_lpi_3_dfm_1), (~ return_add_generic_AC_RND_CONV_false_20_m_r_50_0_lpi_3_dfm_1),
      fsm_output[41]);
  assign nl_acc_22_nl = ({1'b1 , (stage_PE_1_x_re_d_sva[51:0]) , 1'b1}) + conv_u2u_53_54({return_add_generic_AC_RND_CONV_false_9_ma1_lt_ma2_mux_4_nl
      , return_add_generic_AC_RND_CONV_false_9_ma1_lt_ma2_mux_5_nl , 1'b1});
  assign acc_22_nl = nl_acc_22_nl[53:0];
  assign z_out_33_52 = readslicef_54_1_53(acc_22_nl);
  assign return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_mux1h_4_nl = MUX1HOT_s_1_4_2((~
      return_add_generic_AC_RND_CONV_false_21_m_r_51_lpi_3_dfm_mx0), (~ (out_f_d_rsci_q_d[51])),
      (~ return_add_generic_AC_RND_CONV_false_8_m_r_51_lpi_3_dfm_mx0), (~ (in_f_d_rsci_q_d[51])),
      {(fsm_output[43]) , (fsm_output[7]) , (fsm_output[18]) , (fsm_output[32])});
  assign return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_mux1h_5_nl = MUX1HOT_v_51_4_2((~
      return_add_generic_AC_RND_CONV_false_21_m_r_50_0_lpi_3_dfm_1), (~ (out_f_d_rsci_q_d[50:0])),
      (~ return_add_generic_AC_RND_CONV_false_8_m_r_50_0_lpi_3_dfm_1), (~ (in_f_d_rsci_q_d[50:0])),
      {(fsm_output[43]) , (fsm_output[7]) , (fsm_output[18]) , (fsm_output[32])});
  assign nl_acc_23_nl = ({1'b1 , (stage_PE_1_x_im_d_sva[51:0]) , 1'b1}) + conv_u2u_53_54({return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_mux1h_4_nl
      , return_add_generic_AC_RND_CONV_false_23_ma1_lt_ma2_mux1h_5_nl , 1'b1});
  assign acc_23_nl = nl_acc_23_nl[53:0];
  assign z_out_34_52 = readslicef_54_1_53(acc_23_nl);
  assign nl_acc_24_nl = ({1'b1 , return_add_generic_AC_RND_CONV_false_11_mux_2_itm
      , return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_0 , return_add_generic_AC_RND_CONV_false_17_m_r_50_0_lpi_3_dfm_rsp_1
      , 1'b1}) + conv_u2u_53_54({return_add_generic_AC_RND_CONV_false_20_ma1_lt_ma2_mux_1_cse
      , return_add_generic_AC_RND_CONV_false_20_ma1_lt_ma2_mux_4_cse , 1'b1});
  assign acc_24_nl = nl_acc_24_nl[53:0];
  assign z_out_35_52 = readslicef_54_1_53(acc_24_nl);
  assign nl_z_out_36 = return_mult_generic_AC_RND_CONV_false_exp_1_11_0_lpi_3_dfm_1
      + 12'b000000000001;
  assign z_out_36 = nl_z_out_36[11:0];
  assign operator_6_false_8_mux1h_12_nl = MUX1HOT_v_6_5_2((signext_6_1(operator_6_false_8_acc_itm[5])),
      (signext_6_1(exs_26_itm_5_0[5])), BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_0,
      (~ (z_out_45[16:11])), (signext_6_1(exs_27_itm_5_0[5])), {(fsm_output[3]) ,
      or_38_cse , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse
      , (fsm_output[28])});
  assign operator_6_false_8_mux1h_13_nl = MUX1HOT_s_1_5_2((operator_6_false_8_acc_itm[5]),
      (exs_26_itm_5_0[5]), BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_1, (~ (z_out_45[10])),
      (exs_27_itm_5_0[5]), {(fsm_output[3]) , or_38_cse , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse , (fsm_output[28])});
  assign operator_6_false_8_mux1h_14_nl = MUX1HOT_s_1_5_2((operator_6_false_8_acc_itm[5]),
      (exs_26_itm_5_0[5]), reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd, (~ (z_out_45[9])),
      (exs_27_itm_5_0[5]), {(fsm_output[3]) , or_38_cse , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse , (fsm_output[28])});
  assign operator_6_false_8_mux1h_15_nl = MUX1HOT_v_4_5_2((signext_4_2(operator_6_false_8_acc_itm[5:4])),
      (signext_4_2(exs_26_itm_5_0[5:4])), reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1,
      (~ (z_out_45[8:5])), (signext_4_2(exs_27_itm_5_0[5:4])), {(fsm_output[3]) ,
      or_38_cse , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse
      , (fsm_output[28])});
  assign operator_6_false_8_mux1h_16_nl = MUX1HOT_v_4_5_2((operator_6_false_8_acc_itm[3:0]),
      (exs_26_itm_5_0[3:0]), reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2, (~ (z_out_45[4:1])),
      (exs_27_itm_5_0[3:0]), {(fsm_output[3]) , or_38_cse , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse , (fsm_output[28])});
  assign operator_6_false_8_or_3_nl = (fsm_output[3]) | or_38_cse | (fsm_output[28]);
  assign operator_6_false_8_mux1h_17_nl = MUX1HOT_s_1_3_2((~ (rtn_out[0])), reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3,
      (~ (z_out_45[0])), {operator_6_false_8_or_3_nl , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse});
  assign operator_6_false_8_or_4_nl = (~((fsm_output[3]) | or_38_cse | (fsm_output[5])
      | (fsm_output[28]) | (fsm_output[30]))) | return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse;
  assign operator_6_false_8_mux1h_18_nl = MUX1HOT_v_5_3_2((out_u_rsci_q_d[15:11]),
      BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0, (in_u_rsci_q_d[15:11]),
      {(fsm_output[5]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse
      , (fsm_output[30])});
  assign operator_6_false_8_and_2_nl = MUX_v_5_2_2(5'b00000, operator_6_false_8_mux1h_18_nl,
      operator_6_false_8_nor_1_cse);
  assign operator_6_false_8_mux1h_19_nl = MUX1HOT_s_1_3_2((out_u_rsci_q_d[10]), (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1[1]),
      (in_u_rsci_q_d[10]), {(fsm_output[5]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse
      , (fsm_output[30])});
  assign operator_6_false_8_and_3_nl = operator_6_false_8_mux1h_19_nl & operator_6_false_8_nor_1_cse;
  assign operator_6_false_8_mux1h_20_nl = MUX1HOT_s_1_5_2((drf_qr_lval_4_smx_9_0_lpi_3_dfm_mx0[9]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd, (out_u_rsci_q_d[9]), (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1[0]),
      (in_u_rsci_q_d[9]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , or_38_cse , (fsm_output[5]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse
      , (fsm_output[30])});
  assign operator_6_false_8_mux1h_21_nl = MUX1HOT_v_4_5_2((drf_qr_lval_4_smx_9_0_lpi_3_dfm_mx0[8:5]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1, (out_u_rsci_q_d[8:5]), (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[8:5]),
      (in_u_rsci_q_d[8:5]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , or_38_cse , (fsm_output[5]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse
      , (fsm_output[30])});
  assign operator_6_false_8_mux1h_22_nl = MUX1HOT_v_4_5_2((drf_qr_lval_4_smx_9_0_lpi_3_dfm_mx0[4:1]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2, (out_u_rsci_q_d[4:1]), (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[4:1]),
      (in_u_rsci_q_d[4:1]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , or_38_cse , (fsm_output[5]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse
      , (fsm_output[30])});
  assign operator_6_false_8_mux1h_23_nl = MUX1HOT_s_1_5_2((drf_qr_lval_4_smx_9_0_lpi_3_dfm_mx0[0]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3, (out_u_rsci_q_d[0]), (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[0]),
      (in_u_rsci_q_d[0]), {return_add_generic_AC_RND_CONV_false_11_op_bigger_or_3_cse
      , or_38_cse , (fsm_output[5]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_5_cse
      , (fsm_output[30])});
  assign nl_acc_26_nl = conv_s2u_18_19({operator_6_false_8_mux1h_12_nl , operator_6_false_8_mux1h_13_nl
      , operator_6_false_8_mux1h_14_nl , operator_6_false_8_mux1h_15_nl , operator_6_false_8_mux1h_16_nl
      , operator_6_false_8_mux1h_17_nl , operator_6_false_8_or_4_nl}) + conv_u2u_17_19({operator_6_false_8_and_2_nl
      , operator_6_false_8_and_3_nl , operator_6_false_8_mux1h_20_nl , operator_6_false_8_mux1h_21_nl
      , operator_6_false_8_mux1h_22_nl , operator_6_false_8_mux1h_23_nl , 1'b1});
  assign acc_26_nl = nl_acc_26_nl[18:0];
  assign z_out_37 = readslicef_19_18_1(acc_26_nl);
  assign BUTTERFLY_1_else_1_if_BUTTERFLY_1_else_1_if_mux_4_nl = MUX_v_16_2_2((z_out_37[15:0]),
      (z_out_45[15:0]), return_extract_26_exception_or_3_cse);
  assign nl_z_out_38 = BUTTERFLY_1_else_1_if_BUTTERFLY_1_else_1_if_mux_4_nl + conv_u2u_14_16(signext_14_13({BUTTERFLY_1_else_1_if_BUTTERFLY_1_else_1_if_mux_2_cse
      , 11'b00000000000 , BUTTERFLY_1_else_1_if_BUTTERFLY_1_else_1_if_mux_2_cse}));
  assign z_out_38 = nl_z_out_38[15:0];
  assign return_mult_generic_AC_RND_CONV_false_exp_return_mult_generic_AC_RND_CONV_false_exp_mux_4_nl
      = MUX_v_10_2_2(drf_qr_lval_13_smx_10_1_lpi_3_dfm, drf_qr_lval_14_smx_10_1_lpi_3_dfm,
      or_dcpl_404);
  assign return_mult_generic_AC_RND_CONV_false_exp_return_mult_generic_AC_RND_CONV_false_exp_mux_5_nl
      = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_17_e_r_qr_0_lpi_3_dfm, return_add_generic_AC_RND_CONV_false_18_e_r_qr_0_lpi_3_dfm,
      or_dcpl_404);
  assign return_mult_generic_AC_RND_CONV_false_exp_mux1h_18_nl = MUX1HOT_s_1_4_2((~
      return_extract_12_return_extract_12_or_1_cse_sva_1), (~ return_extract_13_return_extract_13_or_1_cse_sva_1),
      (~ return_extract_44_return_extract_44_or_1_cse_sva_1), (~ return_extract_45_return_extract_45_or_1_cse_sva_1),
      {(fsm_output[10]) , (fsm_output[12]) , (fsm_output[35]) , (fsm_output[37])});
  assign nl_acc_28_nl = conv_u2u_12_13({return_mult_generic_AC_RND_CONV_false_exp_return_mult_generic_AC_RND_CONV_false_exp_mux_4_nl
      , return_mult_generic_AC_RND_CONV_false_exp_return_mult_generic_AC_RND_CONV_false_exp_mux_5_nl
      , 1'b1}) + conv_s2u_12_13({10'b1000000000 , return_mult_generic_AC_RND_CONV_false_exp_mux1h_18_nl
      , 1'b1});
  assign acc_28_nl = nl_acc_28_nl[12:0];
  assign z_out_39 = readslicef_13_12_1(acc_28_nl);
  assign stage_u_add_or_4_nl = (fsm_output[4]) | or_dcpl_401 | (fsm_output[29]) |
      return_extract_26_exception_or_3_cse;
  assign stage_u_add_mux1h_8_nl = MUX1HOT_v_16_3_2(16'b1100111111111111, out_u_rsci_q_d,
      in_u_rsci_q_d, {stage_u_add_or_4_nl , (fsm_output[5]) , (fsm_output[30])});
  assign stage_u_add_or_5_nl = (~((fsm_output[4]) | or_dcpl_401 | (fsm_output[29])
      | return_extract_26_exception_or_3_cse)) | (fsm_output[5]) | (fsm_output[30]);
  assign stage_u_add_mux1h_9_nl = MUX1HOT_v_2_5_2((out_u_rsci_q_d[15:14]), BUTTERFLY_1_else_3_else_acc_4_itm_15_14,
      (in_u_rsci_q_d[15:14]), (~ (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0[4:3])),
      (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0[4:3]), {(fsm_output[4])
      , or_dcpl_401 , (fsm_output[29]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_extract_26_exception_or_3_cse});
  assign stage_u_add_mux1h_10_nl = MUX1HOT_v_3_5_2((out_u_rsci_q_d[13:11]), BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_0,
      (in_u_rsci_q_d[13:11]), (~ (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0[2:0])),
      (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_0[2:0]), {(fsm_output[4])
      , or_dcpl_401 , (fsm_output[29]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_extract_26_exception_or_3_cse});
  assign stage_u_add_mux1h_11_nl = MUX1HOT_s_1_5_2((out_u_rsci_q_d[10]), BUTTERFLY_1_else_3_else_acc_4_itm_13_0_rsp_1,
      (in_u_rsci_q_d[10]), (~ (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1[1])),
      (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1[1]), {(fsm_output[4])
      , or_dcpl_401 , (fsm_output[29]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_extract_26_exception_or_3_cse});
  assign stage_u_add_mux1h_12_nl = MUX1HOT_s_1_5_2((out_u_rsci_q_d[9]), (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[4]),
      (in_u_rsci_q_d[9]), (~ (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1[0])),
      (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_1[0]), {(fsm_output[4])
      , or_dcpl_401 , (fsm_output[29]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_extract_26_exception_or_3_cse});
  assign stage_u_add_mux1h_13_nl = MUX1HOT_v_4_5_2((out_u_rsci_q_d[8:5]), (reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd[3:0]),
      (in_u_rsci_q_d[8:5]), (~ (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[8:5])),
      (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[8:5]), {(fsm_output[4])
      , or_dcpl_401 , (fsm_output[29]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_extract_26_exception_or_3_cse});
  assign stage_u_add_mux1h_14_nl = MUX1HOT_v_5_5_2((out_u_rsci_q_d[4:0]), reg_BUTTERFLY_1_else_3_else_acc_4_3_ftd_1,
      (in_u_rsci_q_d[4:0]), (~ (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[4:0])),
      (BUTTERFLY_1_else_1_if_slc_in_u_16_15_0_ncse_sva_rsp_2[4:0]), {(fsm_output[4])
      , or_dcpl_401 , (fsm_output[29]) , return_add_generic_AC_RND_CONV_false_15_e_dif_sat_or_cse
      , return_extract_26_exception_or_3_cse});
  assign nl_acc_29_nl = ({1'b1 , stage_u_add_mux1h_8_nl , stage_u_add_or_5_nl}) +
      conv_u2u_17_18({stage_u_add_mux1h_9_nl , stage_u_add_mux1h_10_nl , stage_u_add_mux1h_11_nl
      , stage_u_add_mux1h_12_nl , stage_u_add_mux1h_13_nl , stage_u_add_mux1h_14_nl
      , 1'b1});
  assign acc_29_nl = nl_acc_29_nl[17:0];
  assign z_out_40 = readslicef_18_17_1(acc_29_nl);
  assign return_mult_generic_AC_RND_CONV_false_2_exp_mux_3_nl = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qr_10_1_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_19_e_r_qr_10_1_lpi_3_dfm_1, fsm_output[39]);
  assign return_mult_generic_AC_RND_CONV_false_2_exp_mux_4_nl = MUX_s_1_2_2(return_add_generic_AC_RND_CONV_false_6_e_r_qr_0_lpi_3_dfm_1,
      return_add_generic_AC_RND_CONV_false_19_e_r_qr_0_lpi_3_dfm_1, fsm_output[39]);
  assign nl_acc_31_nl = conv_u2u_12_13({return_mult_generic_AC_RND_CONV_false_2_exp_mux_3_nl
      , return_mult_generic_AC_RND_CONV_false_2_exp_mux_4_nl , 1'b1}) + conv_u2u_2_13({(~
      BUTTERFLY_1_fiy_slc_BUTTERFLY_1_fiy_acc_1_sdt_9_itm) , 1'b1});
  assign acc_31_nl = nl_acc_31_nl[12:0];
  assign z_out_44 = readslicef_13_12_1(acc_31_nl);
  assign BUTTERFLY_else_2_mux_14_nl = MUX_v_6_2_2(BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_0,
      (z_out_40[16:11]), return_extract_26_exception_or_3_cse);
  assign BUTTERFLY_else_2_mux_15_nl = MUX_s_1_2_2(BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_1,
      (z_out_40[10]), return_extract_26_exception_or_3_cse);
  assign BUTTERFLY_else_2_mux_16_nl = MUX_s_1_2_2(reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd,
      (z_out_40[9]), return_extract_26_exception_or_3_cse);
  assign BUTTERFLY_else_2_mux_17_nl = MUX_v_4_2_2(reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1,
      (z_out_40[8:5]), return_extract_26_exception_or_3_cse);
  assign BUTTERFLY_else_2_mux_18_nl = MUX_v_4_2_2(reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2,
      (z_out_40[4:1]), return_extract_26_exception_or_3_cse);
  assign BUTTERFLY_else_2_mux_19_nl = MUX_s_1_2_2(reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3,
      (z_out_40[0]), return_extract_26_exception_or_3_cse);
  assign BUTTERFLY_else_2_BUTTERFLY_else_2_and_6_nl = MUX_v_3_2_2(3'b000, (BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_0[5:3]),
      return_extract_26_exception_or_3_cse);
  assign BUTTERFLY_else_2_mux_20_nl = MUX_v_2_2_2((signext_2_1(BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_0[5])),
      (BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_0[2:1]), return_extract_26_exception_or_3_cse);
  assign BUTTERFLY_else_2_BUTTERFLY_else_2_and_7_nl = (BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_0[0])
      & return_extract_26_exception_or_3_cse;
  assign BUTTERFLY_else_2_BUTTERFLY_else_2_and_8_nl = BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_1
      & return_extract_26_exception_or_3_cse;
  assign BUTTERFLY_else_2_BUTTERFLY_else_2_and_9_nl = reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd
      & return_extract_26_exception_or_3_cse;
  assign BUTTERFLY_else_2_BUTTERFLY_else_2_and_10_nl = MUX_v_4_2_2(4'b0000, reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_1,
      return_extract_26_exception_or_3_cse);
  assign BUTTERFLY_else_2_BUTTERFLY_else_2_and_11_nl = MUX_v_4_2_2(4'b0000, reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_2,
      return_extract_26_exception_or_3_cse);
  assign BUTTERFLY_else_2_mux_21_nl = MUX_s_1_2_2((BUTTERFLY_1_else_2_acc_1_psp_16_0_sva_rsp_0[5]),
      reg_BUTTERFLY_1_else_2_acc_1_psp_16_0_2_ftd_3, return_extract_26_exception_or_3_cse);
  assign nl_z_out_45 = conv_s2u_17_18({BUTTERFLY_else_2_mux_14_nl , BUTTERFLY_else_2_mux_15_nl
      , BUTTERFLY_else_2_mux_16_nl , BUTTERFLY_else_2_mux_17_nl , BUTTERFLY_else_2_mux_18_nl
      , BUTTERFLY_else_2_mux_19_nl}) + conv_s2u_17_18({BUTTERFLY_else_2_BUTTERFLY_else_2_and_6_nl
      , BUTTERFLY_else_2_mux_20_nl , BUTTERFLY_else_2_BUTTERFLY_else_2_and_7_nl ,
      BUTTERFLY_else_2_BUTTERFLY_else_2_and_8_nl , BUTTERFLY_else_2_BUTTERFLY_else_2_and_9_nl
      , BUTTERFLY_else_2_BUTTERFLY_else_2_and_10_nl , BUTTERFLY_else_2_BUTTERFLY_else_2_and_11_nl
      , BUTTERFLY_else_2_mux_21_nl});
  assign z_out_45 = nl_z_out_45[17:0];
  assign z_out_9 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_11,
      (return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_5_cse[9:0]),
      reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd);
  assign return_add_generic_AC_RND_CONV_false_mux_36_nl = MUX_s_1_2_2(reg_return_add_generic_AC_RND_CONV_false_10_res_rounded_ftd,
      (z_out_6[53]), return_extract_26_exception_or_3_cse);
  assign z_out_10 = MUX_v_10_2_2(return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_11,
      (return_add_generic_AC_RND_CONV_false_return_add_generic_AC_RND_CONV_false_and_5_cse[9:0]),
      return_add_generic_AC_RND_CONV_false_mux_36_nl);
  assign z_out_11 = MUX_v_51_2_2(stage_PE_1_gm_re_d_mux_cse, stage_PE_1_gm_im_d_mux_2_cse,
      or_590_cse);
  assign return_mult_generic_AC_RND_CONV_false_if_mux_6_ssc = MUX_s_1_2_2(return_extract_12_return_extract_12_or_1_cse_sva_1,
      return_extract_44_return_extract_44_or_1_cse_sva_1, fsm_output[35]);

  function automatic [8:0] div_9_u9_u16;
    input [8:0] l;
    input [15:0] r;
    reg [8:0] rdiv;
    reg [16:0] diff;
    reg [17:0] diff_tmp;
    reg [24:0] lbuf;
    integer i; 
  begin
    lbuf = 25'b0;
    lbuf[8:0] = l;
    for(i=8; i>=0; i=i-1)
    begin
      diff_tmp = (lbuf[24:8] - {1'b0,r});
      diff = diff_tmp[16:0];
      rdiv[i] = ~diff[16];
      if(diff[16] == 0)
        lbuf[24:8] = diff;
      lbuf[24:1] = lbuf[23:0];
    end
    div_9_u9_u16 = rdiv;
  end
  endfunction


  function automatic  MUX1HOT_s_1_10_2;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [9:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    MUX1HOT_s_1_10_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_11_2;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [10:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    MUX1HOT_s_1_11_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_12_2;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [11:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    MUX1HOT_s_1_12_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_13_2;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [12:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    MUX1HOT_s_1_13_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_14_2;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [13:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    MUX1HOT_s_1_14_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_15_2;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [14:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    MUX1HOT_s_1_15_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_16_2;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [15:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    MUX1HOT_s_1_16_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_17_2;
    input  input_16;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [16:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    MUX1HOT_s_1_17_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_18_2;
    input  input_17;
    input  input_16;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [17:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    MUX1HOT_s_1_18_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_20_2;
    input  input_19;
    input  input_18;
    input  input_17;
    input  input_16;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [19:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    result = result | (input_18 & sel[18]);
    result = result | (input_19 & sel[19]);
    MUX1HOT_s_1_20_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_22_2;
    input  input_21;
    input  input_20;
    input  input_19;
    input  input_18;
    input  input_17;
    input  input_16;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [21:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    result = result | (input_18 & sel[18]);
    result = result | (input_19 & sel[19]);
    result = result | (input_20 & sel[20]);
    result = result | (input_21 & sel[21]);
    MUX1HOT_s_1_22_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_30_2;
    input  input_29;
    input  input_28;
    input  input_27;
    input  input_26;
    input  input_25;
    input  input_24;
    input  input_23;
    input  input_22;
    input  input_21;
    input  input_20;
    input  input_19;
    input  input_18;
    input  input_17;
    input  input_16;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [29:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    result = result | (input_18 & sel[18]);
    result = result | (input_19 & sel[19]);
    result = result | (input_20 & sel[20]);
    result = result | (input_21 & sel[21]);
    result = result | (input_22 & sel[22]);
    result = result | (input_23 & sel[23]);
    result = result | (input_24 & sel[24]);
    result = result | (input_25 & sel[25]);
    result = result | (input_26 & sel[26]);
    result = result | (input_27 & sel[27]);
    result = result | (input_28 & sel[28]);
    result = result | (input_29 & sel[29]);
    MUX1HOT_s_1_30_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_5_2;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [4:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_6_2;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [5:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_7_2;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [6:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_8_2;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [7:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    MUX1HOT_s_1_8_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_9_2;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [8:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    MUX1HOT_s_1_9_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_13_2;
    input [9:0] input_12;
    input [9:0] input_11;
    input [9:0] input_10;
    input [9:0] input_9;
    input [9:0] input_8;
    input [9:0] input_7;
    input [9:0] input_6;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [12:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    result = result | (input_3 & {10{sel[3]}});
    result = result | (input_4 & {10{sel[4]}});
    result = result | (input_5 & {10{sel[5]}});
    result = result | (input_6 & {10{sel[6]}});
    result = result | (input_7 & {10{sel[7]}});
    result = result | (input_8 & {10{sel[8]}});
    result = result | (input_9 & {10{sel[9]}});
    result = result | (input_10 & {10{sel[10]}});
    result = result | (input_11 & {10{sel[11]}});
    result = result | (input_12 & {10{sel[12]}});
    MUX1HOT_v_10_13_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_3_2;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [2:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    MUX1HOT_v_10_3_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_5_2;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [4:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    result = result | (input_3 & {10{sel[3]}});
    result = result | (input_4 & {10{sel[4]}});
    MUX1HOT_v_10_5_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_6_2;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [5:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | (input_1 & {10{sel[1]}});
    result = result | (input_2 & {10{sel[2]}});
    result = result | (input_3 & {10{sel[3]}});
    result = result | (input_4 & {10{sel[4]}});
    result = result | (input_5 & {10{sel[5]}});
    MUX1HOT_v_10_6_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_13_2;
    input [10:0] input_12;
    input [10:0] input_11;
    input [10:0] input_10;
    input [10:0] input_9;
    input [10:0] input_8;
    input [10:0] input_7;
    input [10:0] input_6;
    input [10:0] input_5;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [12:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    result = result | (input_3 & {11{sel[3]}});
    result = result | (input_4 & {11{sel[4]}});
    result = result | (input_5 & {11{sel[5]}});
    result = result | (input_6 & {11{sel[6]}});
    result = result | (input_7 & {11{sel[7]}});
    result = result | (input_8 & {11{sel[8]}});
    result = result | (input_9 & {11{sel[9]}});
    result = result | (input_10 & {11{sel[10]}});
    result = result | (input_11 & {11{sel[11]}});
    result = result | (input_12 & {11{sel[12]}});
    MUX1HOT_v_11_13_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_3_2;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [2:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    MUX1HOT_v_11_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_5_2;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [4:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    MUX1HOT_v_2_5_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_6_2;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [5:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    MUX1HOT_v_2_6_2 = result;
  end
  endfunction


  function automatic [29:0] MUX1HOT_v_30_12_2;
    input [29:0] input_11;
    input [29:0] input_10;
    input [29:0] input_9;
    input [29:0] input_8;
    input [29:0] input_7;
    input [29:0] input_6;
    input [29:0] input_5;
    input [29:0] input_4;
    input [29:0] input_3;
    input [29:0] input_2;
    input [29:0] input_1;
    input [29:0] input_0;
    input [11:0] sel;
    reg [29:0] result;
  begin
    result = input_0 & {30{sel[0]}};
    result = result | (input_1 & {30{sel[1]}});
    result = result | (input_2 & {30{sel[2]}});
    result = result | (input_3 & {30{sel[3]}});
    result = result | (input_4 & {30{sel[4]}});
    result = result | (input_5 & {30{sel[5]}});
    result = result | (input_6 & {30{sel[6]}});
    result = result | (input_7 & {30{sel[7]}});
    result = result | (input_8 & {30{sel[8]}});
    result = result | (input_9 & {30{sel[9]}});
    result = result | (input_10 & {30{sel[10]}});
    result = result | (input_11 & {30{sel[11]}});
    MUX1HOT_v_30_12_2 = result;
  end
  endfunction


  function automatic [32:0] MUX1HOT_v_33_5_2;
    input [32:0] input_4;
    input [32:0] input_3;
    input [32:0] input_2;
    input [32:0] input_1;
    input [32:0] input_0;
    input [4:0] sel;
    reg [32:0] result;
  begin
    result = input_0 & {33{sel[0]}};
    result = result | (input_1 & {33{sel[1]}});
    result = result | (input_2 & {33{sel[2]}});
    result = result | (input_3 & {33{sel[3]}});
    result = result | (input_4 & {33{sel[4]}});
    MUX1HOT_v_33_5_2 = result;
  end
  endfunction


  function automatic [36:0] MUX1HOT_v_37_5_2;
    input [36:0] input_4;
    input [36:0] input_3;
    input [36:0] input_2;
    input [36:0] input_1;
    input [36:0] input_0;
    input [4:0] sel;
    reg [36:0] result;
  begin
    result = input_0 & {37{sel[0]}};
    result = result | (input_1 & {37{sel[1]}});
    result = result | (input_2 & {37{sel[2]}});
    result = result | (input_3 & {37{sel[3]}});
    result = result | (input_4 & {37{sel[4]}});
    MUX1HOT_v_37_5_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_10_2;
    input [2:0] input_9;
    input [2:0] input_8;
    input [2:0] input_7;
    input [2:0] input_6;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [9:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    result = result | (input_5 & {3{sel[5]}});
    result = result | (input_6 & {3{sel[6]}});
    result = result | (input_7 & {3{sel[7]}});
    result = result | (input_8 & {3{sel[8]}});
    result = result | (input_9 & {3{sel[9]}});
    MUX1HOT_v_3_10_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_17_2;
    input [2:0] input_16;
    input [2:0] input_15;
    input [2:0] input_14;
    input [2:0] input_13;
    input [2:0] input_12;
    input [2:0] input_11;
    input [2:0] input_10;
    input [2:0] input_9;
    input [2:0] input_8;
    input [2:0] input_7;
    input [2:0] input_6;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [16:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    result = result | (input_5 & {3{sel[5]}});
    result = result | (input_6 & {3{sel[6]}});
    result = result | (input_7 & {3{sel[7]}});
    result = result | (input_8 & {3{sel[8]}});
    result = result | (input_9 & {3{sel[9]}});
    result = result | (input_10 & {3{sel[10]}});
    result = result | (input_11 & {3{sel[11]}});
    result = result | (input_12 & {3{sel[12]}});
    result = result | (input_13 & {3{sel[13]}});
    result = result | (input_14 & {3{sel[14]}});
    result = result | (input_15 & {3{sel[15]}});
    result = result | (input_16 & {3{sel[16]}});
    MUX1HOT_v_3_17_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_5_2;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [4:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    MUX1HOT_v_3_5_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_6_2;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [5:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    result = result | (input_5 & {3{sel[5]}});
    MUX1HOT_v_3_6_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_7_2;
    input [2:0] input_6;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [6:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    result = result | (input_5 & {3{sel[5]}});
    result = result | (input_6 & {3{sel[6]}});
    MUX1HOT_v_3_7_2 = result;
  end
  endfunction


  function automatic [44:0] MUX1HOT_v_45_13_2;
    input [44:0] input_12;
    input [44:0] input_11;
    input [44:0] input_10;
    input [44:0] input_9;
    input [44:0] input_8;
    input [44:0] input_7;
    input [44:0] input_6;
    input [44:0] input_5;
    input [44:0] input_4;
    input [44:0] input_3;
    input [44:0] input_2;
    input [44:0] input_1;
    input [44:0] input_0;
    input [12:0] sel;
    reg [44:0] result;
  begin
    result = input_0 & {45{sel[0]}};
    result = result | (input_1 & {45{sel[1]}});
    result = result | (input_2 & {45{sel[2]}});
    result = result | (input_3 & {45{sel[3]}});
    result = result | (input_4 & {45{sel[4]}});
    result = result | (input_5 & {45{sel[5]}});
    result = result | (input_6 & {45{sel[6]}});
    result = result | (input_7 & {45{sel[7]}});
    result = result | (input_8 & {45{sel[8]}});
    result = result | (input_9 & {45{sel[9]}});
    result = result | (input_10 & {45{sel[10]}});
    result = result | (input_11 & {45{sel[11]}});
    result = result | (input_12 & {45{sel[12]}});
    MUX1HOT_v_45_13_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_12_2;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [11:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    MUX1HOT_v_4_12_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_20_2;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [19:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    MUX1HOT_v_4_20_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_5_2;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [4:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    MUX1HOT_v_4_5_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_6_2;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [5:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    MUX1HOT_v_4_6_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_7_2;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [6:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    MUX1HOT_v_4_7_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_8_2;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [7:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    MUX1HOT_v_4_8_2 = result;
  end
  endfunction


  function automatic [49:0] MUX1HOT_v_50_11_2;
    input [49:0] input_10;
    input [49:0] input_9;
    input [49:0] input_8;
    input [49:0] input_7;
    input [49:0] input_6;
    input [49:0] input_5;
    input [49:0] input_4;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [10:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    result = result | (input_3 & {50{sel[3]}});
    result = result | (input_4 & {50{sel[4]}});
    result = result | (input_5 & {50{sel[5]}});
    result = result | (input_6 & {50{sel[6]}});
    result = result | (input_7 & {50{sel[7]}});
    result = result | (input_8 & {50{sel[8]}});
    result = result | (input_9 & {50{sel[9]}});
    result = result | (input_10 & {50{sel[10]}});
    MUX1HOT_v_50_11_2 = result;
  end
  endfunction


  function automatic [49:0] MUX1HOT_v_50_12_2;
    input [49:0] input_11;
    input [49:0] input_10;
    input [49:0] input_9;
    input [49:0] input_8;
    input [49:0] input_7;
    input [49:0] input_6;
    input [49:0] input_5;
    input [49:0] input_4;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [11:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    result = result | (input_3 & {50{sel[3]}});
    result = result | (input_4 & {50{sel[4]}});
    result = result | (input_5 & {50{sel[5]}});
    result = result | (input_6 & {50{sel[6]}});
    result = result | (input_7 & {50{sel[7]}});
    result = result | (input_8 & {50{sel[8]}});
    result = result | (input_9 & {50{sel[9]}});
    result = result | (input_10 & {50{sel[10]}});
    result = result | (input_11 & {50{sel[11]}});
    MUX1HOT_v_50_12_2 = result;
  end
  endfunction


  function automatic [49:0] MUX1HOT_v_50_15_2;
    input [49:0] input_14;
    input [49:0] input_13;
    input [49:0] input_12;
    input [49:0] input_11;
    input [49:0] input_10;
    input [49:0] input_9;
    input [49:0] input_8;
    input [49:0] input_7;
    input [49:0] input_6;
    input [49:0] input_5;
    input [49:0] input_4;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [14:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    result = result | (input_3 & {50{sel[3]}});
    result = result | (input_4 & {50{sel[4]}});
    result = result | (input_5 & {50{sel[5]}});
    result = result | (input_6 & {50{sel[6]}});
    result = result | (input_7 & {50{sel[7]}});
    result = result | (input_8 & {50{sel[8]}});
    result = result | (input_9 & {50{sel[9]}});
    result = result | (input_10 & {50{sel[10]}});
    result = result | (input_11 & {50{sel[11]}});
    result = result | (input_12 & {50{sel[12]}});
    result = result | (input_13 & {50{sel[13]}});
    result = result | (input_14 & {50{sel[14]}});
    MUX1HOT_v_50_15_2 = result;
  end
  endfunction


  function automatic [49:0] MUX1HOT_v_50_3_2;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [2:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    MUX1HOT_v_50_3_2 = result;
  end
  endfunction


  function automatic [49:0] MUX1HOT_v_50_4_2;
    input [49:0] input_3;
    input [49:0] input_2;
    input [49:0] input_1;
    input [49:0] input_0;
    input [3:0] sel;
    reg [49:0] result;
  begin
    result = input_0 & {50{sel[0]}};
    result = result | (input_1 & {50{sel[1]}});
    result = result | (input_2 & {50{sel[2]}});
    result = result | (input_3 & {50{sel[3]}});
    MUX1HOT_v_50_4_2 = result;
  end
  endfunction


  function automatic [50:0] MUX1HOT_v_51_3_2;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [2:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | (input_1 & {51{sel[1]}});
    result = result | (input_2 & {51{sel[2]}});
    MUX1HOT_v_51_3_2 = result;
  end
  endfunction


  function automatic [50:0] MUX1HOT_v_51_4_2;
    input [50:0] input_3;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [3:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | (input_1 & {51{sel[1]}});
    result = result | (input_2 & {51{sel[2]}});
    result = result | (input_3 & {51{sel[3]}});
    MUX1HOT_v_51_4_2 = result;
  end
  endfunction


  function automatic [50:0] MUX1HOT_v_51_5_2;
    input [50:0] input_4;
    input [50:0] input_3;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [4:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | (input_1 & {51{sel[1]}});
    result = result | (input_2 & {51{sel[2]}});
    result = result | (input_3 & {51{sel[3]}});
    result = result | (input_4 & {51{sel[4]}});
    MUX1HOT_v_51_5_2 = result;
  end
  endfunction


  function automatic [50:0] MUX1HOT_v_51_8_2;
    input [50:0] input_7;
    input [50:0] input_6;
    input [50:0] input_5;
    input [50:0] input_4;
    input [50:0] input_3;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [7:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | (input_1 & {51{sel[1]}});
    result = result | (input_2 & {51{sel[2]}});
    result = result | (input_3 & {51{sel[3]}});
    result = result | (input_4 & {51{sel[4]}});
    result = result | (input_5 & {51{sel[5]}});
    result = result | (input_6 & {51{sel[6]}});
    result = result | (input_7 & {51{sel[7]}});
    MUX1HOT_v_51_8_2 = result;
  end
  endfunction


  function automatic [51:0] MUX1HOT_v_52_8_2;
    input [51:0] input_7;
    input [51:0] input_6;
    input [51:0] input_5;
    input [51:0] input_4;
    input [51:0] input_3;
    input [51:0] input_2;
    input [51:0] input_1;
    input [51:0] input_0;
    input [7:0] sel;
    reg [51:0] result;
  begin
    result = input_0 & {52{sel[0]}};
    result = result | (input_1 & {52{sel[1]}});
    result = result | (input_2 & {52{sel[2]}});
    result = result | (input_3 & {52{sel[3]}});
    result = result | (input_4 & {52{sel[4]}});
    result = result | (input_5 & {52{sel[5]}});
    result = result | (input_6 & {52{sel[6]}});
    result = result | (input_7 & {52{sel[7]}});
    MUX1HOT_v_52_8_2 = result;
  end
  endfunction


  function automatic [52:0] MUX1HOT_v_53_3_2;
    input [52:0] input_2;
    input [52:0] input_1;
    input [52:0] input_0;
    input [2:0] sel;
    reg [52:0] result;
  begin
    result = input_0 & {53{sel[0]}};
    result = result | (input_1 & {53{sel[1]}});
    result = result | (input_2 & {53{sel[2]}});
    MUX1HOT_v_53_3_2 = result;
  end
  endfunction


  function automatic [56:0] MUX1HOT_v_57_3_2;
    input [56:0] input_2;
    input [56:0] input_1;
    input [56:0] input_0;
    input [2:0] sel;
    reg [56:0] result;
  begin
    result = input_0 & {57{sel[0]}};
    result = result | (input_1 & {57{sel[1]}});
    result = result | (input_2 & {57{sel[2]}});
    MUX1HOT_v_57_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_13_2;
    input [4:0] input_12;
    input [4:0] input_11;
    input [4:0] input_10;
    input [4:0] input_9;
    input [4:0] input_8;
    input [4:0] input_7;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [12:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    result = result | (input_7 & {5{sel[7]}});
    result = result | (input_8 & {5{sel[8]}});
    result = result | (input_9 & {5{sel[9]}});
    result = result | (input_10 & {5{sel[10]}});
    result = result | (input_11 & {5{sel[11]}});
    result = result | (input_12 & {5{sel[12]}});
    MUX1HOT_v_5_13_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_4_2;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [3:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    MUX1HOT_v_5_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_5_2;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [4:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    MUX1HOT_v_5_5_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_6_2;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [5:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    MUX1HOT_v_5_6_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_7_2;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [6:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    MUX1HOT_v_5_7_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_13_2;
    input [5:0] input_12;
    input [5:0] input_11;
    input [5:0] input_10;
    input [5:0] input_9;
    input [5:0] input_8;
    input [5:0] input_7;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [12:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    result = result | (input_6 & {6{sel[6]}});
    result = result | (input_7 & {6{sel[7]}});
    result = result | (input_8 & {6{sel[8]}});
    result = result | (input_9 & {6{sel[9]}});
    result = result | (input_10 & {6{sel[10]}});
    result = result | (input_11 & {6{sel[11]}});
    result = result | (input_12 & {6{sel[12]}});
    MUX1HOT_v_6_13_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_5_2;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [4:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    MUX1HOT_v_6_5_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_6_2;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [5:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    MUX1HOT_v_6_6_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_7_2;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [6:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    result = result | (input_6 & {6{sel[6]}});
    MUX1HOT_v_6_7_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_8_2;
    input [5:0] input_7;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [7:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    result = result | (input_6 & {6{sel[6]}});
    result = result | (input_7 & {6{sel[7]}});
    MUX1HOT_v_6_8_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_3_2;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [2:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | (input_1 & {9{sel[1]}});
    result = result | (input_2 & {9{sel[2]}});
    MUX1HOT_v_9_3_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_4_2;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [3:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | (input_1 & {9{sel[1]}});
    result = result | (input_2 & {9{sel[2]}});
    result = result | (input_3 & {9{sel[3]}});
    MUX1HOT_v_9_4_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_5_2;
    input [8:0] input_4;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [4:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | (input_1 & {9{sel[1]}});
    result = result | (input_2 & {9{sel[2]}});
    result = result | (input_3 & {9{sel[3]}});
    result = result | (input_4 & {9{sel[4]}});
    MUX1HOT_v_9_5_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input  sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input  sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input  sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [29:0] MUX_v_30_2_2;
    input [29:0] input_0;
    input [29:0] input_1;
    input  sel;
    reg [29:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_30_2_2 = result;
  end
  endfunction


  function automatic [32:0] MUX_v_33_2_2;
    input [32:0] input_0;
    input [32:0] input_1;
    input  sel;
    reg [32:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_33_2_2 = result;
  end
  endfunction


  function automatic [36:0] MUX_v_37_2_2;
    input [36:0] input_0;
    input [36:0] input_1;
    input  sel;
    reg [36:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_37_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [49:0] MUX_v_50_2_2;
    input [49:0] input_0;
    input [49:0] input_1;
    input  sel;
    reg [49:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_50_2_2 = result;
  end
  endfunction


  function automatic [50:0] MUX_v_51_2_2;
    input [50:0] input_0;
    input [50:0] input_1;
    input  sel;
    reg [50:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_51_2_2 = result;
  end
  endfunction


  function automatic [51:0] MUX_v_52_2_2;
    input [51:0] input_0;
    input [51:0] input_1;
    input  sel;
    reg [51:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_52_2_2 = result;
  end
  endfunction


  function automatic [55:0] MUX_v_56_2_2;
    input [55:0] input_0;
    input [55:0] input_1;
    input  sel;
    reg [55:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_56_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [10:0] readslicef_12_11_1;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_12_11_1 = tmp[10:0];
  end
  endfunction


  function automatic [0:0] readslicef_12_1_11;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_12_1_11 = tmp[0:0];
  end
  endfunction


  function automatic [11:0] readslicef_13_12_1;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_13_12_1 = tmp[11:0];
  end
  endfunction


  function automatic [0:0] readslicef_13_1_12;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 12;
    readslicef_13_1_12 = tmp[0:0];
  end
  endfunction


  function automatic [12:0] readslicef_14_13_1;
    input [13:0] vector;
    reg [13:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_14_13_1 = tmp[12:0];
  end
  endfunction


  function automatic [16:0] readslicef_18_17_1;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_18_17_1 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_19_18_1;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_19_18_1 = tmp[17:0];
  end
  endfunction


  function automatic [15:0] readslicef_32_16_16;
    input [31:0] vector;
    reg [31:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_32_16_16 = tmp[15:0];
  end
  endfunction


  function automatic [0:0] readslicef_53_1_52;
    input [52:0] vector;
    reg [52:0] tmp;
  begin
    tmp = vector >> 52;
    readslicef_53_1_52 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_54_1_53;
    input [53:0] vector;
    reg [53:0] tmp;
  begin
    tmp = vector >> 53;
    readslicef_54_1_53 = tmp[0:0];
  end
  endfunction


  function automatic [56:0] readslicef_58_57_1;
    input [57:0] vector;
    reg [57:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_58_57_1 = tmp[56:0];
  end
  endfunction


  function automatic [13:0] signext_14_13;
    input [12:0] vector;
  begin
    signext_14_13= {{1{vector[12]}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input  vector;
  begin
    signext_2_1= {{1{vector}}, vector};
  end
  endfunction


  function automatic [32:0] signext_33_1;
    input  vector;
  begin
    signext_33_1= {{32{vector}}, vector};
  end
  endfunction


  function automatic [44:0] signext_45_11;
    input [10:0] vector;
  begin
    signext_45_11= {{34{vector[10]}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_2;
    input [1:0] vector;
  begin
    signext_4_2= {{2{vector[1]}}, vector};
  end
  endfunction


  function automatic [54:0] signext_55_54;
    input [53:0] vector;
  begin
    signext_55_54= {{1{vector[53]}}, vector};
  end
  endfunction


  function automatic [5:0] signext_6_1;
    input  vector;
  begin
    signext_6_1= {{5{vector}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2u_7_13 ;
    input [6:0]  vector ;
  begin
    conv_s2u_7_13 = {{6{vector[6]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2u_8_12 ;
    input [7:0]  vector ;
  begin
    conv_s2u_8_12 = {{4{vector[7]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2u_8_13 ;
    input [7:0]  vector ;
  begin
    conv_s2u_8_13 = {{5{vector[7]}}, vector};
  end
  endfunction


  function automatic [13:0] conv_s2u_8_14 ;
    input [7:0]  vector ;
  begin
    conv_s2u_8_14 = {{6{vector[7]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [12:0] conv_s2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_s2u_12_13 = {vector[11], vector};
  end
  endfunction


  function automatic [13:0] conv_s2u_13_14 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_14 = {vector[12], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_19 = {vector[17], vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [14:0] conv_u2s_14_15 ;
    input [13:0]  vector ;
  begin
    conv_u2s_14_15 =  {1'b0, vector};
  end
  endfunction


  function automatic [53:0] conv_u2s_53_54 ;
    input [52:0]  vector ;
  begin
    conv_u2s_53_54 =  {1'b0, vector};
  end
  endfunction


  function automatic [53:0] conv_u2u_1_54 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_54 = {{53{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_2_13 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_13 = {{11{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_4_11 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_11 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_11_13 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_13 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_u2u_12_13 = {1'b0, vector};
  end
  endfunction


  function automatic [13:0] conv_u2u_13_14 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_14 = {1'b0, vector};
  end
  endfunction


  function automatic [15:0] conv_u2u_14_16 ;
    input [13:0]  vector ;
  begin
    conv_u2u_14_16 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [17:0] conv_u2u_14_18 ;
    input [13:0]  vector ;
  begin
    conv_u2u_14_18 = {{4{1'b0}}, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_16_32 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_32 = {{16{1'b0}}, vector};
  end
  endfunction


  function automatic [17:0] conv_u2u_17_18 ;
    input [16:0]  vector ;
  begin
    conv_u2u_17_18 = {1'b0, vector};
  end
  endfunction


  function automatic [18:0] conv_u2u_17_19 ;
    input [16:0]  vector ;
  begin
    conv_u2u_17_19 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_28_32 ;
    input [27:0]  vector ;
  begin
    conv_u2u_28_32 = {{4{1'b0}}, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_30_32 ;
    input [29:0]  vector ;
  begin
    conv_u2u_30_32 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [52:0] conv_u2u_52_53 ;
    input [51:0]  vector ;
  begin
    conv_u2u_52_53 = {1'b0, vector};
  end
  endfunction


  function automatic [53:0] conv_u2u_53_54 ;
    input [52:0]  vector ;
  begin
    conv_u2u_53_54 = {1'b0, vector};
  end
  endfunction


  function automatic [57:0] conv_u2u_57_58 ;
    input [56:0]  vector ;
  begin
    conv_u2u_57_58 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage_struct
// ------------------------------------------------------------------


module stage_struct (
  clk, rst, arst_n, ap_start_rsc_dat, ap_start_rsc_vld, ap_start_rsc_rdy, ap_done_rsc_dat,
      ap_done_rsc_vld, ap_done_rsc_rdy, mode1_rsc_dat, mode1_triosy_lz, in_f_d_rsc_adr,
      in_f_d_rsc_d, in_f_d_rsc_we, in_f_d_rsc_q, in_f_d_rsc_en, in_f_d_triosy_lz,
      in_u_rsc_adr, in_u_rsc_d, in_u_rsc_we, in_u_rsc_q, in_u_rsc_en, in_u_triosy_lz,
      out_f_d_rsc_adr, out_f_d_rsc_d, out_f_d_rsc_we, out_f_d_rsc_q, out_f_d_rsc_en,
      out_f_d_triosy_lz, out_u_rsc_adr, out_u_rsc_d, out_u_rsc_we, out_u_rsc_q, out_u_rsc_en,
      out_u_triosy_lz, out1_rsc_dat_u, out1_rsc_dat_d, out1_rsc_vld, out1_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input [15:0] mode1_rsc_dat;
  output mode1_triosy_lz;
  output [9:0] in_f_d_rsc_adr;
  output [63:0] in_f_d_rsc_d;
  output in_f_d_rsc_we;
  input [63:0] in_f_d_rsc_q;
  output in_f_d_rsc_en;
  output in_f_d_triosy_lz;
  output [9:0] in_u_rsc_adr;
  output [15:0] in_u_rsc_d;
  output in_u_rsc_we;
  input [15:0] in_u_rsc_q;
  output in_u_rsc_en;
  output in_u_triosy_lz;
  output [9:0] out_f_d_rsc_adr;
  output [63:0] out_f_d_rsc_d;
  output out_f_d_rsc_we;
  input [63:0] out_f_d_rsc_q;
  output out_f_d_rsc_en;
  output out_f_d_triosy_lz;
  output [9:0] out_u_rsc_adr;
  output [15:0] out_u_rsc_d;
  output out_u_rsc_we;
  input [15:0] out_u_rsc_q;
  output out_u_rsc_en;
  output out_u_triosy_lz;
  output [15:0] out1_rsc_dat_u;
  output [63:0] out1_rsc_dat_d;
  output out1_rsc_vld;
  input out1_rsc_rdy;


  // Interconnect Declarations
  wire [9:0] in_f_d_rsci_adr_d;
  wire [63:0] in_f_d_rsci_d_d;
  wire in_f_d_rsci_en_d;
  wire [63:0] in_f_d_rsci_q_d;
  wire in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [9:0] in_u_rsci_adr_d;
  wire [15:0] in_u_rsci_d_d;
  wire in_u_rsci_en_d;
  wire [15:0] in_u_rsci_q_d;
  wire in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [9:0] out_f_d_rsci_adr_d;
  wire [63:0] out_f_d_rsci_d_d;
  wire out_f_d_rsci_en_d;
  wire [63:0] out_f_d_rsci_q_d;
  wire out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [9:0] out_u_rsci_adr_d;
  wire [15:0] out_u_rsci_d_d;
  wire out_u_rsci_en_d;
  wire [15:0] out_u_rsci_q_d;
  wire out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [79:0] out1_rsc_dat;
  wire in_f_d_rsci_we_d_iff;
  wire in_u_rsci_we_d_iff;
  wire out_f_d_rsci_we_d_iff;
  wire out_u_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_4_64_10_1024_1024_64_5_gen
      in_f_d_rsci (
      .en(in_f_d_rsc_en),
      .q(in_f_d_rsc_q),
      .we(in_f_d_rsc_we),
      .d(in_f_d_rsc_d),
      .adr(in_f_d_rsc_adr),
      .adr_d(in_f_d_rsci_adr_d),
      .d_d(in_f_d_rsci_d_d),
      .en_d(in_f_d_rsci_en_d),
      .we_d(in_f_d_rsci_we_d_iff),
      .q_d(in_f_d_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(in_f_d_rsci_we_d_iff)
    );
  stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_5_16_10_1024_1024_16_5_gen
      in_u_rsci (
      .en(in_u_rsc_en),
      .q(in_u_rsc_q),
      .we(in_u_rsc_we),
      .d(in_u_rsc_d),
      .adr(in_u_rsc_adr),
      .adr_d(in_u_rsci_adr_d),
      .d_d(in_u_rsci_d_d),
      .en_d(in_u_rsci_en_d),
      .we_d(in_u_rsci_we_d_iff),
      .q_d(in_u_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(in_u_rsci_we_d_iff)
    );
  stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_6_64_10_1024_1024_64_5_gen
      out_f_d_rsci (
      .en(out_f_d_rsc_en),
      .q(out_f_d_rsc_q),
      .we(out_f_d_rsc_we),
      .d(out_f_d_rsc_d),
      .adr(out_f_d_rsc_adr),
      .adr_d(out_f_d_rsci_adr_d),
      .d_d(out_f_d_rsci_d_d),
      .en_d(out_f_d_rsci_en_d),
      .we_d(out_f_d_rsci_we_d_iff),
      .q_d(out_f_d_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(out_f_d_rsci_we_d_iff)
    );
  stage_ccs_sample_mem_ccs_ram_sync_singleport_rwport_en_7_16_10_1024_1024_16_5_gen
      out_u_rsci (
      .en(out_u_rsc_en),
      .q(out_u_rsc_q),
      .we(out_u_rsc_we),
      .d(out_u_rsc_d),
      .adr(out_u_rsc_adr),
      .adr_d(out_u_rsci_adr_d),
      .d_d(out_u_rsci_d_d),
      .en_d(out_u_rsci_en_d),
      .we_d(out_u_rsci_we_d_iff),
      .q_d(out_u_rsci_q_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(out_u_rsci_we_d_iff)
    );
  stage_run stage_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .ap_start_rsc_dat(ap_start_rsc_dat),
      .ap_start_rsc_vld(ap_start_rsc_vld),
      .ap_start_rsc_rdy(ap_start_rsc_rdy),
      .ap_done_rsc_dat(ap_done_rsc_dat),
      .ap_done_rsc_vld(ap_done_rsc_vld),
      .ap_done_rsc_rdy(ap_done_rsc_rdy),
      .mode1_rsc_dat(mode1_rsc_dat),
      .mode1_triosy_lz(mode1_triosy_lz),
      .in_f_d_triosy_lz(in_f_d_triosy_lz),
      .in_u_triosy_lz(in_u_triosy_lz),
      .out_f_d_triosy_lz(out_f_d_triosy_lz),
      .out_u_triosy_lz(out_u_triosy_lz),
      .out1_rsc_dat(out1_rsc_dat),
      .out1_rsc_vld(out1_rsc_vld),
      .out1_rsc_rdy(out1_rsc_rdy),
      .in_f_d_rsci_adr_d(in_f_d_rsci_adr_d),
      .in_f_d_rsci_d_d(in_f_d_rsci_d_d),
      .in_f_d_rsci_en_d(in_f_d_rsci_en_d),
      .in_f_d_rsci_q_d(in_f_d_rsci_q_d),
      .in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(in_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .in_u_rsci_adr_d(in_u_rsci_adr_d),
      .in_u_rsci_d_d(in_u_rsci_d_d),
      .in_u_rsci_en_d(in_u_rsci_en_d),
      .in_u_rsci_q_d(in_u_rsci_q_d),
      .in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(in_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .out_f_d_rsci_adr_d(out_f_d_rsci_adr_d),
      .out_f_d_rsci_d_d(out_f_d_rsci_d_d),
      .out_f_d_rsci_en_d(out_f_d_rsci_en_d),
      .out_f_d_rsci_q_d(out_f_d_rsci_q_d),
      .out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(out_f_d_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .out_u_rsci_adr_d(out_u_rsci_adr_d),
      .out_u_rsci_d_d(out_u_rsci_d_d),
      .out_u_rsci_en_d(out_u_rsci_en_d),
      .out_u_rsci_q_d(out_u_rsci_q_d),
      .out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(out_u_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .in_f_d_rsci_we_d_pff(in_f_d_rsci_we_d_iff),
      .in_u_rsci_we_d_pff(in_u_rsci_we_d_iff),
      .out_f_d_rsci_we_d_pff(out_f_d_rsci_we_d_iff),
      .out_u_rsci_we_d_pff(out_u_rsci_we_d_iff)
    );
  assign out1_rsc_dat_d = out1_rsc_dat[63:0];
  assign out1_rsc_dat_u = out1_rsc_dat[79:64];
endmodule

// ------------------------------------------------------------------
//  Design Unit:    stage
// ------------------------------------------------------------------


module fiFFNTT (
  clk, rst, arst_n, ap_start_rsc_dat, ap_start_rsc_vld, ap_start_rsc_rdy, ap_done_rsc_dat,
      ap_done_rsc_vld, ap_done_rsc_rdy, mode1_rsc_dat, mode1_triosy_lz, in_f_d_rsc_adr,
      in_f_d_rsc_d, in_f_d_rsc_we, in_f_d_rsc_q, in_f_d_rsc_en, in_f_d_triosy_lz,
      in_u_rsc_adr, in_u_rsc_d, in_u_rsc_we, in_u_rsc_q, in_u_rsc_en, in_u_triosy_lz,
      out_f_d_rsc_adr, out_f_d_rsc_d, out_f_d_rsc_we, out_f_d_rsc_q, out_f_d_rsc_en,
      out_f_d_triosy_lz, out_u_rsc_adr, out_u_rsc_d, out_u_rsc_we, out_u_rsc_q, out_u_rsc_en,
      out_u_triosy_lz, out1_rsc_dat, out1_rsc_vld, out1_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input ap_start_rsc_dat;
  input ap_start_rsc_vld;
  output ap_start_rsc_rdy;
  output ap_done_rsc_dat;
  output ap_done_rsc_vld;
  input ap_done_rsc_rdy;
  input [15:0] mode1_rsc_dat;
  output mode1_triosy_lz;
  output [9:0] in_f_d_rsc_adr;
  output [63:0] in_f_d_rsc_d;
  output in_f_d_rsc_we;
  input [63:0] in_f_d_rsc_q;
  output in_f_d_rsc_en;
  output in_f_d_triosy_lz;
  output [9:0] in_u_rsc_adr;
  output [15:0] in_u_rsc_d;
  output in_u_rsc_we;
  input [15:0] in_u_rsc_q;
  output in_u_rsc_en;
  output in_u_triosy_lz;
  output [9:0] out_f_d_rsc_adr;
  output [63:0] out_f_d_rsc_d;
  output out_f_d_rsc_we;
  input [63:0] out_f_d_rsc_q;
  output out_f_d_rsc_en;
  output out_f_d_triosy_lz;
  output [9:0] out_u_rsc_adr;
  output [15:0] out_u_rsc_d;
  output out_u_rsc_we;
  input [15:0] out_u_rsc_q;
  output out_u_rsc_en;
  output out_u_triosy_lz;
  output [79:0] out1_rsc_dat;
  output out1_rsc_vld;
  input out1_rsc_rdy;


  // Interconnect Declarations
  wire [15:0] out1_rsc_dat_u;
  wire [63:0] out1_rsc_dat_d;


  // Interconnect Declarations for Component Instantiations 
  stage_struct stage_struct_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .ap_start_rsc_dat(ap_start_rsc_dat),
      .ap_start_rsc_vld(ap_start_rsc_vld),
      .ap_start_rsc_rdy(ap_start_rsc_rdy),
      .ap_done_rsc_dat(ap_done_rsc_dat),
      .ap_done_rsc_vld(ap_done_rsc_vld),
      .ap_done_rsc_rdy(ap_done_rsc_rdy),
      .mode1_rsc_dat(mode1_rsc_dat),
      .mode1_triosy_lz(mode1_triosy_lz),
      .in_f_d_rsc_adr(in_f_d_rsc_adr),
      .in_f_d_rsc_d(in_f_d_rsc_d),
      .in_f_d_rsc_we(in_f_d_rsc_we),
      .in_f_d_rsc_q(in_f_d_rsc_q),
      .in_f_d_rsc_en(in_f_d_rsc_en),
      .in_f_d_triosy_lz(in_f_d_triosy_lz),
      .in_u_rsc_adr(in_u_rsc_adr),
      .in_u_rsc_d(in_u_rsc_d),
      .in_u_rsc_we(in_u_rsc_we),
      .in_u_rsc_q(in_u_rsc_q),
      .in_u_rsc_en(in_u_rsc_en),
      .in_u_triosy_lz(in_u_triosy_lz),
      .out_f_d_rsc_adr(out_f_d_rsc_adr),
      .out_f_d_rsc_d(out_f_d_rsc_d),
      .out_f_d_rsc_we(out_f_d_rsc_we),
      .out_f_d_rsc_q(out_f_d_rsc_q),
      .out_f_d_rsc_en(out_f_d_rsc_en),
      .out_f_d_triosy_lz(out_f_d_triosy_lz),
      .out_u_rsc_adr(out_u_rsc_adr),
      .out_u_rsc_d(out_u_rsc_d),
      .out_u_rsc_we(out_u_rsc_we),
      .out_u_rsc_q(out_u_rsc_q),
      .out_u_rsc_en(out_u_rsc_en),
      .out_u_triosy_lz(out_u_triosy_lz),
      .out1_rsc_dat_u(out1_rsc_dat_u),
      .out1_rsc_dat_d(out1_rsc_dat_d),
      .out1_rsc_vld(out1_rsc_vld),
      .out1_rsc_rdy(out1_rsc_rdy)
    );
  assign out1_rsc_dat = {out1_rsc_dat_u , out1_rsc_dat_d};
endmodule



